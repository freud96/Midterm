/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:23 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module cynw_cm_float_mul_inst_cellmath__64_2WWMM_bdw3636473930_bdw (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
wire  inst_cellmath__17,
	inst_cellmath__18,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23,
	inst_cellmath__24,
	inst_cellmath__25,
	inst_cellmath__26,
	inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__32,
	inst_cellmath__33;
wire [9:0] inst_cellmath__34;
wire  inst_cellmath__37,
	inst_cellmath__38,
	inst_cellmath__41,
	inst_cellmath__42;
wire [47:0] inst_cellmath__43;
wire [7:0] inst_cellmath__50,
	inst_cellmath__54;
wire  inst_cellmath__56,
	inst_cellmath__60,
	inst_cellmath__61;
wire N267,N268,N269,N270,N271,N272,N273 
	,N274,N275,N276,N277,N380;
cynw_cm_float_mul_inst_cellmath__33_0_bdw3636473930_bdw cynw_cm_float_mul_I0 (.inst_cellmath__33_0_out0(inst_cellmath__33), .inst_cellmath__33_0_in0(b_sign), .inst_cellmath__33_0_in1(a_sign));
cynw_cm_float_mul_inst_cellmath__26__8__bdw3636473930_bdw cynw_cm_float_mul_I1 (.inst_cellmath__26__8__out0(inst_cellmath__26), .inst_cellmath__26__8__in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_inst_cellmath__17_0_bdw3636473930_bdw cynw_cm_float_mul_I2 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_inst_cellmath__19__5__bdw3636473930_bdw cynw_cm_float_mul_I3 (.inst_cellmath__19__5__out0(inst_cellmath__19), .inst_cellmath__19__5__in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_inst_cellmath__23_0_bdw3636473930_bdw cynw_cm_float_mul_I4 (.inst_cellmath__23_0_out0(inst_cellmath__23), .inst_cellmath__23_0_in0(inst_cellmath__19), .inst_cellmath__23_0_in1(inst_cellmath__17));
cynw_cm_float_mul_inst_cellmath__29__10__bdw3636473930_bdw cynw_cm_float_mul_I5 (.inst_cellmath__29__10__out0({N268}), .inst_cellmath__29__10__in0(inst_cellmath__26), .inst_cellmath__29__10__in1(inst_cellmath__23));
cynw_cm_float_mul_inst_cellmath__25__7__bdw3636473930_bdw cynw_cm_float_mul_I6 (.inst_cellmath__25__7__out0(inst_cellmath__25), .inst_cellmath__25__7__in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_inst_cellmath__18_0_bdw3636473930_bdw cynw_cm_float_mul_I7 (.inst_cellmath__18_0_out0(inst_cellmath__18), .inst_cellmath__18_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_inst_cellmath__20__6__bdw3636473930_bdw cynw_cm_float_mul_I8 (.inst_cellmath__20__6__out0(inst_cellmath__20), .inst_cellmath__20__6__in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}));
cynw_cm_float_mul_inst_cellmath__24_0_bdw3636473930_bdw cynw_cm_float_mul_I9 (.inst_cellmath__24_0_out0(inst_cellmath__24), .inst_cellmath__24_0_in0(inst_cellmath__20), .inst_cellmath__24_0_in1(inst_cellmath__18));
cynw_cm_float_mul_inst_cellmath__29__9__bdw3636473930_bdw cynw_cm_float_mul_I10 (.inst_cellmath__29__9__out0({N267}), .inst_cellmath__29__9__in0(inst_cellmath__25), .inst_cellmath__29__9__in1(inst_cellmath__24));
cynw_cm_float_mul_inst_cellmath__21_0_bdw3636473930_bdw cynw_cm_float_mul_I11 (.inst_cellmath__21_0_out0(inst_cellmath__21), .inst_cellmath__21_0_in0(inst_cellmath__19), .inst_cellmath__21_0_in1(inst_cellmath__17));
cynw_cm_float_mul_inst_cellmath__22_0_bdw3636473930_bdw cynw_cm_float_mul_I12 (.inst_cellmath__22_0_out0(inst_cellmath__22), .inst_cellmath__22_0_in0(inst_cellmath__20), .inst_cellmath__22_0_in1(inst_cellmath__18));
cynw_cm_float_mul_inst_cellmath__29_0_bdw3636473930_bdw cynw_cm_float_mul_I13 (.inst_cellmath__29_0_out0(inst_cellmath__29), .inst_cellmath__29_0_in0({N267}), .inst_cellmath__29_0_in1({N268}), .inst_cellmath__29_0_in2(inst_cellmath__22), .inst_cellmath__29_0_in3(inst_cellmath__21));
cynw_cm_float_mul_inst_cellmath__53_0_bdw3636473930_bdw cynw_cm_float_mul_I14 (.inst_cellmath__53_0_out0(x[31]), .inst_cellmath__53_0_in0(inst_cellmath__33), .inst_cellmath__53_0_in1(inst_cellmath__29));
cynw_cm_float_mul_inst_cellmath__43_0_bdw3636473930_bdw cynw_cm_float_mul_I15 (.inst_cellmath__43_0_out0({inst_cellmath__43[47], inst_cellmath__43[46], inst_cellmath__43[45], inst_cellmath__43[44], inst_cellmath__43[43], inst_cellmath__43[42], inst_cellmath__43[41], inst_cellmath__43[40], inst_cellmath__43[39], inst_cellmath__43[38], inst_cellmath__43[37], inst_cellmath__43[36], inst_cellmath__43[35], inst_cellmath__43[34], inst_cellmath__43[33], inst_cellmath__43[32], inst_cellmath__43[31], inst_cellmath__43[30], inst_cellmath__43[29], inst_cellmath__43[28], inst_cellmath__43[27], inst_cellmath__43[26], inst_cellmath__43[25], inst_cellmath__43[24], inst_cellmath__43[23], inst_cellmath__43[22], inst_cellmath__43[21], inst_cellmath__43[20], inst_cellmath__43[19], inst_cellmath__43[18], inst_cellmath__43[17], inst_cellmath__43[16], inst_cellmath__43[15], inst_cellmath__43[14], inst_cellmath__43[13], inst_cellmath__43[12], inst_cellmath__43[11], inst_cellmath__43[10], inst_cellmath__43[9], inst_cellmath__43[8], inst_cellmath__43[7], inst_cellmath__43[6], inst_cellmath__43[5], inst_cellmath__43[4], inst_cellmath__43[3], inst_cellmath__43[2], inst_cellmath__43[1], inst_cellmath__43[0]}), .inst_cellmath__43_0_in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__43_0_in1({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_inst_cellmath__30__13__bdw3636473930_bdw cynw_cm_float_mul_I16 (.inst_cellmath__30__13__out0({N271}), .inst_cellmath__30__13__in0(inst_cellmath__26), .inst_cellmath__30__13__in1(inst_cellmath__23), .inst_cellmath__30__13__in2(inst_cellmath__22));
cynw_cm_float_mul_inst_cellmath__30__14__bdw3636473930_bdw cynw_cm_float_mul_I17 (.inst_cellmath__30__14__out0({N272}), .inst_cellmath__30__14__in0(inst_cellmath__25), .inst_cellmath__30__14__in1(inst_cellmath__24), .inst_cellmath__30__14__in2(inst_cellmath__21));
cynw_cm_float_mul_inst_cellmath__30_0_bdw3636473930_bdw cynw_cm_float_mul_I18 (.inst_cellmath__30_0_out0(inst_cellmath__30), .inst_cellmath__30_0_in0({N272}), .inst_cellmath__30_0_in1({N271}));
cynw_cm_float_mul_inst_cellmath__34_0_bdw3636473930_bdw cynw_cm_float_mul_I19 (.inst_cellmath__34_0_out0({inst_cellmath__34[9], inst_cellmath__34[8], inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2], inst_cellmath__34[1], inst_cellmath__34[0]}), .inst_cellmath__34_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}), .inst_cellmath__34_0_in1({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_inst_cellmath__41__24__bdw3636473930_bdw cynw_cm_float_mul_I20 (.inst_cellmath__41__24__out0({N276}), .inst_cellmath__41__24__in0({inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2], inst_cellmath__34[1], inst_cellmath__34[0]}));
cynw_cm_float_mul_inst_cellmath__41__23__bdw3636473930_bdw cynw_cm_float_mul_I21 (.inst_cellmath__41__23__out0({N277}), .inst_cellmath__41__23__in0({N276}), .inst_cellmath__41__23__in1({inst_cellmath__34[8]}));
cynw_cm_float_mul_inst_cellmath__41_0_bdw3636473930_bdw cynw_cm_float_mul_I22 (.inst_cellmath__41_0_out0(inst_cellmath__41), .inst_cellmath__41_0_in0({N277}), .inst_cellmath__41_0_in1({inst_cellmath__34[9]}));
cynw_cm_float_mul_inst_cellmath__37_0_bdw3636473930_bdw cynw_cm_float_mul_I23 (.inst_cellmath__37_0_out0(inst_cellmath__37), .inst_cellmath__37_0_in0(inst_cellmath__41), .inst_cellmath__37_0_in1(inst_cellmath__30));
cynw_cm_float_mul_inst_cellmath__35__16__bdw3636473930_bdw cynw_cm_float_mul_I24 (.inst_cellmath__35__16__out0({N273}), .inst_cellmath__35__16__in0({inst_cellmath__34[9], inst_cellmath__34[8], inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2], inst_cellmath__34[1], inst_cellmath__34[0]}));
cynw_cm_float_mul_inst_cellmath__32__11__bdw3636473930_bdw cynw_cm_float_mul_I25 (.inst_cellmath__32__11__out0({N269}), .inst_cellmath__32__11__in0(inst_cellmath__25), .inst_cellmath__32__11__in1(inst_cellmath__24), .inst_cellmath__32__11__in2(inst_cellmath__22));
cynw_cm_float_mul_inst_cellmath__32__12__bdw3636473930_bdw cynw_cm_float_mul_I26 (.inst_cellmath__32__12__out0({N270}), .inst_cellmath__32__12__in0(inst_cellmath__26), .inst_cellmath__32__12__in1(inst_cellmath__23), .inst_cellmath__32__12__in2(inst_cellmath__21));
cynw_cm_float_mul_inst_cellmath__32_0_bdw3636473930_bdw cynw_cm_float_mul_I27 (.inst_cellmath__32_0_out0(inst_cellmath__32), .inst_cellmath__32_0_in0({N270}), .inst_cellmath__32_0_in1({N269}));
cynw_cm_float_mul_inst_cellmath__60_0_bdw3636473930_bdw cynw_cm_float_mul_I28 (.inst_cellmath__60_0_out0(inst_cellmath__60), .inst_cellmath__60_0_in0(inst_cellmath__37), .inst_cellmath__60_0_in1({N273}), .inst_cellmath__60_0_in2({inst_cellmath__34[9]}), .inst_cellmath__60_0_in3(inst_cellmath__32), .inst_cellmath__60_0_in4(inst_cellmath__29));
cynw_cm_float_mul_inst_cellmath__42__22__bdw3636473930_bdw cynw_cm_float_mul_I29 (.inst_cellmath__42__22__out0({N274}), .inst_cellmath__42__22__in0({inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2], inst_cellmath__34[1]}));
cynw_cm_float_mul_inst_cellmath__42__21__bdw3636473930_bdw cynw_cm_float_mul_I30 (.inst_cellmath__42__21__out0({N275}), .inst_cellmath__42__21__in0({N274}), .inst_cellmath__42__21__in1({inst_cellmath__34[8]}));
cynw_cm_float_mul_inst_cellmath__42_0_bdw3636473930_bdw cynw_cm_float_mul_I31 (.inst_cellmath__42_0_out0(inst_cellmath__42), .inst_cellmath__42_0_in0({N275}), .inst_cellmath__42_0_in1({inst_cellmath__34[9]}));
cynw_cm_float_mul_inst_cellmath__38_0_bdw3636473930_bdw cynw_cm_float_mul_I32 (.inst_cellmath__38_0_out0(inst_cellmath__38), .inst_cellmath__38_0_in0(inst_cellmath__42), .inst_cellmath__38_0_in1(inst_cellmath__30));
cynw_cm_float_mul_inst_cellmath__61_0_bdw3636473930_bdw cynw_cm_float_mul_I33 (.inst_cellmath__61_0_out0(inst_cellmath__61), .inst_cellmath__61_0_in0(inst_cellmath__38), .inst_cellmath__61_0_in1({inst_cellmath__34[9]}), .inst_cellmath__61_0_in2(inst_cellmath__32), .inst_cellmath__61_0_in3(inst_cellmath__29));
cynw_cm_float_mul_inst_cellmath__56_1_bdw3636473930_bdw cynw_cm_float_mul_I34 (.inst_cellmath__56_1_out0(inst_cellmath__56), .inst_cellmath__56_1_in0(inst_cellmath__61), .inst_cellmath__56_1_in1(inst_cellmath__60), .inst_cellmath__56_1_in2({inst_cellmath__43[47]}));
cynw_cm_float_mul_inst_cellmath__50_0_bdw3636473930_bdw cynw_cm_float_mul_I35 (.inst_cellmath__50_0_out0({inst_cellmath__50[7], inst_cellmath__50[6], inst_cellmath__50[5], inst_cellmath__50[4], inst_cellmath__50[3], inst_cellmath__50[2], inst_cellmath__50[1], inst_cellmath__50[0]}), .inst_cellmath__50_0_in0({inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2], inst_cellmath__34[1], inst_cellmath__34[0]}));
cynw_cm_float_mul_inst_cellmath__54_7_bdw3636473930_bdw cynw_cm_float_mul_I36 (.inst_cellmath__54_7_out0({inst_cellmath__54[7]}), .inst_cellmath__54_7_in0(inst_cellmath__38), .inst_cellmath__54_7_in1(inst_cellmath__37), .inst_cellmath__54_7_in2(inst_cellmath__29));
cynw_cm_float_mul_inst_cellmath__54__30__bdw3636473930_bdw cynw_cm_float_mul_I37 (.inst_cellmath__54__30__out0({N380}), .inst_cellmath__54__30__in0(inst_cellmath__38), .inst_cellmath__54__30__in1(inst_cellmath__37), .inst_cellmath__54__30__in2(inst_cellmath__29));
cynw_cm_float_mul_inst_cellmath__64_2WWMM_bdw3636473930_bdw cynw_cm_float_mul_I38 (.inst_cellmath__64_2WWMM_out0({x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__64_2WWMM_in0(inst_cellmath__56), .inst_cellmath__64_2WWMM_in1({N380}), .inst_cellmath__64_2WWMM_in2({inst_cellmath__54[7]}), .inst_cellmath__64_2WWMM_in3({inst_cellmath__50[7], inst_cellmath__50[6], inst_cellmath__50[5], inst_cellmath__50[4], inst_cellmath__50[3], inst_cellmath__50[2], inst_cellmath__50[1], inst_cellmath__50[0]}), .inst_cellmath__64_2WWMM_in4({inst_cellmath__43[47], inst_cellmath__43[46], inst_cellmath__43[45], inst_cellmath__43[44], inst_cellmath__43[43], inst_cellmath__43[42], inst_cellmath__43[41], inst_cellmath__43[40], inst_cellmath__43[39], inst_cellmath__43[38], inst_cellmath__43[37], inst_cellmath__43[36], inst_cellmath__43[35], inst_cellmath__43[34], inst_cellmath__43[33], inst_cellmath__43[32], inst_cellmath__43[31], inst_cellmath__43[30], inst_cellmath__43[29], inst_cellmath__43[28], inst_cellmath__43[27], inst_cellmath__43[26], inst_cellmath__43[25], inst_cellmath__43[24], inst_cellmath__43[23]}), .inst_cellmath__64_2WWMM_in5({inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2], inst_cellmath__34[1], inst_cellmath__34[0]}), .inst_cellmath__64_2WWMM_in6(inst_cellmath__29));
assign inst_cellmath__54[0] = 1'B0;
assign inst_cellmath__54[1] = 1'B0;
assign inst_cellmath__54[2] = 1'B0;
assign inst_cellmath__54[3] = 1'B0;
assign inst_cellmath__54[4] = 1'B0;
assign inst_cellmath__54[5] = 1'B0;
assign inst_cellmath__54[6] = 1'B0;
endmodule

module cynw_cm_float_mul_inst_cellmath__33_0_bdw3636473930_bdw (
	inst_cellmath__33_0_out0,
	inst_cellmath__33_0_in0,
	inst_cellmath__33_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__33_0_out0;
input  inst_cellmath__33_0_in0,
	inst_cellmath__33_0_in1;
XOR2XL inst_cellmath__33_0_I0 (.Y(inst_cellmath__33_0_out0), .A(inst_cellmath__33_0_in1), .B(inst_cellmath__33_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__26__8__bdw3636473930_bdw (
	inst_cellmath__26__8__out0,
	inst_cellmath__26__8__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__26__8__out0;
input [7:0] inst_cellmath__26__8__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__26__8__I0 (.Y(N11), .A(inst_cellmath__26__8__in0[0]), .B(inst_cellmath__26__8__in0[1]));
NOR2XL inst_cellmath__26__8__I1 (.Y(N12), .A(inst_cellmath__26__8__in0[7]), .B(inst_cellmath__26__8__in0[6]));
NOR2XL inst_cellmath__26__8__I2 (.Y(N13), .A(inst_cellmath__26__8__in0[5]), .B(inst_cellmath__26__8__in0[4]));
NOR2XL inst_cellmath__26__8__I3 (.Y(N14), .A(inst_cellmath__26__8__in0[3]), .B(inst_cellmath__26__8__in0[2]));
NAND2XL inst_cellmath__26__8__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__26__8__I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__26__8__I6 (.Y(inst_cellmath__26__8__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_inst_cellmath__17_0_bdw3636473930_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[0]), .B(inst_cellmath__17_0_in0[1]));
NAND2XL inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[6]));
NAND2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[5]), .B(inst_cellmath__17_0_in0[4]));
NAND2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[3]), .B(inst_cellmath__17_0_in0[2]));
NOR2XL inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_inst_cellmath__19__5__bdw3636473930_bdw (
	inst_cellmath__19__5__out0,
	inst_cellmath__19__5__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19__5__out0;
input [22:0] inst_cellmath__19__5__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__19__5__I1 (.Y(N27), .A(inst_cellmath__19__5__in0[22]), .B(inst_cellmath__19__5__in0[21]));
NOR2XL inst_cellmath__19__5__I2 (.Y(N28), .A(inst_cellmath__19__5__in0[20]), .B(inst_cellmath__19__5__in0[19]));
NOR2XL inst_cellmath__19__5__I3 (.Y(N29), .A(inst_cellmath__19__5__in0[18]), .B(inst_cellmath__19__5__in0[17]));
NOR2XL inst_cellmath__19__5__I4 (.Y(N30), .A(inst_cellmath__19__5__in0[16]), .B(inst_cellmath__19__5__in0[15]));
NOR2XL inst_cellmath__19__5__I5 (.Y(N31), .A(inst_cellmath__19__5__in0[14]), .B(inst_cellmath__19__5__in0[13]));
NOR2XL inst_cellmath__19__5__I6 (.Y(N32), .A(inst_cellmath__19__5__in0[12]), .B(inst_cellmath__19__5__in0[11]));
NOR2XL inst_cellmath__19__5__I7 (.Y(N33), .A(inst_cellmath__19__5__in0[10]), .B(inst_cellmath__19__5__in0[9]));
NOR2XL inst_cellmath__19__5__I8 (.Y(N34), .A(inst_cellmath__19__5__in0[8]), .B(inst_cellmath__19__5__in0[7]));
NOR2XL inst_cellmath__19__5__I9 (.Y(N35), .A(inst_cellmath__19__5__in0[6]), .B(inst_cellmath__19__5__in0[5]));
NOR2XL inst_cellmath__19__5__I10 (.Y(N36), .A(inst_cellmath__19__5__in0[4]), .B(inst_cellmath__19__5__in0[3]));
NAND2XL inst_cellmath__19__5__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__19__5__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__19__5__I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__19__5__I25 (.Y(N44), .A(inst_cellmath__19__5__in0[0]), .B(inst_cellmath__19__5__in0[1]), .C(inst_cellmath__19__5__in0[2]), .D(N39));
NOR2XL inst_cellmath__19__5__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__19__5__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__19__5__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__19__5__I23 (.Y(inst_cellmath__19__5__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_inst_cellmath__23_0_bdw3636473930_bdw (
	inst_cellmath__23_0_out0,
	inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__23_0_out0;
input  inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1;
AND2XL inst_cellmath__23_0_I0 (.Y(inst_cellmath__23_0_out0), .A(inst_cellmath__23_0_in1), .B(inst_cellmath__23_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__29__10__bdw3636473930_bdw (
	inst_cellmath__29__10__out0,
	inst_cellmath__29__10__in0,
	inst_cellmath__29__10__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__29__10__out0;
input  inst_cellmath__29__10__in0,
	inst_cellmath__29__10__in1;
AND2XL inst_cellmath__29__10__I0 (.Y(inst_cellmath__29__10__out0[0]), .A(inst_cellmath__29__10__in0), .B(inst_cellmath__29__10__in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__25__7__bdw3636473930_bdw (
	inst_cellmath__25__7__out0,
	inst_cellmath__25__7__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__25__7__out0;
input [7:0] inst_cellmath__25__7__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__25__7__I0 (.Y(N11), .A(inst_cellmath__25__7__in0[0]), .B(inst_cellmath__25__7__in0[1]));
NOR2XL inst_cellmath__25__7__I1 (.Y(N12), .A(inst_cellmath__25__7__in0[7]), .B(inst_cellmath__25__7__in0[6]));
NOR2XL inst_cellmath__25__7__I2 (.Y(N13), .A(inst_cellmath__25__7__in0[5]), .B(inst_cellmath__25__7__in0[4]));
NOR2XL inst_cellmath__25__7__I3 (.Y(N14), .A(inst_cellmath__25__7__in0[3]), .B(inst_cellmath__25__7__in0[2]));
NAND2XL inst_cellmath__25__7__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__25__7__I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__25__7__I6 (.Y(inst_cellmath__25__7__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_inst_cellmath__18_0_bdw3636473930_bdw (
	inst_cellmath__18_0_out0,
	inst_cellmath__18_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__18_0_out0;
input [7:0] inst_cellmath__18_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__18_0_I0 (.Y(N11), .A(inst_cellmath__18_0_in0[0]), .B(inst_cellmath__18_0_in0[1]));
NAND2XL inst_cellmath__18_0_I1 (.Y(N12), .A(inst_cellmath__18_0_in0[7]), .B(inst_cellmath__18_0_in0[6]));
NAND2XL inst_cellmath__18_0_I2 (.Y(N13), .A(inst_cellmath__18_0_in0[5]), .B(inst_cellmath__18_0_in0[4]));
NAND2XL inst_cellmath__18_0_I3 (.Y(N14), .A(inst_cellmath__18_0_in0[3]), .B(inst_cellmath__18_0_in0[2]));
NOR2XL inst_cellmath__18_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__18_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__18_0_I6 (.Y(inst_cellmath__18_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_inst_cellmath__20__6__bdw3636473930_bdw (
	inst_cellmath__20__6__out0,
	inst_cellmath__20__6__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__20__6__out0;
input [22:0] inst_cellmath__20__6__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__20__6__I1 (.Y(N27), .A(inst_cellmath__20__6__in0[22]), .B(inst_cellmath__20__6__in0[21]));
NOR2XL inst_cellmath__20__6__I2 (.Y(N28), .A(inst_cellmath__20__6__in0[20]), .B(inst_cellmath__20__6__in0[19]));
NOR2XL inst_cellmath__20__6__I3 (.Y(N29), .A(inst_cellmath__20__6__in0[18]), .B(inst_cellmath__20__6__in0[17]));
NOR2XL inst_cellmath__20__6__I4 (.Y(N30), .A(inst_cellmath__20__6__in0[16]), .B(inst_cellmath__20__6__in0[15]));
NOR2XL inst_cellmath__20__6__I5 (.Y(N31), .A(inst_cellmath__20__6__in0[14]), .B(inst_cellmath__20__6__in0[13]));
NOR2XL inst_cellmath__20__6__I6 (.Y(N32), .A(inst_cellmath__20__6__in0[12]), .B(inst_cellmath__20__6__in0[11]));
NOR2XL inst_cellmath__20__6__I7 (.Y(N33), .A(inst_cellmath__20__6__in0[10]), .B(inst_cellmath__20__6__in0[9]));
NOR2XL inst_cellmath__20__6__I8 (.Y(N34), .A(inst_cellmath__20__6__in0[8]), .B(inst_cellmath__20__6__in0[7]));
NOR2XL inst_cellmath__20__6__I9 (.Y(N35), .A(inst_cellmath__20__6__in0[6]), .B(inst_cellmath__20__6__in0[5]));
NOR2XL inst_cellmath__20__6__I10 (.Y(N36), .A(inst_cellmath__20__6__in0[4]), .B(inst_cellmath__20__6__in0[3]));
NAND2XL inst_cellmath__20__6__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__20__6__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__20__6__I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__20__6__I25 (.Y(N44), .A(inst_cellmath__20__6__in0[0]), .B(inst_cellmath__20__6__in0[1]), .C(inst_cellmath__20__6__in0[2]), .D(N39));
NOR2XL inst_cellmath__20__6__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__20__6__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__20__6__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__20__6__I23 (.Y(inst_cellmath__20__6__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_inst_cellmath__24_0_bdw3636473930_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__24_0_out0;
input  inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1;
AND2XL inst_cellmath__24_0_I0 (.Y(inst_cellmath__24_0_out0), .A(inst_cellmath__24_0_in1), .B(inst_cellmath__24_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__29__9__bdw3636473930_bdw (
	inst_cellmath__29__9__out0,
	inst_cellmath__29__9__in0,
	inst_cellmath__29__9__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__29__9__out0;
input  inst_cellmath__29__9__in0,
	inst_cellmath__29__9__in1;
AND2XL inst_cellmath__29__9__I0 (.Y(inst_cellmath__29__9__out0[0]), .A(inst_cellmath__29__9__in0), .B(inst_cellmath__29__9__in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__21_0_bdw3636473930_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__21_0_out0;
input  inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1;
NOR2BX1 inst_cellmath__21_0_I2 (.Y(inst_cellmath__21_0_out0), .AN(inst_cellmath__21_0_in1), .B(inst_cellmath__21_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__22_0_bdw3636473930_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__22_0_out0;
input  inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1;
NOR2BX1 inst_cellmath__22_0_I2 (.Y(inst_cellmath__22_0_out0), .AN(inst_cellmath__22_0_in1), .B(inst_cellmath__22_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__29_0_bdw3636473930_bdw (
	inst_cellmath__29_0_out0,
	inst_cellmath__29_0_in0,
	inst_cellmath__29_0_in1,
	inst_cellmath__29_0_in2,
	inst_cellmath__29_0_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__29_0_out0;
input [0:0] inst_cellmath__29_0_in0,
	inst_cellmath__29_0_in1;
input  inst_cellmath__29_0_in2,
	inst_cellmath__29_0_in3;
OR4X1 inst_cellmath__29_0_I6 (.Y(inst_cellmath__29_0_out0), .A(inst_cellmath__29_0_in2), .B(inst_cellmath__29_0_in3), .C(inst_cellmath__29_0_in1[0]), .D(inst_cellmath__29_0_in0[0]));
endmodule

module cynw_cm_float_mul_inst_cellmath__53_0_bdw3636473930_bdw (
	inst_cellmath__53_0_out0,
	inst_cellmath__53_0_in0,
	inst_cellmath__53_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__53_0_out0;
input  inst_cellmath__53_0_in0,
	inst_cellmath__53_0_in1;
NOR2BX1 inst_cellmath__53_0_I2 (.Y(inst_cellmath__53_0_out0), .AN(inst_cellmath__53_0_in0), .B(inst_cellmath__53_0_in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__43_0_bdw3636473930_bdw (
	inst_cellmath__43_0_out0,
	inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__43_0_out0;
input [22:0] inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1;
wire N383,N385,N387,N389,N391,N393,N395 
	,N397,N399,N401,N403,N405,N407,N409,N411 
	,N413,N415,N417,N419,N421,N423,N425,N427 
	,N440,N442,N444,N446,N448,N450,N452,N454 
	,N456,N458,N460,N462,N464,N466,N468,N470 
	,N472,N474,N476,N478,N480,N482,N484,N486 
	,N499,N501,N503,N505,N507,N509,N511,N513 
	,N515,N517,N519,N521,N523,N525,N527,N529 
	,N531,N533,N535,N537,N539,N541,N543,N545 
	,N558,N560,N562,N564,N566,N568,N570,N572 
	,N574,N576,N578,N580,N582,N584,N586,N588 
	,N590,N592,N594,N596,N598,N600,N602,N604 
	,N617,N619,N621,N623,N625,N627,N629,N631 
	,N633,N635,N637,N639,N641,N643,N645,N647 
	,N649,N651,N653,N655,N657,N659,N661,N663 
	,N676,N678,N680,N682,N684,N686,N688,N690 
	,N692,N694,N696,N698,N700,N702,N704,N706 
	,N708,N710,N712,N714,N716,N718,N720,N722 
	,N735,N737,N739,N741,N743,N745,N747,N749 
	,N751,N753,N755,N757,N759,N761,N763,N765 
	,N767,N769,N771,N773,N775,N777,N779,N781 
	,N794,N796,N798,N800,N802,N804,N806,N808 
	,N810,N812,N814,N816,N818,N820,N822,N824 
	,N826,N828,N830,N832,N834,N836,N838,N840 
	,N853,N855,N857,N859,N861,N863,N865,N867 
	,N869,N871,N873,N875,N877,N879,N881,N883 
	,N885,N887,N889,N891,N893,N895,N897,N899 
	,N912,N914,N916,N918,N920,N922,N924,N926 
	,N928,N930,N932,N934,N936,N938,N940,N942 
	,N944,N946,N948,N950,N952,N954,N956,N958 
	,N971,N973,N975,N977,N979,N981,N983,N985 
	,N987,N989,N991,N993,N995,N997,N999,N1001 
	,N1003,N1005,N1007,N1009,N1011,N1013,N1015,N1017 
	,N1030,N1032,N1034,N1036,N1038,N1040,N1042,N1044 
	,N1046,N1048,N1050,N1052,N1054,N1056,N1058,N1060 
	,N1062,N1064,N1066,N1068,N1070,N1072,N1074,N1076 
	,N1089,N1091,N1093,N1095,N1097,N1099,N1101,N1103 
	,N1105,N1107,N1109,N1111,N1113,N1115,N1117,N1119 
	,N1121,N1123,N1125,N1127,N1129,N1131,N1133,N1135 
	,N1148,N1150,N1152,N1154,N1156,N1158,N1160,N1162 
	,N1164,N1166,N1168,N1170,N1172,N1174,N1176,N1178 
	,N1180,N1182,N1184,N1186,N1188,N1190,N1192,N1194 
	,N1207,N1209,N1211,N1213,N1215,N1217,N1219,N1221 
	,N1223,N1225,N1227,N1229,N1231,N1233,N1235,N1237 
	,N1239,N1241,N1243,N1245,N1247,N1249,N1251,N1253 
	,N1266,N1268,N1270,N1272,N1274,N1276,N1278,N1280 
	,N1282,N1284,N1286,N1288,N1290,N1292,N1294,N1296 
	,N1298,N1300,N1302,N1304,N1306,N1308,N1310,N1312 
	,N1325,N1327,N1329,N1331,N1333,N1335,N1337,N1339 
	,N1341,N1343,N1345,N1347,N1349,N1351,N1353,N1355 
	,N1357,N1359,N1361,N1363,N1365,N1367,N1369,N1371 
	,N1384,N1386,N1388,N1390,N1392,N1394,N1396,N1398 
	,N1400,N1402,N1404,N1406,N1408,N1410,N1412,N1414 
	,N1416,N1418,N1420,N1422,N1424,N1426,N1428,N1430 
	,N1443,N1445,N1447,N1449,N1451,N1453,N1455,N1457 
	,N1459,N1461,N1463,N1465,N1467,N1469,N1471,N1473 
	,N1475,N1477,N1479,N1481,N1483,N1485,N1487,N1489 
	,N1502,N1504,N1506,N1508,N1510,N1512,N1514,N1516 
	,N1518,N1520,N1522,N1524,N1526,N1528,N1530,N1532 
	,N1534,N1536,N1538,N1540,N1542,N1544,N1546,N1548 
	,N1561,N1563,N1565,N1567,N1569,N1571,N1573,N1575 
	,N1577,N1579,N1581,N1583,N1585,N1587,N1589,N1591 
	,N1593,N1595,N1597,N1599,N1601,N1603,N1605,N1607 
	,N1620,N1622,N1624,N1626,N1628,N1630,N1632,N1634 
	,N1636,N1638,N1640,N1642,N1644,N1646,N1648,N1650 
	,N1652,N1654,N1656,N1658,N1660,N1662,N1664,N1666 
	,N1679,N1681,N1683,N1685,N1687,N1689,N1691,N1693 
	,N1695,N1697,N1699,N1701,N1703,N1705,N1707,N1709 
	,N1711,N1713,N1715,N1717,N1719,N1721,N1723,N1725 
	,N1734,N1736,N1738,N1740,N1742,N1744,N1746,N1748 
	,N1750,N1752,N1754,N1756,N1758,N1760,N1762,N1764 
	,N1766,N1768,N1770,N1772,N1774,N1776,N1778,N1812 
	,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820 
	,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828 
	,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836 
	,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844 
	,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852 
	,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860 
	,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868 
	,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876 
	,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884 
	,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892 
	,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900 
	,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908 
	,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916 
	,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924 
	,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932 
	,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940 
	,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948 
	,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956 
	,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964 
	,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972 
	,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980 
	,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988 
	,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996 
	,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004 
	,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012 
	,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020 
	,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028 
	,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036 
	,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044 
	,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052 
	,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060 
	,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068 
	,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076 
	,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084 
	,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092 
	,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100 
	,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108 
	,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116 
	,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124 
	,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132 
	,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140 
	,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148 
	,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156 
	,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164 
	,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172 
	,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180 
	,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188 
	,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196 
	,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204 
	,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212 
	,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220 
	,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228 
	,N2229,N2230,N2231,N2232,N2233,N2236,N2237,N2238 
	,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246 
	,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254 
	,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262 
	,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270 
	,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278 
	,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286 
	,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294 
	,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302 
	,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310 
	,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318 
	,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326 
	,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334 
	,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342 
	,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350 
	,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358 
	,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366 
	,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374 
	,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382 
	,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390 
	,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398 
	,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406 
	,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414 
	,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422 
	,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430 
	,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438 
	,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446 
	,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454 
	,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462 
	,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470 
	,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478 
	,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486 
	,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494 
	,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502 
	,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510 
	,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518 
	,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526 
	,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534 
	,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542 
	,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550 
	,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558 
	,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566 
	,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574 
	,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582 
	,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590 
	,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598 
	,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606 
	,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614 
	,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622 
	,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630 
	,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638 
	,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646 
	,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654 
	,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662 
	,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670 
	,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678 
	,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686 
	,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694 
	,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702 
	,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710 
	,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718 
	,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726 
	,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734 
	,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742 
	,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750 
	,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758 
	,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766 
	,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774 
	,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782 
	,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790 
	,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798 
	,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806 
	,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814 
	,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822 
	,N2823,N2824,N2826,N2827,N2828,N2829,N2830,N2831 
	,N2832,N2833,N2835,N2836,N2837,N2838,N2839,N2840 
	,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848 
	,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856 
	,N2859,N2867,N2875,N2887,N2899,N2915,N2931,N2935 
	,N2936,N2955,N2959,N2985,N2987,N2991,N2992,N3019 
	,N3057,N3059,N3082,N3085,N3088,N3091,N3094,N3097 
	,N3100,N3103,N3106,N3109,N3112,N3115,N3118,N3121 
	,N3124,N3141,N3143,N3144,N3145,N3146,N3147,N3148 
	,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156 
	,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164 
	,N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172 
	,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180 
	,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188 
	,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196 
	,N3197,N3198,N3199,N3200,N3202,N3204,N3205,N3206 
	,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214 
	,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222 
	,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230 
	,N3232,N3234,N3235,N3236,N3237,N3238,N3239,N3240 
	,N3241,N3242,N3243,N3246,N3248,N3249,N3250,N3252 
	,N3255,N3256,N3258,N3259,N3260,N3264,N3269,N3270 
	,N3272,N3273,N3274,N3278,N3282,N3283,N3284,N3288 
	,N3292,N3296,N3297,N3298,N3303,N3304,N3306,N3307 
	,N3308,N3312,N3316,N3317,N3318,N3322,N3326,N3330 
	,N3331,N3332,N3336,N3337,N3338,N3342,N3346,N3350 
	,N3354,N3358,N3359,N3360,N3364,N3365,N3366,N3370 
	,N3371,N3372,N3376,N3585,N3586,N3587,N3588,N3589 
	,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597 
	,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605 
	,N3606,N3607,N3608,N3609,N3615,N3616,N3617,N3618 
	,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626 
	,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634 
	,N3635,N3636,N3639,N3640,N3646,N3657,N3658,N3690 
	,N3724,N3734,N3738,N3742,N3743,N3744,N3745,N3746 
	,N3747,N3748,N3749,N3757,N3764;
INVXL inst_cellmath__43_0_I1991 (.Y(N3585), .A(inst_cellmath__43_0_in0[0]));
INVXL inst_cellmath__43_0_I1992 (.Y(N3586), .A(inst_cellmath__43_0_in0[1]));
INVXL inst_cellmath__43_0_I1993 (.Y(N3587), .A(inst_cellmath__43_0_in0[2]));
INVXL inst_cellmath__43_0_I1994 (.Y(N3588), .A(inst_cellmath__43_0_in0[3]));
INVXL inst_cellmath__43_0_I1995 (.Y(N3589), .A(inst_cellmath__43_0_in0[4]));
INVXL inst_cellmath__43_0_I1996 (.Y(N3590), .A(inst_cellmath__43_0_in0[5]));
INVXL inst_cellmath__43_0_I1997 (.Y(N3591), .A(inst_cellmath__43_0_in0[6]));
INVXL inst_cellmath__43_0_I1998 (.Y(N3592), .A(inst_cellmath__43_0_in0[7]));
INVXL inst_cellmath__43_0_I1999 (.Y(N3593), .A(inst_cellmath__43_0_in0[8]));
INVXL inst_cellmath__43_0_I2000 (.Y(N3594), .A(inst_cellmath__43_0_in0[9]));
INVXL inst_cellmath__43_0_I2001 (.Y(N3595), .A(inst_cellmath__43_0_in0[10]));
INVXL inst_cellmath__43_0_I2002 (.Y(N3596), .A(inst_cellmath__43_0_in0[11]));
INVXL inst_cellmath__43_0_I2003 (.Y(N3597), .A(inst_cellmath__43_0_in0[12]));
INVXL inst_cellmath__43_0_I2004 (.Y(N3598), .A(inst_cellmath__43_0_in0[13]));
INVXL inst_cellmath__43_0_I2005 (.Y(N3599), .A(inst_cellmath__43_0_in0[14]));
INVXL inst_cellmath__43_0_I2006 (.Y(N3600), .A(inst_cellmath__43_0_in0[15]));
INVXL inst_cellmath__43_0_I2007 (.Y(N3601), .A(inst_cellmath__43_0_in0[16]));
INVXL inst_cellmath__43_0_I2008 (.Y(N3602), .A(inst_cellmath__43_0_in0[17]));
INVXL inst_cellmath__43_0_I2009 (.Y(N3603), .A(inst_cellmath__43_0_in0[18]));
INVXL inst_cellmath__43_0_I2010 (.Y(N3604), .A(inst_cellmath__43_0_in0[19]));
INVXL inst_cellmath__43_0_I2011 (.Y(N3605), .A(inst_cellmath__43_0_in0[20]));
INVXL inst_cellmath__43_0_I2012 (.Y(N3606), .A(inst_cellmath__43_0_in0[21]));
INVXL inst_cellmath__43_0_I2013 (.Y(N3607), .A(inst_cellmath__43_0_in0[22]));
INVXL inst_cellmath__43_0_I2014 (.Y(N3608), .A(inst_cellmath__43_0_in1[0]));
NOR2XL inst_cellmath__43_0_I87 (.Y(inst_cellmath__43_0_out0[0]), .A(N3608), .B(N3585));
NOR2XL inst_cellmath__43_0_I88 (.Y(N383), .A(N3608), .B(N3586));
NOR2XL inst_cellmath__43_0_I89 (.Y(N385), .A(N3608), .B(N3587));
NOR2XL inst_cellmath__43_0_I90 (.Y(N387), .A(N3608), .B(N3588));
NOR2XL inst_cellmath__43_0_I91 (.Y(N389), .A(N3608), .B(N3589));
NOR2XL inst_cellmath__43_0_I92 (.Y(N391), .A(N3608), .B(N3590));
NOR2XL inst_cellmath__43_0_I93 (.Y(N393), .A(N3608), .B(N3591));
NOR2XL inst_cellmath__43_0_I94 (.Y(N395), .A(N3608), .B(N3592));
NOR2XL inst_cellmath__43_0_I95 (.Y(N397), .A(N3608), .B(N3593));
NOR2XL inst_cellmath__43_0_I96 (.Y(N399), .A(N3608), .B(N3594));
NOR2XL inst_cellmath__43_0_I97 (.Y(N401), .A(N3608), .B(N3595));
NOR2XL inst_cellmath__43_0_I98 (.Y(N403), .A(N3608), .B(N3596));
NOR2XL inst_cellmath__43_0_I99 (.Y(N405), .A(N3608), .B(N3597));
NOR2XL inst_cellmath__43_0_I100 (.Y(N407), .A(N3608), .B(N3598));
NOR2XL inst_cellmath__43_0_I101 (.Y(N409), .A(N3608), .B(N3599));
NOR2XL inst_cellmath__43_0_I102 (.Y(N411), .A(N3608), .B(N3600));
NOR2XL inst_cellmath__43_0_I103 (.Y(N413), .A(N3608), .B(N3601));
NOR2XL inst_cellmath__43_0_I104 (.Y(N415), .A(N3608), .B(N3602));
NOR2XL inst_cellmath__43_0_I105 (.Y(N417), .A(N3608), .B(N3603));
NOR2XL inst_cellmath__43_0_I106 (.Y(N419), .A(N3608), .B(N3604));
NOR2XL inst_cellmath__43_0_I107 (.Y(N421), .A(N3608), .B(N3605));
NOR2XL inst_cellmath__43_0_I108 (.Y(N423), .A(N3608), .B(N3606));
NOR2XL inst_cellmath__43_0_I109 (.Y(N425), .A(N3608), .B(N3607));
INVXL inst_cellmath__43_0_I110 (.Y(N427), .A(N3608));
INVXL inst_cellmath__43_0_I2015 (.Y(N3609), .A(inst_cellmath__43_0_in1[1]));
NOR2XL inst_cellmath__43_0_I116 (.Y(N440), .A(N3609), .B(N3585));
NOR2XL inst_cellmath__43_0_I117 (.Y(N442), .A(N3609), .B(N3586));
NOR2XL inst_cellmath__43_0_I118 (.Y(N444), .A(N3609), .B(N3587));
NOR2XL inst_cellmath__43_0_I119 (.Y(N446), .A(N3609), .B(N3588));
NOR2XL inst_cellmath__43_0_I120 (.Y(N448), .A(N3609), .B(N3589));
NOR2XL inst_cellmath__43_0_I121 (.Y(N450), .A(N3609), .B(N3590));
NOR2XL inst_cellmath__43_0_I122 (.Y(N452), .A(N3609), .B(N3591));
NOR2XL inst_cellmath__43_0_I123 (.Y(N454), .A(N3609), .B(N3592));
NOR2XL inst_cellmath__43_0_I124 (.Y(N456), .A(N3609), .B(N3593));
NOR2XL inst_cellmath__43_0_I125 (.Y(N458), .A(N3609), .B(N3594));
NOR2XL inst_cellmath__43_0_I126 (.Y(N460), .A(N3609), .B(N3595));
NOR2XL inst_cellmath__43_0_I127 (.Y(N462), .A(N3609), .B(N3596));
NOR2XL inst_cellmath__43_0_I128 (.Y(N464), .A(N3609), .B(N3597));
NOR2XL inst_cellmath__43_0_I129 (.Y(N466), .A(N3609), .B(N3598));
NOR2XL inst_cellmath__43_0_I130 (.Y(N468), .A(N3609), .B(N3599));
NOR2XL inst_cellmath__43_0_I131 (.Y(N470), .A(N3609), .B(N3600));
NOR2XL inst_cellmath__43_0_I132 (.Y(N472), .A(N3609), .B(N3601));
NOR2XL inst_cellmath__43_0_I133 (.Y(N474), .A(N3609), .B(N3602));
NOR2XL inst_cellmath__43_0_I134 (.Y(N476), .A(N3609), .B(N3603));
NOR2XL inst_cellmath__43_0_I135 (.Y(N478), .A(N3609), .B(N3604));
NOR2XL inst_cellmath__43_0_I136 (.Y(N480), .A(N3609), .B(N3605));
NOR2XL inst_cellmath__43_0_I137 (.Y(N482), .A(N3609), .B(N3606));
NOR2XL inst_cellmath__43_0_I138 (.Y(N484), .A(N3609), .B(N3607));
INVXL inst_cellmath__43_0_I139 (.Y(N486), .A(N3609));
INVXL inst_cellmath__43_0_I2163 (.Y(N3615), .A(inst_cellmath__43_0_in1[2]));
NOR2XL inst_cellmath__43_0_I145 (.Y(N499), .A(N3615), .B(N3585));
NOR2XL inst_cellmath__43_0_I146 (.Y(N501), .A(N3615), .B(N3586));
NOR2XL inst_cellmath__43_0_I147 (.Y(N503), .A(N3615), .B(N3587));
NOR2XL inst_cellmath__43_0_I148 (.Y(N505), .A(N3615), .B(N3588));
NOR2XL inst_cellmath__43_0_I149 (.Y(N507), .A(N3615), .B(N3589));
NOR2XL inst_cellmath__43_0_I150 (.Y(N509), .A(N3615), .B(N3590));
NOR2XL inst_cellmath__43_0_I151 (.Y(N511), .A(N3615), .B(N3591));
NOR2XL inst_cellmath__43_0_I152 (.Y(N513), .A(N3615), .B(N3592));
NOR2XL inst_cellmath__43_0_I153 (.Y(N515), .A(N3615), .B(N3593));
NOR2XL inst_cellmath__43_0_I154 (.Y(N517), .A(N3615), .B(N3594));
NOR2XL inst_cellmath__43_0_I155 (.Y(N519), .A(N3615), .B(N3595));
NOR2XL inst_cellmath__43_0_I156 (.Y(N521), .A(N3615), .B(N3596));
NOR2XL inst_cellmath__43_0_I157 (.Y(N523), .A(N3615), .B(N3597));
NOR2XL inst_cellmath__43_0_I158 (.Y(N525), .A(N3615), .B(N3598));
NOR2XL inst_cellmath__43_0_I159 (.Y(N527), .A(N3615), .B(N3599));
NOR2XL inst_cellmath__43_0_I160 (.Y(N529), .A(N3615), .B(N3600));
NOR2XL inst_cellmath__43_0_I161 (.Y(N531), .A(N3615), .B(N3601));
NOR2XL inst_cellmath__43_0_I162 (.Y(N533), .A(N3615), .B(N3602));
NOR2XL inst_cellmath__43_0_I163 (.Y(N535), .A(N3615), .B(N3603));
NOR2XL inst_cellmath__43_0_I164 (.Y(N537), .A(N3615), .B(N3604));
NOR2XL inst_cellmath__43_0_I165 (.Y(N539), .A(N3615), .B(N3605));
NOR2XL inst_cellmath__43_0_I166 (.Y(N541), .A(N3615), .B(N3606));
NOR2XL inst_cellmath__43_0_I167 (.Y(N543), .A(N3615), .B(N3607));
INVXL inst_cellmath__43_0_I168 (.Y(N545), .A(N3615));
INVXL inst_cellmath__43_0_I2022 (.Y(N3616), .A(inst_cellmath__43_0_in1[3]));
NOR2XL inst_cellmath__43_0_I174 (.Y(N558), .A(N3616), .B(N3585));
NOR2XL inst_cellmath__43_0_I175 (.Y(N560), .A(N3616), .B(N3586));
NOR2XL inst_cellmath__43_0_I176 (.Y(N562), .A(N3616), .B(N3587));
NOR2XL inst_cellmath__43_0_I177 (.Y(N564), .A(N3616), .B(N3588));
NOR2XL inst_cellmath__43_0_I178 (.Y(N566), .A(N3616), .B(N3589));
NOR2XL inst_cellmath__43_0_I179 (.Y(N568), .A(N3616), .B(N3590));
NOR2XL inst_cellmath__43_0_I180 (.Y(N570), .A(N3616), .B(N3591));
NOR2XL inst_cellmath__43_0_I181 (.Y(N572), .A(N3616), .B(N3592));
NOR2XL inst_cellmath__43_0_I182 (.Y(N574), .A(N3616), .B(N3593));
NOR2XL inst_cellmath__43_0_I183 (.Y(N576), .A(N3616), .B(N3594));
NOR2XL inst_cellmath__43_0_I184 (.Y(N578), .A(N3616), .B(N3595));
NOR2XL inst_cellmath__43_0_I185 (.Y(N580), .A(N3616), .B(N3596));
NOR2XL inst_cellmath__43_0_I186 (.Y(N582), .A(N3616), .B(N3597));
NOR2XL inst_cellmath__43_0_I187 (.Y(N584), .A(N3616), .B(N3598));
NOR2XL inst_cellmath__43_0_I188 (.Y(N586), .A(N3616), .B(N3599));
NOR2XL inst_cellmath__43_0_I189 (.Y(N588), .A(N3616), .B(N3600));
NOR2XL inst_cellmath__43_0_I190 (.Y(N590), .A(N3616), .B(N3601));
NOR2XL inst_cellmath__43_0_I191 (.Y(N592), .A(N3616), .B(N3602));
NOR2XL inst_cellmath__43_0_I192 (.Y(N594), .A(N3616), .B(N3603));
NOR2XL inst_cellmath__43_0_I193 (.Y(N596), .A(N3616), .B(N3604));
NOR2XL inst_cellmath__43_0_I194 (.Y(N598), .A(N3616), .B(N3605));
NOR2XL inst_cellmath__43_0_I195 (.Y(N600), .A(N3616), .B(N3606));
NOR2XL inst_cellmath__43_0_I196 (.Y(N602), .A(N3616), .B(N3607));
INVXL inst_cellmath__43_0_I197 (.Y(N604), .A(N3616));
INVXL inst_cellmath__43_0_I2023 (.Y(N3617), .A(inst_cellmath__43_0_in1[4]));
NOR2XL inst_cellmath__43_0_I203 (.Y(N617), .A(N3617), .B(N3585));
NOR2XL inst_cellmath__43_0_I204 (.Y(N619), .A(N3617), .B(N3586));
NOR2XL inst_cellmath__43_0_I205 (.Y(N621), .A(N3617), .B(N3587));
NOR2XL inst_cellmath__43_0_I206 (.Y(N623), .A(N3617), .B(N3588));
NOR2XL inst_cellmath__43_0_I207 (.Y(N625), .A(N3617), .B(N3589));
NOR2XL inst_cellmath__43_0_I208 (.Y(N627), .A(N3617), .B(N3590));
NOR2XL inst_cellmath__43_0_I209 (.Y(N629), .A(N3617), .B(N3591));
NOR2XL inst_cellmath__43_0_I210 (.Y(N631), .A(N3617), .B(N3592));
NOR2XL inst_cellmath__43_0_I211 (.Y(N633), .A(N3617), .B(N3593));
NOR2XL inst_cellmath__43_0_I212 (.Y(N635), .A(N3617), .B(N3594));
NOR2XL inst_cellmath__43_0_I213 (.Y(N637), .A(N3617), .B(N3595));
NOR2XL inst_cellmath__43_0_I214 (.Y(N639), .A(N3617), .B(N3596));
NOR2XL inst_cellmath__43_0_I215 (.Y(N641), .A(N3617), .B(N3597));
NOR2XL inst_cellmath__43_0_I216 (.Y(N643), .A(N3617), .B(N3598));
NOR2XL inst_cellmath__43_0_I217 (.Y(N645), .A(N3617), .B(N3599));
NOR2XL inst_cellmath__43_0_I218 (.Y(N647), .A(N3617), .B(N3600));
NOR2XL inst_cellmath__43_0_I219 (.Y(N649), .A(N3617), .B(N3601));
NOR2XL inst_cellmath__43_0_I220 (.Y(N651), .A(N3617), .B(N3602));
NOR2XL inst_cellmath__43_0_I221 (.Y(N653), .A(N3617), .B(N3603));
NOR2XL inst_cellmath__43_0_I222 (.Y(N655), .A(N3617), .B(N3604));
NOR2XL inst_cellmath__43_0_I223 (.Y(N657), .A(N3617), .B(N3605));
NOR2XL inst_cellmath__43_0_I224 (.Y(N659), .A(N3617), .B(N3606));
NOR2XL inst_cellmath__43_0_I225 (.Y(N661), .A(N3617), .B(N3607));
INVXL inst_cellmath__43_0_I226 (.Y(N663), .A(N3617));
INVXL inst_cellmath__43_0_I2024 (.Y(N3618), .A(inst_cellmath__43_0_in1[5]));
NOR2XL inst_cellmath__43_0_I232 (.Y(N676), .A(N3618), .B(N3585));
NOR2XL inst_cellmath__43_0_I233 (.Y(N678), .A(N3618), .B(N3586));
NOR2XL inst_cellmath__43_0_I234 (.Y(N680), .A(N3618), .B(N3587));
NOR2XL inst_cellmath__43_0_I235 (.Y(N682), .A(N3618), .B(N3588));
NOR2XL inst_cellmath__43_0_I236 (.Y(N684), .A(N3618), .B(N3589));
NOR2XL inst_cellmath__43_0_I237 (.Y(N686), .A(N3618), .B(N3590));
NOR2XL inst_cellmath__43_0_I238 (.Y(N688), .A(N3618), .B(N3591));
NOR2XL inst_cellmath__43_0_I239 (.Y(N690), .A(N3618), .B(N3592));
NOR2XL inst_cellmath__43_0_I240 (.Y(N692), .A(N3618), .B(N3593));
NOR2XL inst_cellmath__43_0_I241 (.Y(N694), .A(N3618), .B(N3594));
NOR2XL inst_cellmath__43_0_I242 (.Y(N696), .A(N3618), .B(N3595));
NOR2XL inst_cellmath__43_0_I243 (.Y(N698), .A(N3618), .B(N3596));
NOR2XL inst_cellmath__43_0_I244 (.Y(N700), .A(N3618), .B(N3597));
NOR2XL inst_cellmath__43_0_I245 (.Y(N702), .A(N3618), .B(N3598));
NOR2XL inst_cellmath__43_0_I246 (.Y(N704), .A(N3618), .B(N3599));
NOR2XL inst_cellmath__43_0_I247 (.Y(N706), .A(N3618), .B(N3600));
NOR2XL inst_cellmath__43_0_I248 (.Y(N708), .A(N3618), .B(N3601));
NOR2XL inst_cellmath__43_0_I249 (.Y(N710), .A(N3618), .B(N3602));
NOR2XL inst_cellmath__43_0_I250 (.Y(N712), .A(N3618), .B(N3603));
NOR2XL inst_cellmath__43_0_I251 (.Y(N714), .A(N3618), .B(N3604));
NOR2XL inst_cellmath__43_0_I252 (.Y(N716), .A(N3618), .B(N3605));
NOR2XL inst_cellmath__43_0_I253 (.Y(N718), .A(N3618), .B(N3606));
NOR2XL inst_cellmath__43_0_I254 (.Y(N720), .A(N3618), .B(N3607));
INVXL inst_cellmath__43_0_I255 (.Y(N722), .A(N3618));
INVXL inst_cellmath__43_0_I2025 (.Y(N3619), .A(inst_cellmath__43_0_in1[6]));
NOR2XL inst_cellmath__43_0_I261 (.Y(N735), .A(N3619), .B(N3585));
NOR2XL inst_cellmath__43_0_I262 (.Y(N737), .A(N3619), .B(N3586));
NOR2XL inst_cellmath__43_0_I263 (.Y(N739), .A(N3619), .B(N3587));
NOR2XL inst_cellmath__43_0_I264 (.Y(N741), .A(N3619), .B(N3588));
NOR2XL inst_cellmath__43_0_I265 (.Y(N743), .A(N3619), .B(N3589));
NOR2XL inst_cellmath__43_0_I266 (.Y(N745), .A(N3619), .B(N3590));
NOR2XL inst_cellmath__43_0_I267 (.Y(N747), .A(N3619), .B(N3591));
NOR2XL inst_cellmath__43_0_I268 (.Y(N749), .A(N3619), .B(N3592));
NOR2XL inst_cellmath__43_0_I269 (.Y(N751), .A(N3619), .B(N3593));
NOR2XL inst_cellmath__43_0_I270 (.Y(N753), .A(N3619), .B(N3594));
NOR2XL inst_cellmath__43_0_I271 (.Y(N755), .A(N3619), .B(N3595));
NOR2XL inst_cellmath__43_0_I272 (.Y(N757), .A(N3619), .B(N3596));
NOR2XL inst_cellmath__43_0_I273 (.Y(N759), .A(N3619), .B(N3597));
NOR2XL inst_cellmath__43_0_I274 (.Y(N761), .A(N3619), .B(N3598));
NOR2XL inst_cellmath__43_0_I275 (.Y(N763), .A(N3619), .B(N3599));
NOR2XL inst_cellmath__43_0_I276 (.Y(N765), .A(N3619), .B(N3600));
NOR2XL inst_cellmath__43_0_I277 (.Y(N767), .A(N3619), .B(N3601));
NOR2XL inst_cellmath__43_0_I278 (.Y(N769), .A(N3619), .B(N3602));
NOR2XL inst_cellmath__43_0_I279 (.Y(N771), .A(N3619), .B(N3603));
NOR2XL inst_cellmath__43_0_I280 (.Y(N773), .A(N3619), .B(N3604));
NOR2XL inst_cellmath__43_0_I281 (.Y(N775), .A(N3619), .B(N3605));
NOR2XL inst_cellmath__43_0_I282 (.Y(N777), .A(N3619), .B(N3606));
NOR2XL inst_cellmath__43_0_I283 (.Y(N779), .A(N3619), .B(N3607));
INVXL inst_cellmath__43_0_I284 (.Y(N781), .A(N3619));
INVXL inst_cellmath__43_0_I2026 (.Y(N3620), .A(inst_cellmath__43_0_in1[7]));
NOR2XL inst_cellmath__43_0_I290 (.Y(N794), .A(N3620), .B(N3585));
NOR2XL inst_cellmath__43_0_I291 (.Y(N796), .A(N3620), .B(N3586));
NOR2XL inst_cellmath__43_0_I292 (.Y(N798), .A(N3620), .B(N3587));
NOR2XL inst_cellmath__43_0_I293 (.Y(N800), .A(N3620), .B(N3588));
NOR2XL inst_cellmath__43_0_I294 (.Y(N802), .A(N3620), .B(N3589));
NOR2XL inst_cellmath__43_0_I295 (.Y(N804), .A(N3620), .B(N3590));
NOR2XL inst_cellmath__43_0_I296 (.Y(N806), .A(N3620), .B(N3591));
NOR2XL inst_cellmath__43_0_I297 (.Y(N808), .A(N3620), .B(N3592));
NOR2XL inst_cellmath__43_0_I298 (.Y(N810), .A(N3620), .B(N3593));
NOR2XL inst_cellmath__43_0_I299 (.Y(N812), .A(N3620), .B(N3594));
NOR2XL inst_cellmath__43_0_I300 (.Y(N814), .A(N3620), .B(N3595));
NOR2XL inst_cellmath__43_0_I301 (.Y(N816), .A(N3620), .B(N3596));
NOR2XL inst_cellmath__43_0_I302 (.Y(N818), .A(N3620), .B(N3597));
NOR2XL inst_cellmath__43_0_I303 (.Y(N820), .A(N3620), .B(N3598));
NOR2XL inst_cellmath__43_0_I304 (.Y(N822), .A(N3620), .B(N3599));
NOR2XL inst_cellmath__43_0_I305 (.Y(N824), .A(N3620), .B(N3600));
NOR2XL inst_cellmath__43_0_I306 (.Y(N826), .A(N3620), .B(N3601));
NOR2XL inst_cellmath__43_0_I307 (.Y(N828), .A(N3620), .B(N3602));
NOR2XL inst_cellmath__43_0_I308 (.Y(N830), .A(N3620), .B(N3603));
NOR2XL inst_cellmath__43_0_I309 (.Y(N832), .A(N3620), .B(N3604));
NOR2XL inst_cellmath__43_0_I310 (.Y(N834), .A(N3620), .B(N3605));
NOR2XL inst_cellmath__43_0_I311 (.Y(N836), .A(N3620), .B(N3606));
NOR2XL inst_cellmath__43_0_I312 (.Y(N838), .A(N3620), .B(N3607));
INVXL inst_cellmath__43_0_I313 (.Y(N840), .A(N3620));
INVXL inst_cellmath__43_0_I2027 (.Y(N3621), .A(inst_cellmath__43_0_in1[8]));
NOR2XL inst_cellmath__43_0_I319 (.Y(N853), .A(N3621), .B(N3585));
NOR2XL inst_cellmath__43_0_I320 (.Y(N855), .A(N3621), .B(N3586));
NOR2XL inst_cellmath__43_0_I321 (.Y(N857), .A(N3621), .B(N3587));
NOR2XL inst_cellmath__43_0_I322 (.Y(N859), .A(N3621), .B(N3588));
NOR2XL inst_cellmath__43_0_I323 (.Y(N861), .A(N3621), .B(N3589));
NOR2XL inst_cellmath__43_0_I324 (.Y(N863), .A(N3621), .B(N3590));
NOR2XL inst_cellmath__43_0_I325 (.Y(N865), .A(N3621), .B(N3591));
NOR2XL inst_cellmath__43_0_I326 (.Y(N867), .A(N3621), .B(N3592));
NOR2XL inst_cellmath__43_0_I327 (.Y(N869), .A(N3621), .B(N3593));
NOR2XL inst_cellmath__43_0_I328 (.Y(N871), .A(N3621), .B(N3594));
NOR2XL inst_cellmath__43_0_I329 (.Y(N873), .A(N3621), .B(N3595));
NOR2XL inst_cellmath__43_0_I330 (.Y(N875), .A(N3621), .B(N3596));
NOR2XL inst_cellmath__43_0_I331 (.Y(N877), .A(N3621), .B(N3597));
NOR2XL inst_cellmath__43_0_I332 (.Y(N879), .A(N3621), .B(N3598));
NOR2XL inst_cellmath__43_0_I333 (.Y(N881), .A(N3621), .B(N3599));
NOR2XL inst_cellmath__43_0_I334 (.Y(N883), .A(N3621), .B(N3600));
NOR2XL inst_cellmath__43_0_I335 (.Y(N885), .A(N3621), .B(N3601));
NOR2XL inst_cellmath__43_0_I336 (.Y(N887), .A(N3621), .B(N3602));
NOR2XL inst_cellmath__43_0_I337 (.Y(N889), .A(N3621), .B(N3603));
NOR2XL inst_cellmath__43_0_I338 (.Y(N891), .A(N3621), .B(N3604));
NOR2XL inst_cellmath__43_0_I339 (.Y(N893), .A(N3621), .B(N3605));
NOR2XL inst_cellmath__43_0_I340 (.Y(N895), .A(N3621), .B(N3606));
NOR2XL inst_cellmath__43_0_I341 (.Y(N897), .A(N3621), .B(N3607));
INVXL inst_cellmath__43_0_I342 (.Y(N899), .A(N3621));
INVXL inst_cellmath__43_0_I2028 (.Y(N3622), .A(inst_cellmath__43_0_in1[9]));
NOR2XL inst_cellmath__43_0_I348 (.Y(N912), .A(N3622), .B(N3585));
NOR2XL inst_cellmath__43_0_I349 (.Y(N914), .A(N3622), .B(N3586));
NOR2XL inst_cellmath__43_0_I350 (.Y(N916), .A(N3622), .B(N3587));
NOR2XL inst_cellmath__43_0_I351 (.Y(N918), .A(N3622), .B(N3588));
NOR2XL inst_cellmath__43_0_I352 (.Y(N920), .A(N3622), .B(N3589));
NOR2XL inst_cellmath__43_0_I353 (.Y(N922), .A(N3622), .B(N3590));
NOR2XL inst_cellmath__43_0_I354 (.Y(N924), .A(N3622), .B(N3591));
NOR2XL inst_cellmath__43_0_I355 (.Y(N926), .A(N3622), .B(N3592));
NOR2XL inst_cellmath__43_0_I356 (.Y(N928), .A(N3622), .B(N3593));
NOR2XL inst_cellmath__43_0_I357 (.Y(N930), .A(N3622), .B(N3594));
NOR2XL inst_cellmath__43_0_I358 (.Y(N932), .A(N3622), .B(N3595));
NOR2XL inst_cellmath__43_0_I359 (.Y(N934), .A(N3622), .B(N3596));
NOR2XL inst_cellmath__43_0_I360 (.Y(N936), .A(N3622), .B(N3597));
NOR2XL inst_cellmath__43_0_I361 (.Y(N938), .A(N3622), .B(N3598));
NOR2XL inst_cellmath__43_0_I362 (.Y(N940), .A(N3622), .B(N3599));
NOR2XL inst_cellmath__43_0_I363 (.Y(N942), .A(N3622), .B(N3600));
NOR2XL inst_cellmath__43_0_I364 (.Y(N944), .A(N3622), .B(N3601));
NOR2XL inst_cellmath__43_0_I365 (.Y(N946), .A(N3622), .B(N3602));
NOR2XL inst_cellmath__43_0_I366 (.Y(N948), .A(N3622), .B(N3603));
NOR2XL inst_cellmath__43_0_I367 (.Y(N950), .A(N3622), .B(N3604));
NOR2XL inst_cellmath__43_0_I368 (.Y(N952), .A(N3622), .B(N3605));
NOR2XL inst_cellmath__43_0_I369 (.Y(N954), .A(N3622), .B(N3606));
NOR2XL inst_cellmath__43_0_I370 (.Y(N956), .A(N3622), .B(N3607));
INVXL inst_cellmath__43_0_I371 (.Y(N958), .A(N3622));
INVXL inst_cellmath__43_0_I2029 (.Y(N3623), .A(inst_cellmath__43_0_in1[10]));
NOR2XL inst_cellmath__43_0_I377 (.Y(N971), .A(N3623), .B(N3585));
NOR2XL inst_cellmath__43_0_I378 (.Y(N973), .A(N3623), .B(N3586));
NOR2XL inst_cellmath__43_0_I379 (.Y(N975), .A(N3623), .B(N3587));
NOR2XL inst_cellmath__43_0_I380 (.Y(N977), .A(N3623), .B(N3588));
NOR2XL inst_cellmath__43_0_I381 (.Y(N979), .A(N3623), .B(N3589));
NOR2XL inst_cellmath__43_0_I382 (.Y(N981), .A(N3623), .B(N3590));
NOR2XL inst_cellmath__43_0_I383 (.Y(N983), .A(N3623), .B(N3591));
NOR2XL inst_cellmath__43_0_I384 (.Y(N985), .A(N3623), .B(N3592));
NOR2XL inst_cellmath__43_0_I385 (.Y(N987), .A(N3623), .B(N3593));
NOR2XL inst_cellmath__43_0_I386 (.Y(N989), .A(N3623), .B(N3594));
NOR2XL inst_cellmath__43_0_I387 (.Y(N991), .A(N3623), .B(N3595));
NOR2XL inst_cellmath__43_0_I388 (.Y(N993), .A(N3623), .B(N3596));
NOR2XL inst_cellmath__43_0_I389 (.Y(N995), .A(N3623), .B(N3597));
NOR2XL inst_cellmath__43_0_I390 (.Y(N997), .A(N3623), .B(N3598));
NOR2XL inst_cellmath__43_0_I391 (.Y(N999), .A(N3623), .B(N3599));
NOR2XL inst_cellmath__43_0_I392 (.Y(N1001), .A(N3623), .B(N3600));
NOR2XL inst_cellmath__43_0_I393 (.Y(N1003), .A(N3623), .B(N3601));
NOR2XL inst_cellmath__43_0_I394 (.Y(N1005), .A(N3623), .B(N3602));
NOR2XL inst_cellmath__43_0_I395 (.Y(N1007), .A(N3623), .B(N3603));
NOR2XL inst_cellmath__43_0_I396 (.Y(N1009), .A(N3623), .B(N3604));
NOR2XL inst_cellmath__43_0_I397 (.Y(N1011), .A(N3623), .B(N3605));
NOR2XL inst_cellmath__43_0_I398 (.Y(N1013), .A(N3623), .B(N3606));
NOR2XL inst_cellmath__43_0_I399 (.Y(N1015), .A(N3623), .B(N3607));
INVXL inst_cellmath__43_0_I400 (.Y(N1017), .A(N3623));
INVXL inst_cellmath__43_0_I2030 (.Y(N3624), .A(inst_cellmath__43_0_in1[11]));
NOR2XL inst_cellmath__43_0_I406 (.Y(N1030), .A(N3624), .B(N3585));
NOR2XL inst_cellmath__43_0_I407 (.Y(N1032), .A(N3624), .B(N3586));
NOR2XL inst_cellmath__43_0_I408 (.Y(N1034), .A(N3624), .B(N3587));
NOR2XL inst_cellmath__43_0_I409 (.Y(N1036), .A(N3624), .B(N3588));
NOR2XL inst_cellmath__43_0_I410 (.Y(N1038), .A(N3624), .B(N3589));
NOR2XL inst_cellmath__43_0_I411 (.Y(N1040), .A(N3624), .B(N3590));
NOR2XL inst_cellmath__43_0_I412 (.Y(N1042), .A(N3624), .B(N3591));
NOR2XL inst_cellmath__43_0_I413 (.Y(N1044), .A(N3624), .B(N3592));
NOR2XL inst_cellmath__43_0_I414 (.Y(N1046), .A(N3624), .B(N3593));
NOR2XL inst_cellmath__43_0_I415 (.Y(N1048), .A(N3624), .B(N3594));
NOR2XL inst_cellmath__43_0_I416 (.Y(N1050), .A(N3624), .B(N3595));
NOR2XL inst_cellmath__43_0_I417 (.Y(N1052), .A(N3624), .B(N3596));
NOR2XL inst_cellmath__43_0_I418 (.Y(N1054), .A(N3624), .B(N3597));
NOR2XL inst_cellmath__43_0_I419 (.Y(N1056), .A(N3624), .B(N3598));
NOR2XL inst_cellmath__43_0_I420 (.Y(N1058), .A(N3624), .B(N3599));
NOR2XL inst_cellmath__43_0_I421 (.Y(N1060), .A(N3624), .B(N3600));
NOR2XL inst_cellmath__43_0_I422 (.Y(N1062), .A(N3624), .B(N3601));
NOR2XL inst_cellmath__43_0_I423 (.Y(N1064), .A(N3624), .B(N3602));
NOR2XL inst_cellmath__43_0_I424 (.Y(N1066), .A(N3624), .B(N3603));
NOR2XL inst_cellmath__43_0_I425 (.Y(N1068), .A(N3624), .B(N3604));
NOR2XL inst_cellmath__43_0_I426 (.Y(N1070), .A(N3624), .B(N3605));
NOR2XL inst_cellmath__43_0_I427 (.Y(N1072), .A(N3624), .B(N3606));
NOR2XL inst_cellmath__43_0_I428 (.Y(N1074), .A(N3624), .B(N3607));
INVXL inst_cellmath__43_0_I429 (.Y(N1076), .A(N3624));
INVXL inst_cellmath__43_0_I2031 (.Y(N3625), .A(inst_cellmath__43_0_in1[12]));
NOR2XL inst_cellmath__43_0_I435 (.Y(N1089), .A(N3625), .B(N3585));
NOR2XL inst_cellmath__43_0_I436 (.Y(N1091), .A(N3625), .B(N3586));
NOR2XL inst_cellmath__43_0_I437 (.Y(N1093), .A(N3625), .B(N3587));
NOR2XL inst_cellmath__43_0_I438 (.Y(N1095), .A(N3625), .B(N3588));
NOR2XL inst_cellmath__43_0_I439 (.Y(N1097), .A(N3625), .B(N3589));
NOR2XL inst_cellmath__43_0_I440 (.Y(N1099), .A(N3625), .B(N3590));
NOR2XL inst_cellmath__43_0_I441 (.Y(N1101), .A(N3625), .B(N3591));
NOR2XL inst_cellmath__43_0_I442 (.Y(N1103), .A(N3625), .B(N3592));
NOR2XL inst_cellmath__43_0_I443 (.Y(N1105), .A(N3625), .B(N3593));
NOR2XL inst_cellmath__43_0_I444 (.Y(N1107), .A(N3625), .B(N3594));
NOR2XL inst_cellmath__43_0_I445 (.Y(N1109), .A(N3625), .B(N3595));
NOR2XL inst_cellmath__43_0_I446 (.Y(N1111), .A(N3625), .B(N3596));
NOR2XL inst_cellmath__43_0_I447 (.Y(N1113), .A(N3625), .B(N3597));
NOR2XL inst_cellmath__43_0_I448 (.Y(N1115), .A(N3625), .B(N3598));
NOR2XL inst_cellmath__43_0_I449 (.Y(N1117), .A(N3625), .B(N3599));
NOR2XL inst_cellmath__43_0_I450 (.Y(N1119), .A(N3625), .B(N3600));
NOR2XL inst_cellmath__43_0_I451 (.Y(N1121), .A(N3625), .B(N3601));
NOR2XL inst_cellmath__43_0_I452 (.Y(N1123), .A(N3625), .B(N3602));
NOR2XL inst_cellmath__43_0_I453 (.Y(N1125), .A(N3625), .B(N3603));
NOR2XL inst_cellmath__43_0_I454 (.Y(N1127), .A(N3625), .B(N3604));
NOR2XL inst_cellmath__43_0_I455 (.Y(N1129), .A(N3625), .B(N3605));
NOR2XL inst_cellmath__43_0_I456 (.Y(N1131), .A(N3625), .B(N3606));
NOR2XL inst_cellmath__43_0_I457 (.Y(N1133), .A(N3625), .B(N3607));
INVXL inst_cellmath__43_0_I458 (.Y(N1135), .A(N3625));
INVXL inst_cellmath__43_0_I2032 (.Y(N3626), .A(inst_cellmath__43_0_in1[13]));
NOR2XL inst_cellmath__43_0_I464 (.Y(N1148), .A(N3626), .B(N3585));
NOR2XL inst_cellmath__43_0_I465 (.Y(N1150), .A(N3626), .B(N3586));
NOR2XL inst_cellmath__43_0_I466 (.Y(N1152), .A(N3626), .B(N3587));
NOR2XL inst_cellmath__43_0_I467 (.Y(N1154), .A(N3626), .B(N3588));
NOR2XL inst_cellmath__43_0_I468 (.Y(N1156), .A(N3626), .B(N3589));
NOR2XL inst_cellmath__43_0_I469 (.Y(N1158), .A(N3626), .B(N3590));
NOR2XL inst_cellmath__43_0_I470 (.Y(N1160), .A(N3626), .B(N3591));
NOR2XL inst_cellmath__43_0_I471 (.Y(N1162), .A(N3626), .B(N3592));
NOR2XL inst_cellmath__43_0_I472 (.Y(N1164), .A(N3626), .B(N3593));
NOR2XL inst_cellmath__43_0_I473 (.Y(N1166), .A(N3626), .B(N3594));
NOR2XL inst_cellmath__43_0_I474 (.Y(N1168), .A(N3626), .B(N3595));
NOR2XL inst_cellmath__43_0_I475 (.Y(N1170), .A(N3626), .B(N3596));
NOR2XL inst_cellmath__43_0_I476 (.Y(N1172), .A(N3626), .B(N3597));
NOR2XL inst_cellmath__43_0_I477 (.Y(N1174), .A(N3626), .B(N3598));
NOR2XL inst_cellmath__43_0_I478 (.Y(N1176), .A(N3626), .B(N3599));
NOR2XL inst_cellmath__43_0_I479 (.Y(N1178), .A(N3626), .B(N3600));
NOR2XL inst_cellmath__43_0_I480 (.Y(N1180), .A(N3626), .B(N3601));
NOR2XL inst_cellmath__43_0_I481 (.Y(N1182), .A(N3626), .B(N3602));
NOR2XL inst_cellmath__43_0_I482 (.Y(N1184), .A(N3626), .B(N3603));
NOR2XL inst_cellmath__43_0_I483 (.Y(N1186), .A(N3626), .B(N3604));
NOR2XL inst_cellmath__43_0_I484 (.Y(N1188), .A(N3626), .B(N3605));
NOR2XL inst_cellmath__43_0_I485 (.Y(N1190), .A(N3626), .B(N3606));
NOR2XL inst_cellmath__43_0_I486 (.Y(N1192), .A(N3626), .B(N3607));
INVXL inst_cellmath__43_0_I487 (.Y(N1194), .A(N3626));
INVXL inst_cellmath__43_0_I2033 (.Y(N3627), .A(inst_cellmath__43_0_in1[14]));
NOR2XL inst_cellmath__43_0_I493 (.Y(N1207), .A(N3627), .B(N3585));
NOR2XL inst_cellmath__43_0_I494 (.Y(N1209), .A(N3627), .B(N3586));
NOR2XL inst_cellmath__43_0_I495 (.Y(N1211), .A(N3627), .B(N3587));
NOR2XL inst_cellmath__43_0_I496 (.Y(N1213), .A(N3627), .B(N3588));
NOR2XL inst_cellmath__43_0_I497 (.Y(N1215), .A(N3627), .B(N3589));
NOR2XL inst_cellmath__43_0_I498 (.Y(N1217), .A(N3627), .B(N3590));
NOR2XL inst_cellmath__43_0_I499 (.Y(N1219), .A(N3627), .B(N3591));
NOR2XL inst_cellmath__43_0_I500 (.Y(N1221), .A(N3627), .B(N3592));
NOR2XL inst_cellmath__43_0_I501 (.Y(N1223), .A(N3627), .B(N3593));
NOR2XL inst_cellmath__43_0_I502 (.Y(N1225), .A(N3627), .B(N3594));
NOR2XL inst_cellmath__43_0_I503 (.Y(N1227), .A(N3627), .B(N3595));
NOR2XL inst_cellmath__43_0_I504 (.Y(N1229), .A(N3627), .B(N3596));
NOR2XL inst_cellmath__43_0_I505 (.Y(N1231), .A(N3627), .B(N3597));
NOR2XL inst_cellmath__43_0_I506 (.Y(N1233), .A(N3627), .B(N3598));
NOR2XL inst_cellmath__43_0_I507 (.Y(N1235), .A(N3627), .B(N3599));
NOR2XL inst_cellmath__43_0_I508 (.Y(N1237), .A(N3627), .B(N3600));
NOR2XL inst_cellmath__43_0_I509 (.Y(N1239), .A(N3627), .B(N3601));
NOR2XL inst_cellmath__43_0_I510 (.Y(N1241), .A(N3627), .B(N3602));
NOR2XL inst_cellmath__43_0_I511 (.Y(N1243), .A(N3627), .B(N3603));
NOR2XL inst_cellmath__43_0_I512 (.Y(N1245), .A(N3627), .B(N3604));
NOR2XL inst_cellmath__43_0_I513 (.Y(N1247), .A(N3627), .B(N3605));
NOR2XL inst_cellmath__43_0_I514 (.Y(N1249), .A(N3627), .B(N3606));
NOR2XL inst_cellmath__43_0_I515 (.Y(N1251), .A(N3627), .B(N3607));
INVXL inst_cellmath__43_0_I516 (.Y(N1253), .A(N3627));
INVXL inst_cellmath__43_0_I2034 (.Y(N3628), .A(inst_cellmath__43_0_in1[15]));
NOR2XL inst_cellmath__43_0_I522 (.Y(N1266), .A(N3628), .B(N3585));
NOR2XL inst_cellmath__43_0_I523 (.Y(N1268), .A(N3628), .B(N3586));
NOR2XL inst_cellmath__43_0_I524 (.Y(N1270), .A(N3628), .B(N3587));
NOR2XL inst_cellmath__43_0_I525 (.Y(N1272), .A(N3628), .B(N3588));
NOR2XL inst_cellmath__43_0_I526 (.Y(N1274), .A(N3628), .B(N3589));
NOR2XL inst_cellmath__43_0_I527 (.Y(N1276), .A(N3628), .B(N3590));
NOR2XL inst_cellmath__43_0_I528 (.Y(N1278), .A(N3628), .B(N3591));
NOR2XL inst_cellmath__43_0_I529 (.Y(N1280), .A(N3628), .B(N3592));
NOR2XL inst_cellmath__43_0_I530 (.Y(N1282), .A(N3628), .B(N3593));
NOR2XL inst_cellmath__43_0_I531 (.Y(N1284), .A(N3628), .B(N3594));
NOR2XL inst_cellmath__43_0_I532 (.Y(N1286), .A(N3628), .B(N3595));
NOR2XL inst_cellmath__43_0_I533 (.Y(N1288), .A(N3628), .B(N3596));
NOR2XL inst_cellmath__43_0_I534 (.Y(N1290), .A(N3628), .B(N3597));
NOR2XL inst_cellmath__43_0_I535 (.Y(N1292), .A(N3628), .B(N3598));
NOR2XL inst_cellmath__43_0_I536 (.Y(N1294), .A(N3628), .B(N3599));
NOR2XL inst_cellmath__43_0_I537 (.Y(N1296), .A(N3628), .B(N3600));
NOR2XL inst_cellmath__43_0_I538 (.Y(N1298), .A(N3628), .B(N3601));
NOR2XL inst_cellmath__43_0_I539 (.Y(N1300), .A(N3628), .B(N3602));
NOR2XL inst_cellmath__43_0_I540 (.Y(N1302), .A(N3628), .B(N3603));
NOR2XL inst_cellmath__43_0_I541 (.Y(N1304), .A(N3628), .B(N3604));
NOR2XL inst_cellmath__43_0_I542 (.Y(N1306), .A(N3628), .B(N3605));
NOR2XL inst_cellmath__43_0_I543 (.Y(N1308), .A(N3628), .B(N3606));
NOR2XL inst_cellmath__43_0_I544 (.Y(N1310), .A(N3628), .B(N3607));
INVXL inst_cellmath__43_0_I545 (.Y(N1312), .A(N3628));
INVXL inst_cellmath__43_0_I2035 (.Y(N3629), .A(inst_cellmath__43_0_in1[16]));
NOR2XL inst_cellmath__43_0_I551 (.Y(N1325), .A(N3629), .B(N3585));
NOR2XL inst_cellmath__43_0_I552 (.Y(N1327), .A(N3629), .B(N3586));
NOR2XL inst_cellmath__43_0_I553 (.Y(N1329), .A(N3629), .B(N3587));
NOR2XL inst_cellmath__43_0_I554 (.Y(N1331), .A(N3629), .B(N3588));
NOR2XL inst_cellmath__43_0_I555 (.Y(N1333), .A(N3629), .B(N3589));
NOR2XL inst_cellmath__43_0_I556 (.Y(N1335), .A(N3629), .B(N3590));
NOR2XL inst_cellmath__43_0_I557 (.Y(N1337), .A(N3629), .B(N3591));
NOR2XL inst_cellmath__43_0_I558 (.Y(N1339), .A(N3629), .B(N3592));
NOR2XL inst_cellmath__43_0_I559 (.Y(N1341), .A(N3629), .B(N3593));
NOR2XL inst_cellmath__43_0_I560 (.Y(N1343), .A(N3629), .B(N3594));
NOR2XL inst_cellmath__43_0_I561 (.Y(N1345), .A(N3629), .B(N3595));
NOR2XL inst_cellmath__43_0_I562 (.Y(N1347), .A(N3629), .B(N3596));
NOR2XL inst_cellmath__43_0_I563 (.Y(N1349), .A(N3629), .B(N3597));
NOR2XL inst_cellmath__43_0_I564 (.Y(N1351), .A(N3629), .B(N3598));
NOR2XL inst_cellmath__43_0_I565 (.Y(N1353), .A(N3629), .B(N3599));
NOR2XL inst_cellmath__43_0_I566 (.Y(N1355), .A(N3629), .B(N3600));
NOR2XL inst_cellmath__43_0_I567 (.Y(N1357), .A(N3629), .B(N3601));
NOR2XL inst_cellmath__43_0_I568 (.Y(N1359), .A(N3629), .B(N3602));
NOR2XL inst_cellmath__43_0_I569 (.Y(N1361), .A(N3629), .B(N3603));
NOR2XL inst_cellmath__43_0_I570 (.Y(N1363), .A(N3629), .B(N3604));
NOR2XL inst_cellmath__43_0_I571 (.Y(N1365), .A(N3629), .B(N3605));
NOR2XL inst_cellmath__43_0_I572 (.Y(N1367), .A(N3629), .B(N3606));
NOR2XL inst_cellmath__43_0_I573 (.Y(N1369), .A(N3629), .B(N3607));
INVXL inst_cellmath__43_0_I574 (.Y(N1371), .A(N3629));
INVXL inst_cellmath__43_0_I2036 (.Y(N3630), .A(inst_cellmath__43_0_in1[17]));
NOR2XL inst_cellmath__43_0_I580 (.Y(N1384), .A(N3630), .B(N3585));
NOR2XL inst_cellmath__43_0_I581 (.Y(N1386), .A(N3630), .B(N3586));
NOR2XL inst_cellmath__43_0_I582 (.Y(N1388), .A(N3630), .B(N3587));
NOR2XL inst_cellmath__43_0_I583 (.Y(N1390), .A(N3630), .B(N3588));
NOR2XL inst_cellmath__43_0_I584 (.Y(N1392), .A(N3630), .B(N3589));
NOR2XL inst_cellmath__43_0_I585 (.Y(N1394), .A(N3630), .B(N3590));
NOR2XL inst_cellmath__43_0_I586 (.Y(N1396), .A(N3630), .B(N3591));
NOR2XL inst_cellmath__43_0_I587 (.Y(N1398), .A(N3630), .B(N3592));
NOR2XL inst_cellmath__43_0_I588 (.Y(N1400), .A(N3630), .B(N3593));
NOR2XL inst_cellmath__43_0_I589 (.Y(N1402), .A(N3630), .B(N3594));
NOR2XL inst_cellmath__43_0_I590 (.Y(N1404), .A(N3630), .B(N3595));
NOR2XL inst_cellmath__43_0_I591 (.Y(N1406), .A(N3630), .B(N3596));
NOR2XL inst_cellmath__43_0_I592 (.Y(N1408), .A(N3630), .B(N3597));
NOR2XL inst_cellmath__43_0_I593 (.Y(N1410), .A(N3630), .B(N3598));
NOR2XL inst_cellmath__43_0_I594 (.Y(N1412), .A(N3630), .B(N3599));
NOR2XL inst_cellmath__43_0_I595 (.Y(N1414), .A(N3630), .B(N3600));
NOR2XL inst_cellmath__43_0_I596 (.Y(N1416), .A(N3630), .B(N3601));
NOR2XL inst_cellmath__43_0_I597 (.Y(N1418), .A(N3630), .B(N3602));
NOR2XL inst_cellmath__43_0_I598 (.Y(N1420), .A(N3630), .B(N3603));
NOR2XL inst_cellmath__43_0_I599 (.Y(N1422), .A(N3630), .B(N3604));
NOR2XL inst_cellmath__43_0_I600 (.Y(N1424), .A(N3630), .B(N3605));
NOR2XL inst_cellmath__43_0_I601 (.Y(N1426), .A(N3630), .B(N3606));
NOR2XL inst_cellmath__43_0_I602 (.Y(N1428), .A(N3630), .B(N3607));
INVXL inst_cellmath__43_0_I603 (.Y(N1430), .A(N3630));
INVXL inst_cellmath__43_0_I2037 (.Y(N3631), .A(inst_cellmath__43_0_in1[18]));
NOR2XL inst_cellmath__43_0_I609 (.Y(N1443), .A(N3631), .B(N3585));
NOR2XL inst_cellmath__43_0_I610 (.Y(N1445), .A(N3631), .B(N3586));
NOR2XL inst_cellmath__43_0_I611 (.Y(N1447), .A(N3631), .B(N3587));
NOR2XL inst_cellmath__43_0_I612 (.Y(N1449), .A(N3631), .B(N3588));
NOR2XL inst_cellmath__43_0_I613 (.Y(N1451), .A(N3631), .B(N3589));
NOR2XL inst_cellmath__43_0_I614 (.Y(N1453), .A(N3631), .B(N3590));
NOR2XL inst_cellmath__43_0_I615 (.Y(N1455), .A(N3631), .B(N3591));
NOR2XL inst_cellmath__43_0_I616 (.Y(N1457), .A(N3631), .B(N3592));
NOR2XL inst_cellmath__43_0_I617 (.Y(N1459), .A(N3631), .B(N3593));
NOR2XL inst_cellmath__43_0_I618 (.Y(N1461), .A(N3631), .B(N3594));
NOR2XL inst_cellmath__43_0_I619 (.Y(N1463), .A(N3631), .B(N3595));
NOR2XL inst_cellmath__43_0_I620 (.Y(N1465), .A(N3631), .B(N3596));
NOR2XL inst_cellmath__43_0_I621 (.Y(N1467), .A(N3631), .B(N3597));
NOR2XL inst_cellmath__43_0_I622 (.Y(N1469), .A(N3631), .B(N3598));
NOR2XL inst_cellmath__43_0_I623 (.Y(N1471), .A(N3631), .B(N3599));
NOR2XL inst_cellmath__43_0_I624 (.Y(N1473), .A(N3631), .B(N3600));
NOR2XL inst_cellmath__43_0_I625 (.Y(N1475), .A(N3631), .B(N3601));
NOR2XL inst_cellmath__43_0_I626 (.Y(N1477), .A(N3631), .B(N3602));
NOR2XL inst_cellmath__43_0_I627 (.Y(N1479), .A(N3631), .B(N3603));
NOR2XL inst_cellmath__43_0_I628 (.Y(N1481), .A(N3631), .B(N3604));
NOR2XL inst_cellmath__43_0_I629 (.Y(N1483), .A(N3631), .B(N3605));
NOR2XL inst_cellmath__43_0_I630 (.Y(N1485), .A(N3631), .B(N3606));
NOR2XL inst_cellmath__43_0_I631 (.Y(N1487), .A(N3631), .B(N3607));
INVXL inst_cellmath__43_0_I632 (.Y(N1489), .A(N3631));
INVXL inst_cellmath__43_0_I2038 (.Y(N3632), .A(inst_cellmath__43_0_in1[19]));
NOR2XL inst_cellmath__43_0_I638 (.Y(N1502), .A(N3632), .B(N3585));
NOR2XL inst_cellmath__43_0_I639 (.Y(N1504), .A(N3632), .B(N3586));
NOR2XL inst_cellmath__43_0_I640 (.Y(N1506), .A(N3632), .B(N3587));
NOR2XL inst_cellmath__43_0_I641 (.Y(N1508), .A(N3632), .B(N3588));
NOR2XL inst_cellmath__43_0_I642 (.Y(N1510), .A(N3632), .B(N3589));
NOR2XL inst_cellmath__43_0_I643 (.Y(N1512), .A(N3632), .B(N3590));
NOR2XL inst_cellmath__43_0_I644 (.Y(N1514), .A(N3632), .B(N3591));
NOR2XL inst_cellmath__43_0_I645 (.Y(N1516), .A(N3632), .B(N3592));
NOR2XL inst_cellmath__43_0_I646 (.Y(N1518), .A(N3632), .B(N3593));
NOR2XL inst_cellmath__43_0_I647 (.Y(N1520), .A(N3632), .B(N3594));
NOR2XL inst_cellmath__43_0_I648 (.Y(N1522), .A(N3632), .B(N3595));
NOR2XL inst_cellmath__43_0_I649 (.Y(N1524), .A(N3632), .B(N3596));
NOR2XL inst_cellmath__43_0_I650 (.Y(N1526), .A(N3632), .B(N3597));
NOR2XL inst_cellmath__43_0_I651 (.Y(N1528), .A(N3632), .B(N3598));
NOR2XL inst_cellmath__43_0_I652 (.Y(N1530), .A(N3632), .B(N3599));
NOR2XL inst_cellmath__43_0_I653 (.Y(N1532), .A(N3632), .B(N3600));
NOR2XL inst_cellmath__43_0_I654 (.Y(N1534), .A(N3632), .B(N3601));
NOR2XL inst_cellmath__43_0_I655 (.Y(N1536), .A(N3632), .B(N3602));
NOR2XL inst_cellmath__43_0_I656 (.Y(N1538), .A(N3632), .B(N3603));
NOR2XL inst_cellmath__43_0_I657 (.Y(N1540), .A(N3632), .B(N3604));
NOR2XL inst_cellmath__43_0_I658 (.Y(N1542), .A(N3632), .B(N3605));
NOR2XL inst_cellmath__43_0_I659 (.Y(N1544), .A(N3632), .B(N3606));
NOR2XL inst_cellmath__43_0_I660 (.Y(N1546), .A(N3632), .B(N3607));
INVXL inst_cellmath__43_0_I661 (.Y(N1548), .A(N3632));
INVXL inst_cellmath__43_0_I2039 (.Y(N3633), .A(inst_cellmath__43_0_in1[20]));
NOR2XL inst_cellmath__43_0_I667 (.Y(N1561), .A(N3633), .B(N3585));
NOR2XL inst_cellmath__43_0_I668 (.Y(N1563), .A(N3633), .B(N3586));
NOR2XL inst_cellmath__43_0_I669 (.Y(N1565), .A(N3633), .B(N3587));
NOR2XL inst_cellmath__43_0_I670 (.Y(N1567), .A(N3633), .B(N3588));
NOR2XL inst_cellmath__43_0_I671 (.Y(N1569), .A(N3633), .B(N3589));
NOR2XL inst_cellmath__43_0_I672 (.Y(N1571), .A(N3633), .B(N3590));
NOR2XL inst_cellmath__43_0_I673 (.Y(N1573), .A(N3633), .B(N3591));
NOR2XL inst_cellmath__43_0_I674 (.Y(N1575), .A(N3633), .B(N3592));
NOR2XL inst_cellmath__43_0_I675 (.Y(N1577), .A(N3633), .B(N3593));
NOR2XL inst_cellmath__43_0_I676 (.Y(N1579), .A(N3633), .B(N3594));
NOR2XL inst_cellmath__43_0_I677 (.Y(N1581), .A(N3633), .B(N3595));
NOR2XL inst_cellmath__43_0_I678 (.Y(N1583), .A(N3633), .B(N3596));
NOR2XL inst_cellmath__43_0_I679 (.Y(N1585), .A(N3633), .B(N3597));
NOR2XL inst_cellmath__43_0_I680 (.Y(N1587), .A(N3633), .B(N3598));
NOR2XL inst_cellmath__43_0_I681 (.Y(N1589), .A(N3633), .B(N3599));
NOR2XL inst_cellmath__43_0_I682 (.Y(N1591), .A(N3633), .B(N3600));
NOR2XL inst_cellmath__43_0_I683 (.Y(N1593), .A(N3633), .B(N3601));
NOR2XL inst_cellmath__43_0_I684 (.Y(N1595), .A(N3633), .B(N3602));
NOR2XL inst_cellmath__43_0_I685 (.Y(N1597), .A(N3633), .B(N3603));
NOR2XL inst_cellmath__43_0_I686 (.Y(N1599), .A(N3633), .B(N3604));
NOR2XL inst_cellmath__43_0_I687 (.Y(N1601), .A(N3633), .B(N3605));
NOR2XL inst_cellmath__43_0_I688 (.Y(N1603), .A(N3633), .B(N3606));
NOR2XL inst_cellmath__43_0_I689 (.Y(N1605), .A(N3633), .B(N3607));
INVXL inst_cellmath__43_0_I690 (.Y(N1607), .A(N3633));
INVXL inst_cellmath__43_0_I2040 (.Y(N3634), .A(inst_cellmath__43_0_in1[21]));
NOR2XL inst_cellmath__43_0_I696 (.Y(N1620), .A(N3634), .B(N3585));
NOR2XL inst_cellmath__43_0_I697 (.Y(N1622), .A(N3634), .B(N3586));
NOR2XL inst_cellmath__43_0_I698 (.Y(N1624), .A(N3634), .B(N3587));
NOR2XL inst_cellmath__43_0_I699 (.Y(N1626), .A(N3634), .B(N3588));
NOR2XL inst_cellmath__43_0_I700 (.Y(N1628), .A(N3634), .B(N3589));
NOR2XL inst_cellmath__43_0_I701 (.Y(N1630), .A(N3634), .B(N3590));
NOR2XL inst_cellmath__43_0_I702 (.Y(N1632), .A(N3634), .B(N3591));
NOR2XL inst_cellmath__43_0_I703 (.Y(N1634), .A(N3634), .B(N3592));
NOR2XL inst_cellmath__43_0_I704 (.Y(N1636), .A(N3634), .B(N3593));
NOR2XL inst_cellmath__43_0_I705 (.Y(N1638), .A(N3634), .B(N3594));
NOR2XL inst_cellmath__43_0_I706 (.Y(N1640), .A(N3634), .B(N3595));
NOR2XL inst_cellmath__43_0_I707 (.Y(N1642), .A(N3634), .B(N3596));
NOR2XL inst_cellmath__43_0_I708 (.Y(N1644), .A(N3634), .B(N3597));
NOR2XL inst_cellmath__43_0_I709 (.Y(N1646), .A(N3634), .B(N3598));
NOR2XL inst_cellmath__43_0_I710 (.Y(N1648), .A(N3634), .B(N3599));
NOR2XL inst_cellmath__43_0_I711 (.Y(N1650), .A(N3634), .B(N3600));
NOR2XL inst_cellmath__43_0_I712 (.Y(N1652), .A(N3634), .B(N3601));
NOR2XL inst_cellmath__43_0_I713 (.Y(N1654), .A(N3634), .B(N3602));
NOR2XL inst_cellmath__43_0_I714 (.Y(N1656), .A(N3634), .B(N3603));
NOR2XL inst_cellmath__43_0_I715 (.Y(N1658), .A(N3634), .B(N3604));
NOR2XL inst_cellmath__43_0_I716 (.Y(N1660), .A(N3634), .B(N3605));
NOR2XL inst_cellmath__43_0_I717 (.Y(N1662), .A(N3634), .B(N3606));
NOR2XL inst_cellmath__43_0_I718 (.Y(N1664), .A(N3634), .B(N3607));
INVXL inst_cellmath__43_0_I719 (.Y(N1666), .A(N3634));
INVXL inst_cellmath__43_0_I2041 (.Y(N3635), .A(inst_cellmath__43_0_in1[22]));
NOR2XL inst_cellmath__43_0_I725 (.Y(N1679), .A(N3635), .B(N3585));
NOR2XL inst_cellmath__43_0_I726 (.Y(N1681), .A(N3635), .B(N3586));
NOR2XL inst_cellmath__43_0_I727 (.Y(N1683), .A(N3635), .B(N3587));
NOR2XL inst_cellmath__43_0_I728 (.Y(N1685), .A(N3635), .B(N3588));
NOR2XL inst_cellmath__43_0_I729 (.Y(N1687), .A(N3635), .B(N3589));
NOR2XL inst_cellmath__43_0_I730 (.Y(N1689), .A(N3635), .B(N3590));
NOR2XL inst_cellmath__43_0_I731 (.Y(N1691), .A(N3635), .B(N3591));
NOR2XL inst_cellmath__43_0_I732 (.Y(N1693), .A(N3635), .B(N3592));
NOR2XL inst_cellmath__43_0_I733 (.Y(N1695), .A(N3635), .B(N3593));
NOR2XL inst_cellmath__43_0_I734 (.Y(N1697), .A(N3635), .B(N3594));
NOR2XL inst_cellmath__43_0_I735 (.Y(N1699), .A(N3635), .B(N3595));
NOR2XL inst_cellmath__43_0_I736 (.Y(N1701), .A(N3635), .B(N3596));
NOR2XL inst_cellmath__43_0_I737 (.Y(N1703), .A(N3635), .B(N3597));
NOR2XL inst_cellmath__43_0_I738 (.Y(N1705), .A(N3635), .B(N3598));
NOR2XL inst_cellmath__43_0_I739 (.Y(N1707), .A(N3635), .B(N3599));
NOR2XL inst_cellmath__43_0_I740 (.Y(N1709), .A(N3635), .B(N3600));
NOR2XL inst_cellmath__43_0_I741 (.Y(N1711), .A(N3635), .B(N3601));
NOR2XL inst_cellmath__43_0_I742 (.Y(N1713), .A(N3635), .B(N3602));
NOR2XL inst_cellmath__43_0_I743 (.Y(N1715), .A(N3635), .B(N3603));
NOR2XL inst_cellmath__43_0_I744 (.Y(N1717), .A(N3635), .B(N3604));
NOR2XL inst_cellmath__43_0_I745 (.Y(N1719), .A(N3635), .B(N3605));
NOR2XL inst_cellmath__43_0_I746 (.Y(N1721), .A(N3635), .B(N3606));
NOR2XL inst_cellmath__43_0_I747 (.Y(N1723), .A(N3635), .B(N3607));
INVXL inst_cellmath__43_0_I748 (.Y(N1725), .A(N3635));
INVXL inst_cellmath__43_0_I754 (.Y(N1734), .A(N3585));
INVXL inst_cellmath__43_0_I755 (.Y(N1736), .A(N3586));
INVXL inst_cellmath__43_0_I756 (.Y(N1738), .A(N3587));
INVXL inst_cellmath__43_0_I757 (.Y(N1740), .A(N3588));
INVXL inst_cellmath__43_0_I758 (.Y(N1742), .A(N3589));
INVXL inst_cellmath__43_0_I759 (.Y(N1744), .A(N3590));
INVXL inst_cellmath__43_0_I760 (.Y(N1746), .A(N3591));
INVXL inst_cellmath__43_0_I761 (.Y(N1748), .A(N3592));
INVXL inst_cellmath__43_0_I762 (.Y(N1750), .A(N3593));
INVXL inst_cellmath__43_0_I763 (.Y(N1752), .A(N3594));
INVXL inst_cellmath__43_0_I764 (.Y(N1754), .A(N3595));
INVXL inst_cellmath__43_0_I765 (.Y(N1756), .A(N3596));
INVXL inst_cellmath__43_0_I766 (.Y(N1758), .A(N3597));
INVXL inst_cellmath__43_0_I767 (.Y(N1760), .A(N3598));
INVXL inst_cellmath__43_0_I768 (.Y(N1762), .A(N3599));
INVXL inst_cellmath__43_0_I769 (.Y(N1764), .A(N3600));
INVXL inst_cellmath__43_0_I770 (.Y(N1766), .A(N3601));
INVXL inst_cellmath__43_0_I771 (.Y(N1768), .A(N3602));
INVXL inst_cellmath__43_0_I772 (.Y(N1770), .A(N3603));
INVXL inst_cellmath__43_0_I773 (.Y(N1772), .A(N3604));
INVXL inst_cellmath__43_0_I774 (.Y(N1774), .A(N3605));
INVXL inst_cellmath__43_0_I775 (.Y(N1776), .A(N3606));
INVXL inst_cellmath__43_0_I776 (.Y(N1778), .A(N3607));
ADDHX1 inst_cellmath__43_0_I807 (.CO(N1813), .S(N1812), .A(N385), .B(N442));
ADDHX1 inst_cellmath__43_0_I808 (.CO(N1815), .S(N1814), .A(N387), .B(N444));
ADDFX1 inst_cellmath__43_0_I809 (.CO(N1817), .S(N1816), .A(N501), .B(N558), .CI(N1813));
ADDHX1 inst_cellmath__43_0_I810 (.CO(N1819), .S(N1818), .A(N389), .B(N446));
ADDFX1 inst_cellmath__43_0_I811 (.CO(N1821), .S(N1820), .A(N560), .B(N503), .CI(N617));
ADDFX1 inst_cellmath__43_0_I812 (.CO(N1823), .S(N1822), .A(N1818), .B(N1815), .CI(N1817));
ADDHX1 inst_cellmath__43_0_I813 (.CO(N1825), .S(N1824), .A(N391), .B(N448));
ADDFX1 inst_cellmath__43_0_I814 (.CO(N1827), .S(N1826), .A(N562), .B(N505), .CI(N619));
ADDFX1 inst_cellmath__43_0_I815 (.CO(N1829), .S(N1828), .A(N1819), .B(N676), .CI(N1824));
ADDFX1 inst_cellmath__43_0_I816 (.CO(N1831), .S(N1830), .A(N1826), .B(N1821), .CI(N1828));
ADDHX1 inst_cellmath__43_0_I817 (.CO(N1833), .S(N1832), .A(N393), .B(N450));
ADDFX1 inst_cellmath__43_0_I818 (.CO(N1835), .S(N1834), .A(N564), .B(N507), .CI(N621));
ADDFX1 inst_cellmath__43_0_I819 (.CO(N1837), .S(N1836), .A(N735), .B(N678), .CI(N1825));
ADDFX1 inst_cellmath__43_0_I820 (.CO(N1839), .S(N1838), .A(N1827), .B(N1832), .CI(N1834));
ADDFX1 inst_cellmath__43_0_I821 (.CO(N1841), .S(N1840), .A(N1836), .B(N1829), .CI(N1838));
ADDHX1 inst_cellmath__43_0_I822 (.CO(N1843), .S(N1842), .A(N395), .B(N452));
ADDFX1 inst_cellmath__43_0_I823 (.CO(N1845), .S(N1844), .A(N566), .B(N509), .CI(N623));
ADDFX1 inst_cellmath__43_0_I824 (.CO(N1847), .S(N1846), .A(N737), .B(N680), .CI(N794));
ADDFX1 inst_cellmath__43_0_I825 (.CO(N1849), .S(N1848), .A(N1842), .B(N1833), .CI(N1835));
ADDFX1 inst_cellmath__43_0_I826 (.CO(N1851), .S(N1850), .A(N1844), .B(N1837), .CI(N1846));
ADDFX1 inst_cellmath__43_0_I827 (.CO(N1853), .S(N1852), .A(N1848), .B(N1839), .CI(N1850));
ADDHX1 inst_cellmath__43_0_I828 (.CO(N1855), .S(N1854), .A(N397), .B(N454));
ADDFX1 inst_cellmath__43_0_I829 (.CO(N1857), .S(N1856), .A(N568), .B(N511), .CI(N625));
ADDFX1 inst_cellmath__43_0_I830 (.CO(N1859), .S(N1858), .A(N739), .B(N682), .CI(N796));
ADDFX1 inst_cellmath__43_0_I831 (.CO(N1861), .S(N1860), .A(N1843), .B(N853), .CI(N1854));
ADDFX1 inst_cellmath__43_0_I832 (.CO(N1863), .S(N1862), .A(N1847), .B(N1845), .CI(N1856));
ADDFX1 inst_cellmath__43_0_I833 (.CO(N1865), .S(N1864), .A(N1849), .B(N1858), .CI(N1860));
ADDFX1 inst_cellmath__43_0_I834 (.CO(N1867), .S(N1866), .A(N1862), .B(N1851), .CI(N1864));
ADDHX1 inst_cellmath__43_0_I835 (.CO(N1869), .S(N1868), .A(N399), .B(N456));
ADDFX1 inst_cellmath__43_0_I836 (.CO(N1871), .S(N1870), .A(N570), .B(N513), .CI(N627));
ADDFX1 inst_cellmath__43_0_I837 (.CO(N1873), .S(N1872), .A(N741), .B(N684), .CI(N798));
ADDFX1 inst_cellmath__43_0_I838 (.CO(N1875), .S(N1874), .A(N912), .B(N855), .CI(N1855));
ADDFX1 inst_cellmath__43_0_I839 (.CO(N1877), .S(N1876), .A(N1857), .B(N1868), .CI(N1859));
ADDFX1 inst_cellmath__43_0_I840 (.CO(N1879), .S(N1878), .A(N1872), .B(N1870), .CI(N1861));
ADDFX1 inst_cellmath__43_0_I841 (.CO(N1881), .S(N1880), .A(N1863), .B(N1874), .CI(N1876));
ADDFX1 inst_cellmath__43_0_I842 (.CO(N1883), .S(N1882), .A(N1865), .B(N1878), .CI(N1880));
ADDHX1 inst_cellmath__43_0_I843 (.CO(N1885), .S(N1884), .A(N401), .B(N458));
ADDFX1 inst_cellmath__43_0_I844 (.CO(N1887), .S(N1886), .A(N572), .B(N515), .CI(N629));
ADDFX1 inst_cellmath__43_0_I845 (.CO(N1889), .S(N1888), .A(N743), .B(N686), .CI(N800));
ADDFX1 inst_cellmath__43_0_I846 (.CO(N1891), .S(N1890), .A(N914), .B(N857), .CI(N971));
ADDFX1 inst_cellmath__43_0_I847 (.CO(N1893), .S(N1892), .A(N1884), .B(N1869), .CI(N1871));
ADDFX1 inst_cellmath__43_0_I848 (.CO(N1895), .S(N1894), .A(N1875), .B(N1873), .CI(N1886));
ADDFX1 inst_cellmath__43_0_I849 (.CO(N1897), .S(N1896), .A(N1890), .B(N1888), .CI(N1877));
ADDFX1 inst_cellmath__43_0_I850 (.CO(N1899), .S(N1898), .A(N1879), .B(N1892), .CI(N1894));
ADDFX1 inst_cellmath__43_0_I851 (.CO(N1901), .S(N1900), .A(N1881), .B(N1896), .CI(N1898));
ADDHX1 inst_cellmath__43_0_I852 (.CO(N1903), .S(N1902), .A(N403), .B(N460));
ADDFX1 inst_cellmath__43_0_I853 (.CO(N1905), .S(N1904), .A(N574), .B(N517), .CI(N631));
ADDFX1 inst_cellmath__43_0_I854 (.CO(N1907), .S(N1906), .A(N745), .B(N688), .CI(N802));
ADDFX1 inst_cellmath__43_0_I855 (.CO(N1909), .S(N1908), .A(N916), .B(N859), .CI(N973));
ADDFX1 inst_cellmath__43_0_I856 (.CO(N1911), .S(N1910), .A(N1885), .B(N1030), .CI(N1902));
ADDFX1 inst_cellmath__43_0_I857 (.CO(N1913), .S(N1912), .A(N1889), .B(N1887), .CI(N1891));
ADDFX1 inst_cellmath__43_0_I858 (.CO(N1915), .S(N1914), .A(N1906), .B(N1904), .CI(N1908));
ADDFX1 inst_cellmath__43_0_I859 (.CO(N1917), .S(N1916), .A(N1910), .B(N1893), .CI(N1895));
ADDFX1 inst_cellmath__43_0_I860 (.CO(N1919), .S(N1918), .A(N1897), .B(N1912), .CI(N1914));
ADDFX1 inst_cellmath__43_0_I861 (.CO(N1921), .S(N1920), .A(N1899), .B(N1916), .CI(N1918));
ADDHX1 inst_cellmath__43_0_I862 (.CO(N1923), .S(N1922), .A(N405), .B(N462));
ADDFX1 inst_cellmath__43_0_I863 (.CO(N1925), .S(N1924), .A(N576), .B(N519), .CI(N633));
ADDFX1 inst_cellmath__43_0_I864 (.CO(N1927), .S(N1926), .A(N747), .B(N690), .CI(N804));
ADDFX1 inst_cellmath__43_0_I865 (.CO(N1929), .S(N1928), .A(N918), .B(N861), .CI(N975));
ADDFX1 inst_cellmath__43_0_I866 (.CO(N1931), .S(N1930), .A(N1089), .B(N1032), .CI(N1903));
ADDFX1 inst_cellmath__43_0_I867 (.CO(N1933), .S(N1932), .A(N1905), .B(N1922), .CI(N1907));
ADDFX1 inst_cellmath__43_0_I868 (.CO(N1935), .S(N1934), .A(N1924), .B(N1909), .CI(N1926));
ADDFX1 inst_cellmath__43_0_I869 (.CO(N1937), .S(N1936), .A(N1911), .B(N1928), .CI(N1930));
ADDFX1 inst_cellmath__43_0_I870 (.CO(N1939), .S(N1938), .A(N1915), .B(N1913), .CI(N1932));
ADDFX1 inst_cellmath__43_0_I871 (.CO(N1941), .S(N1940), .A(N1917), .B(N1934), .CI(N1936));
ADDFX1 inst_cellmath__43_0_I872 (.CO(N1943), .S(N1942), .A(N1938), .B(N1919), .CI(N1940));
ADDHX1 inst_cellmath__43_0_I873 (.CO(N1945), .S(N1944), .A(N407), .B(N464));
ADDFX1 inst_cellmath__43_0_I874 (.CO(N1947), .S(N1946), .A(N578), .B(N521), .CI(N635));
ADDFX1 inst_cellmath__43_0_I875 (.CO(N1949), .S(N1948), .A(N749), .B(N692), .CI(N806));
ADDFX1 inst_cellmath__43_0_I876 (.CO(N1951), .S(N1950), .A(N920), .B(N863), .CI(N977));
ADDFX1 inst_cellmath__43_0_I877 (.CO(N1953), .S(N1952), .A(N1091), .B(N1034), .CI(N1148));
ADDFX1 inst_cellmath__43_0_I878 (.CO(N1955), .S(N1954), .A(N1944), .B(N1923), .CI(N1925));
ADDFX1 inst_cellmath__43_0_I879 (.CO(N1957), .S(N1956), .A(N1929), .B(N1927), .CI(N1931));
ADDFX1 inst_cellmath__43_0_I880 (.CO(N1959), .S(N1958), .A(N1948), .B(N1946), .CI(N1950));
ADDFX1 inst_cellmath__43_0_I881 (.CO(N1961), .S(N1960), .A(N1933), .B(N1952), .CI(N1954));
ADDFX1 inst_cellmath__43_0_I882 (.CO(N1963), .S(N1962), .A(N1937), .B(N1935), .CI(N1956));
ADDFX1 inst_cellmath__43_0_I883 (.CO(N1965), .S(N1964), .A(N1939), .B(N1958), .CI(N1960));
ADDFX1 inst_cellmath__43_0_I884 (.CO(N1967), .S(N1966), .A(N1941), .B(N1962), .CI(N1964));
ADDHX1 inst_cellmath__43_0_I885 (.CO(N1969), .S(N1968), .A(N409), .B(N466));
ADDFX1 inst_cellmath__43_0_I886 (.CO(N1971), .S(N1970), .A(N580), .B(N523), .CI(N637));
ADDFX1 inst_cellmath__43_0_I887 (.CO(N1973), .S(N1972), .A(N751), .B(N694), .CI(N808));
ADDFX1 inst_cellmath__43_0_I888 (.CO(N1975), .S(N1974), .A(N922), .B(N865), .CI(N979));
ADDFX1 inst_cellmath__43_0_I889 (.CO(N1977), .S(N1976), .A(N1093), .B(N1036), .CI(N1150));
ADDFX1 inst_cellmath__43_0_I890 (.CO(N1979), .S(N1978), .A(N1945), .B(N1207), .CI(N1968));
ADDFX1 inst_cellmath__43_0_I891 (.CO(N1981), .S(N1980), .A(N1949), .B(N1947), .CI(N1951));
ADDFX1 inst_cellmath__43_0_I892 (.CO(N1983), .S(N1982), .A(N1970), .B(N1953), .CI(N1972));
ADDFX1 inst_cellmath__43_0_I893 (.CO(N1985), .S(N1984), .A(N1976), .B(N1974), .CI(N1955));
ADDFX1 inst_cellmath__43_0_I894 (.CO(N1987), .S(N1986), .A(N1957), .B(N1978), .CI(N1959));
ADDFX1 inst_cellmath__43_0_I895 (.CO(N1989), .S(N1988), .A(N1982), .B(N1980), .CI(N1984));
ADDFX1 inst_cellmath__43_0_I896 (.CO(N1991), .S(N1990), .A(N1963), .B(N1961), .CI(N1986));
ADDFX1 inst_cellmath__43_0_I897 (.CO(N1993), .S(N1992), .A(N1965), .B(N1988), .CI(N1990));
ADDHX1 inst_cellmath__43_0_I898 (.CO(N1995), .S(N1994), .A(N411), .B(N468));
ADDFX1 inst_cellmath__43_0_I899 (.CO(N1997), .S(N1996), .A(N582), .B(N525), .CI(N639));
ADDFX1 inst_cellmath__43_0_I900 (.CO(N1999), .S(N1998), .A(N753), .B(N696), .CI(N810));
ADDFX1 inst_cellmath__43_0_I901 (.CO(N2001), .S(N2000), .A(N924), .B(N867), .CI(N981));
ADDFX1 inst_cellmath__43_0_I902 (.CO(N2003), .S(N2002), .A(N1095), .B(N1038), .CI(N1152));
ADDFX1 inst_cellmath__43_0_I903 (.CO(N2005), .S(N2004), .A(N1266), .B(N1209), .CI(N1969));
ADDFX1 inst_cellmath__43_0_I904 (.CO(N2007), .S(N2006), .A(N1971), .B(N1994), .CI(N1973));
ADDFX1 inst_cellmath__43_0_I905 (.CO(N2009), .S(N2008), .A(N1977), .B(N1975), .CI(N1996));
ADDFX1 inst_cellmath__43_0_I906 (.CO(N2011), .S(N2010), .A(N2000), .B(N1998), .CI(N2002));
ADDFX1 inst_cellmath__43_0_I907 (.CO(N2013), .S(N2012), .A(N2004), .B(N1979), .CI(N1981));
ADDFX1 inst_cellmath__43_0_I908 (.CO(N2015), .S(N2014), .A(N2006), .B(N1983), .CI(N1985));
ADDFX1 inst_cellmath__43_0_I909 (.CO(N2017), .S(N2016), .A(N2010), .B(N2008), .CI(N1987));
ADDFX1 inst_cellmath__43_0_I910 (.CO(N2019), .S(N2018), .A(N2014), .B(N2012), .CI(N1989));
ADDFX1 inst_cellmath__43_0_I911 (.CO(N2021), .S(N2020), .A(N1991), .B(N2016), .CI(N2018));
ADDHX1 inst_cellmath__43_0_I912 (.CO(N2023), .S(N2022), .A(N413), .B(N470));
ADDFX1 inst_cellmath__43_0_I913 (.CO(N2025), .S(N2024), .A(N584), .B(N527), .CI(N641));
ADDFX1 inst_cellmath__43_0_I914 (.CO(N2027), .S(N2026), .A(N755), .B(N698), .CI(N812));
ADDFX1 inst_cellmath__43_0_I915 (.CO(N2029), .S(N2028), .A(N926), .B(N869), .CI(N983));
ADDFX1 inst_cellmath__43_0_I916 (.CO(N2031), .S(N2030), .A(N1097), .B(N1040), .CI(N1154));
ADDFX1 inst_cellmath__43_0_I917 (.CO(N2033), .S(N2032), .A(N1268), .B(N1211), .CI(N1325));
ADDFX1 inst_cellmath__43_0_I918 (.CO(N2035), .S(N2034), .A(N2022), .B(N1995), .CI(N1997));
ADDFX1 inst_cellmath__43_0_I919 (.CO(N2037), .S(N2036), .A(N2001), .B(N1999), .CI(N2003));
ADDFX1 inst_cellmath__43_0_I920 (.CO(N2039), .S(N2038), .A(N2024), .B(N2005), .CI(N2026));
ADDFX1 inst_cellmath__43_0_I921 (.CO(N2041), .S(N2040), .A(N2030), .B(N2028), .CI(N2032));
ADDFX1 inst_cellmath__43_0_I922 (.CO(N2043), .S(N2042), .A(N2009), .B(N2007), .CI(N2011));
ADDFX1 inst_cellmath__43_0_I923 (.CO(N2045), .S(N2044), .A(N2036), .B(N2034), .CI(N2013));
ADDFX1 inst_cellmath__43_0_I924 (.CO(N2047), .S(N2046), .A(N2040), .B(N2038), .CI(N2015));
ADDFX1 inst_cellmath__43_0_I925 (.CO(N2049), .S(N2048), .A(N2017), .B(N2042), .CI(N2044));
ADDFX1 inst_cellmath__43_0_I926 (.CO(N2051), .S(N2050), .A(N2019), .B(N2046), .CI(N2048));
ADDHX1 inst_cellmath__43_0_I927 (.CO(N2053), .S(N2052), .A(N415), .B(N472));
ADDFX1 inst_cellmath__43_0_I928 (.CO(N2055), .S(N2054), .A(N586), .B(N529), .CI(N643));
ADDFX1 inst_cellmath__43_0_I929 (.CO(N2057), .S(N2056), .A(N757), .B(N700), .CI(N814));
ADDFX1 inst_cellmath__43_0_I930 (.CO(N2059), .S(N2058), .A(N928), .B(N871), .CI(N985));
ADDFX1 inst_cellmath__43_0_I931 (.CO(N2061), .S(N2060), .A(N1099), .B(N1042), .CI(N1156));
ADDFX1 inst_cellmath__43_0_I932 (.CO(N2063), .S(N2062), .A(N1270), .B(N1213), .CI(N1327));
ADDFX1 inst_cellmath__43_0_I933 (.CO(N2065), .S(N2064), .A(N2023), .B(N1384), .CI(N2052));
ADDFX1 inst_cellmath__43_0_I934 (.CO(N2067), .S(N2066), .A(N2027), .B(N2025), .CI(N2029));
ADDFX1 inst_cellmath__43_0_I935 (.CO(N2069), .S(N2068), .A(N2033), .B(N2031), .CI(N2054));
ADDFX1 inst_cellmath__43_0_I936 (.CO(N2071), .S(N2070), .A(N2058), .B(N2056), .CI(N2060));
ADDFX1 inst_cellmath__43_0_I937 (.CO(N2073), .S(N2072), .A(N2035), .B(N2062), .CI(N2037));
ADDFX1 inst_cellmath__43_0_I938 (.CO(N2075), .S(N2074), .A(N2039), .B(N2064), .CI(N2066));
ADDFX1 inst_cellmath__43_0_I939 (.CO(N2077), .S(N2076), .A(N2068), .B(N2041), .CI(N2070));
ADDFX1 inst_cellmath__43_0_I940 (.CO(N2079), .S(N2078), .A(N2072), .B(N2043), .CI(N2045));
ADDFX1 inst_cellmath__43_0_I941 (.CO(N2081), .S(N2080), .A(N2076), .B(N2074), .CI(N2047));
ADDFX1 inst_cellmath__43_0_I942 (.CO(N2083), .S(N2082), .A(N2049), .B(N2078), .CI(N2080));
ADDHX1 inst_cellmath__43_0_I943 (.CO(N2085), .S(N2084), .A(N417), .B(N474));
ADDFX1 inst_cellmath__43_0_I944 (.CO(N2087), .S(N2086), .A(N588), .B(N531), .CI(N645));
ADDFX1 inst_cellmath__43_0_I945 (.CO(N2089), .S(N2088), .A(N759), .B(N702), .CI(N816));
ADDFX1 inst_cellmath__43_0_I946 (.CO(N2091), .S(N2090), .A(N930), .B(N873), .CI(N987));
ADDFX1 inst_cellmath__43_0_I947 (.CO(N2093), .S(N2092), .A(N1101), .B(N1044), .CI(N1158));
ADDFX1 inst_cellmath__43_0_I948 (.CO(N2095), .S(N2094), .A(N1272), .B(N1215), .CI(N1329));
ADDFX1 inst_cellmath__43_0_I949 (.CO(N2097), .S(N2096), .A(N1443), .B(N1386), .CI(N2053));
ADDFX1 inst_cellmath__43_0_I950 (.CO(N2099), .S(N2098), .A(N2055), .B(N2084), .CI(N2057));
ADDFX1 inst_cellmath__43_0_I951 (.CO(N2101), .S(N2100), .A(N2061), .B(N2059), .CI(N2063));
ADDFX1 inst_cellmath__43_0_I952 (.CO(N2103), .S(N2102), .A(N2088), .B(N2086), .CI(N2090));
ADDFX1 inst_cellmath__43_0_I953 (.CO(N2105), .S(N2104), .A(N2094), .B(N2092), .CI(N2065));
ADDFX1 inst_cellmath__43_0_I954 (.CO(N2107), .S(N2106), .A(N2067), .B(N2096), .CI(N2069));
ADDFX1 inst_cellmath__43_0_I955 (.CO(N2109), .S(N2108), .A(N2098), .B(N2071), .CI(N2100));
ADDFX1 inst_cellmath__43_0_I956 (.CO(N2111), .S(N2110), .A(N2102), .B(N2073), .CI(N2104));
ADDFX1 inst_cellmath__43_0_I957 (.CO(N2113), .S(N2112), .A(N2106), .B(N2075), .CI(N2077));
ADDFX1 inst_cellmath__43_0_I958 (.CO(N2115), .S(N2114), .A(N2110), .B(N2108), .CI(N2079));
ADDFX1 inst_cellmath__43_0_I959 (.CO(N2117), .S(N2116), .A(N2081), .B(N2112), .CI(N2114));
ADDHX1 inst_cellmath__43_0_I960 (.CO(N2119), .S(N2118), .A(N419), .B(N476));
ADDFX1 inst_cellmath__43_0_I961 (.CO(N2121), .S(N2120), .A(N590), .B(N533), .CI(N647));
ADDFX1 inst_cellmath__43_0_I962 (.CO(N2123), .S(N2122), .A(N761), .B(N704), .CI(N818));
ADDFX1 inst_cellmath__43_0_I963 (.CO(N2125), .S(N2124), .A(N932), .B(N875), .CI(N989));
ADDFX1 inst_cellmath__43_0_I964 (.CO(N2127), .S(N2126), .A(N1103), .B(N1046), .CI(N1160));
ADDFX1 inst_cellmath__43_0_I965 (.CO(N2129), .S(N2128), .A(N1274), .B(N1217), .CI(N1331));
ADDFX1 inst_cellmath__43_0_I966 (.CO(N2131), .S(N2130), .A(N1445), .B(N1388), .CI(N1502));
ADDFX1 inst_cellmath__43_0_I967 (.CO(N2133), .S(N2132), .A(N2118), .B(N2085), .CI(N2087));
ADDFX1 inst_cellmath__43_0_I968 (.CO(N2135), .S(N2134), .A(N2091), .B(N2089), .CI(N2093));
ADDFX1 inst_cellmath__43_0_I969 (.CO(N2137), .S(N2136), .A(N2097), .B(N2095), .CI(N2120));
ADDFX1 inst_cellmath__43_0_I970 (.CO(N2139), .S(N2138), .A(N2124), .B(N2122), .CI(N2126));
ADDFX1 inst_cellmath__43_0_I971 (.CO(N2141), .S(N2140), .A(N2130), .B(N2128), .CI(N2099));
ADDFX1 inst_cellmath__43_0_I972 (.CO(N2143), .S(N2142), .A(N2132), .B(N2101), .CI(N2103));
ADDFX1 inst_cellmath__43_0_I973 (.CO(N2145), .S(N2144), .A(N2105), .B(N2134), .CI(N2136));
ADDFX1 inst_cellmath__43_0_I974 (.CO(N2147), .S(N2146), .A(N2107), .B(N2138), .CI(N2140));
ADDFX1 inst_cellmath__43_0_I975 (.CO(N2149), .S(N2148), .A(N2142), .B(N2109), .CI(N2111));
ADDFX1 inst_cellmath__43_0_I976 (.CO(N2151), .S(N2150), .A(N2146), .B(N2144), .CI(N2113));
ADDFX1 inst_cellmath__43_0_I977 (.CO(N2153), .S(N2152), .A(N2115), .B(N2148), .CI(N2150));
ADDHX1 inst_cellmath__43_0_I978 (.CO(N2155), .S(N2154), .A(N421), .B(N478));
ADDFX1 inst_cellmath__43_0_I979 (.CO(N2157), .S(N2156), .A(N592), .B(N535), .CI(N649));
ADDFX1 inst_cellmath__43_0_I980 (.CO(N2159), .S(N2158), .A(N763), .B(N706), .CI(N820));
ADDFX1 inst_cellmath__43_0_I981 (.CO(N2161), .S(N2160), .A(N934), .B(N877), .CI(N991));
ADDFX1 inst_cellmath__43_0_I982 (.CO(N2163), .S(N2162), .A(N1105), .B(N1048), .CI(N1162));
ADDFX1 inst_cellmath__43_0_I983 (.CO(N2165), .S(N2164), .A(N1276), .B(N1219), .CI(N1333));
ADDFX1 inst_cellmath__43_0_I984 (.CO(N2167), .S(N2166), .A(N1447), .B(N1390), .CI(N1504));
ADDFX1 inst_cellmath__43_0_I985 (.CO(N2169), .S(N2168), .A(N2119), .B(N1561), .CI(N2154));
ADDFX1 inst_cellmath__43_0_I986 (.CO(N2171), .S(N2170), .A(N2123), .B(N2121), .CI(N2125));
ADDFX1 inst_cellmath__43_0_I987 (.CO(N2173), .S(N2172), .A(N2129), .B(N2127), .CI(N2131));
ADDFX1 inst_cellmath__43_0_I988 (.CO(N2175), .S(N2174), .A(N2158), .B(N2156), .CI(N2160));
ADDFX1 inst_cellmath__43_0_I989 (.CO(N2177), .S(N2176), .A(N2164), .B(N2162), .CI(N2166));
ADDFX1 inst_cellmath__43_0_I990 (.CO(N2179), .S(N2178), .A(N2135), .B(N2133), .CI(N2168));
ADDFX1 inst_cellmath__43_0_I991 (.CO(N2181), .S(N2180), .A(N2170), .B(N2137), .CI(N2172));
ADDFX1 inst_cellmath__43_0_I992 (.CO(N2183), .S(N2182), .A(N2141), .B(N2139), .CI(N2174));
ADDFX1 inst_cellmath__43_0_I993 (.CO(N2185), .S(N2184), .A(N2143), .B(N2176), .CI(N2178));
ADDFX1 inst_cellmath__43_0_I994 (.CO(N2187), .S(N2186), .A(N2180), .B(N2145), .CI(N2147));
ADDFX1 inst_cellmath__43_0_I995 (.CO(N2189), .S(N2188), .A(N2149), .B(N2182), .CI(N2184));
ADDFX1 inst_cellmath__43_0_I996 (.CO(N2191), .S(N2190), .A(N2151), .B(N2186), .CI(N2188));
ADDHX1 inst_cellmath__43_0_I997 (.CO(N2193), .S(N2192), .A(N423), .B(N480));
ADDFX1 inst_cellmath__43_0_I998 (.CO(N2195), .S(N2194), .A(N594), .B(N537), .CI(N651));
ADDFX1 inst_cellmath__43_0_I999 (.CO(N2197), .S(N2196), .A(N765), .B(N708), .CI(N822));
ADDFX1 inst_cellmath__43_0_I1000 (.CO(N2199), .S(N2198), .A(N936), .B(N879), .CI(N993));
ADDFX1 inst_cellmath__43_0_I1001 (.CO(N2201), .S(N2200), .A(N1107), .B(N1050), .CI(N1164));
ADDFX1 inst_cellmath__43_0_I1002 (.CO(N2203), .S(N2202), .A(N1278), .B(N1221), .CI(N1335));
ADDFX1 inst_cellmath__43_0_I1003 (.CO(N2205), .S(N2204), .A(N1449), .B(N1392), .CI(N1506));
ADDFX1 inst_cellmath__43_0_I1004 (.CO(N2207), .S(N2206), .A(N1620), .B(N1563), .CI(N2155));
ADDFX1 inst_cellmath__43_0_I1005 (.CO(N2209), .S(N2208), .A(N2157), .B(N2192), .CI(N2159));
ADDFX1 inst_cellmath__43_0_I1006 (.CO(N2211), .S(N2210), .A(N2163), .B(N2161), .CI(N2165));
ADDFX1 inst_cellmath__43_0_I1007 (.CO(N2213), .S(N2212), .A(N2194), .B(N2167), .CI(N2196));
ADDFX1 inst_cellmath__43_0_I1008 (.CO(N2215), .S(N2214), .A(N2200), .B(N2198), .CI(N2202));
ADDFX1 inst_cellmath__43_0_I1009 (.CO(N2217), .S(N2216), .A(N2169), .B(N2204), .CI(N2206));
ADDFX1 inst_cellmath__43_0_I1010 (.CO(N2219), .S(N2218), .A(N2173), .B(N2171), .CI(N2175));
ADDFX1 inst_cellmath__43_0_I1011 (.CO(N2221), .S(N2220), .A(N2208), .B(N2177), .CI(N2210));
ADDFX1 inst_cellmath__43_0_I1012 (.CO(N2223), .S(N2222), .A(N2214), .B(N2212), .CI(N2179));
ADDFX1 inst_cellmath__43_0_I1013 (.CO(N2225), .S(N2224), .A(N2181), .B(N2216), .CI(N2218));
ADDFX1 inst_cellmath__43_0_I1014 (.CO(N2227), .S(N2226), .A(N2220), .B(N2183), .CI(N2185));
ADDFX1 inst_cellmath__43_0_I1015 (.CO(N2229), .S(N2228), .A(N2187), .B(N2222), .CI(N2224));
ADDFX1 inst_cellmath__43_0_I1016 (.CO(N2231), .S(N2230), .A(N2189), .B(N2226), .CI(N2228));
XNOR2X1 hap1_A_I1927 (.Y(N2232), .A(N425), .B(N482));
OR2XL hap1_A_I1928 (.Y(N2233), .A(N425), .B(N482));
ADDFX1 inst_cellmath__43_0_I1018 (.CO(N2237), .S(N2236), .A(N596), .B(N539), .CI(N653));
ADDFX1 inst_cellmath__43_0_I1019 (.CO(N2239), .S(N2238), .A(N767), .B(N710), .CI(N824));
ADDFX1 inst_cellmath__43_0_I1020 (.CO(N2241), .S(N2240), .A(N938), .B(N881), .CI(N995));
ADDFX1 inst_cellmath__43_0_I1021 (.CO(N2243), .S(N2242), .A(N1109), .B(N1052), .CI(N1166));
ADDFX1 inst_cellmath__43_0_I1022 (.CO(N2245), .S(N2244), .A(N1280), .B(N1223), .CI(N1337));
ADDFX1 inst_cellmath__43_0_I1023 (.CO(N2247), .S(N2246), .A(N1451), .B(N1394), .CI(N1508));
ADDFX1 inst_cellmath__43_0_I1024 (.CO(N2249), .S(N2248), .A(N1622), .B(N1565), .CI(N1679));
ADDFX1 inst_cellmath__43_0_I1025 (.CO(N2251), .S(N2250), .A(N2232), .B(N2193), .CI(N2195));
ADDFX1 inst_cellmath__43_0_I1026 (.CO(N2253), .S(N2252), .A(N2199), .B(N2197), .CI(N2201));
ADDFX1 inst_cellmath__43_0_I1027 (.CO(N2255), .S(N2254), .A(N2205), .B(N2203), .CI(N2207));
ADDFX1 inst_cellmath__43_0_I1028 (.CO(N2257), .S(N2256), .A(N2238), .B(N2236), .CI(N2240));
ADDFX1 inst_cellmath__43_0_I1029 (.CO(N2259), .S(N2258), .A(N2244), .B(N2242), .CI(N2246));
ADDFX1 inst_cellmath__43_0_I1030 (.CO(N2261), .S(N2260), .A(N2209), .B(N2248), .CI(N2211));
ADDFX1 inst_cellmath__43_0_I1031 (.CO(N2263), .S(N2262), .A(N2213), .B(N2250), .CI(N2252));
ADDFX1 inst_cellmath__43_0_I1032 (.CO(N2265), .S(N2264), .A(N2217), .B(N2215), .CI(N2254));
ADDFX1 inst_cellmath__43_0_I1033 (.CO(N2267), .S(N2266), .A(N2258), .B(N2256), .CI(N2219));
ADDFX1 inst_cellmath__43_0_I1034 (.CO(N2269), .S(N2268), .A(N2260), .B(N2221), .CI(N2262));
ADDFX1 inst_cellmath__43_0_I1035 (.CO(N2271), .S(N2270), .A(N2264), .B(N2223), .CI(N2266));
ADDFX1 inst_cellmath__43_0_I1036 (.CO(N2273), .S(N2272), .A(N2268), .B(N2225), .CI(N2227));
ADDFX1 inst_cellmath__43_0_I1037 (.CO(N2275), .S(N2274), .A(N2229), .B(N2270), .CI(N2272));
ADDHX1 inst_cellmath__43_0_I1038 (.CO(N2277), .S(N2276), .A(N1734), .B(N484));
ADDFX1 inst_cellmath__43_0_I1039 (.CO(N2279), .S(N2278), .A(N541), .B(N427), .CI(N598));
ADDFX1 inst_cellmath__43_0_I1040 (.CO(N2281), .S(N2280), .A(N712), .B(N655), .CI(N769));
ADDFX1 inst_cellmath__43_0_I1041 (.CO(N2283), .S(N2282), .A(N883), .B(N826), .CI(N940));
ADDFX1 inst_cellmath__43_0_I1042 (.CO(N2285), .S(N2284), .A(N1054), .B(N997), .CI(N1111));
ADDFX1 inst_cellmath__43_0_I1043 (.CO(N2287), .S(N2286), .A(N1225), .B(N1168), .CI(N1282));
ADDFX1 inst_cellmath__43_0_I1044 (.CO(N2289), .S(N2288), .A(N1396), .B(N1339), .CI(N1453));
ADDFX1 inst_cellmath__43_0_I1045 (.CO(N2291), .S(N2290), .A(N1567), .B(N1510), .CI(N1624));
ADDFX1 inst_cellmath__43_0_I1046 (.CO(N2293), .S(N2292), .A(N2233), .B(N1681), .CI(N2276));
ADDFX1 inst_cellmath__43_0_I1047 (.CO(N2295), .S(N2294), .A(N2239), .B(N2237), .CI(N2241));
ADDFX1 inst_cellmath__43_0_I1048 (.CO(N2297), .S(N2296), .A(N2245), .B(N2243), .CI(N2247));
ADDFX1 inst_cellmath__43_0_I1049 (.CO(N2299), .S(N2298), .A(N2278), .B(N2249), .CI(N2280));
ADDFX1 inst_cellmath__43_0_I1050 (.CO(N2301), .S(N2300), .A(N2284), .B(N2282), .CI(N2286));
ADDFX1 inst_cellmath__43_0_I1051 (.CO(N2303), .S(N2302), .A(N2290), .B(N2288), .CI(N2251));
ADDFX1 inst_cellmath__43_0_I1052 (.CO(N2305), .S(N2304), .A(N2292), .B(N2253), .CI(N2255));
ADDFX1 inst_cellmath__43_0_I1053 (.CO(N2307), .S(N2306), .A(N2294), .B(N2257), .CI(N2296));
ADDFX1 inst_cellmath__43_0_I1054 (.CO(N2309), .S(N2308), .A(N2298), .B(N2259), .CI(N2300));
ADDFX1 inst_cellmath__43_0_I1055 (.CO(N2311), .S(N2310), .A(N2302), .B(N2261), .CI(N2263));
ADDFX1 inst_cellmath__43_0_I1056 (.CO(N2313), .S(N2312), .A(N2265), .B(N2304), .CI(N2306));
ADDFX1 inst_cellmath__43_0_I1057 (.CO(N2315), .S(N2314), .A(N2308), .B(N2267), .CI(N2310));
ADDFX1 inst_cellmath__43_0_I1058 (.CO(N2317), .S(N2316), .A(N2312), .B(N2269), .CI(N2271));
ADDFX1 inst_cellmath__43_0_I1059 (.CO(N2319), .S(N2318), .A(N2273), .B(N2314), .CI(N2316));
ADDHX1 inst_cellmath__43_0_I1060 (.CO(N2321), .S(N2320), .A(N1736), .B(N543));
ADDFX1 inst_cellmath__43_0_I1061 (.CO(N2323), .S(N2322), .A(N600), .B(N486), .CI(N657));
ADDFX1 inst_cellmath__43_0_I1062 (.CO(N2325), .S(N2324), .A(N771), .B(N714), .CI(N828));
ADDFX1 inst_cellmath__43_0_I1063 (.CO(N2327), .S(N2326), .A(N942), .B(N885), .CI(N999));
ADDFX1 inst_cellmath__43_0_I1064 (.CO(N2329), .S(N2328), .A(N1113), .B(N1056), .CI(N1170));
ADDFX1 inst_cellmath__43_0_I1065 (.CO(N2331), .S(N2330), .A(N1284), .B(N1227), .CI(N1341));
ADDFX1 inst_cellmath__43_0_I1066 (.CO(N2333), .S(N2332), .A(N1455), .B(N1398), .CI(N1512));
ADDFX1 inst_cellmath__43_0_I1067 (.CO(N2335), .S(N2334), .A(N1626), .B(N1569), .CI(N1683));
ADDFX1 inst_cellmath__43_0_I1068 (.CO(N2337), .S(N2336), .A(N2320), .B(N2277), .CI(N2279));
ADDFX1 inst_cellmath__43_0_I1069 (.CO(N2339), .S(N2338), .A(N2283), .B(N2281), .CI(N2285));
ADDFX1 inst_cellmath__43_0_I1070 (.CO(N2341), .S(N2340), .A(N2289), .B(N2287), .CI(N2291));
ADDFX1 inst_cellmath__43_0_I1071 (.CO(N2343), .S(N2342), .A(N2324), .B(N2322), .CI(N2326));
ADDFX1 inst_cellmath__43_0_I1072 (.CO(N2345), .S(N2344), .A(N2330), .B(N2328), .CI(N2332));
ADDFX1 inst_cellmath__43_0_I1073 (.CO(N2347), .S(N2346), .A(N2293), .B(N2334), .CI(N2295));
ADDFX1 inst_cellmath__43_0_I1074 (.CO(N2349), .S(N2348), .A(N2336), .B(N2297), .CI(N2299));
ADDFX1 inst_cellmath__43_0_I1075 (.CO(N2351), .S(N2350), .A(N2338), .B(N2301), .CI(N2340));
ADDFX1 inst_cellmath__43_0_I1076 (.CO(N2353), .S(N2352), .A(N2342), .B(N2303), .CI(N2344));
ADDFX1 inst_cellmath__43_0_I1077 (.CO(N2355), .S(N2354), .A(N2346), .B(N2305), .CI(N2307));
ADDFX1 inst_cellmath__43_0_I1078 (.CO(N2357), .S(N2356), .A(N2350), .B(N2348), .CI(N2309));
ADDFX1 inst_cellmath__43_0_I1079 (.CO(N2359), .S(N2358), .A(N2352), .B(N2311), .CI(N2313));
ADDFX1 inst_cellmath__43_0_I1080 (.CO(N2361), .S(N2360), .A(N2356), .B(N2354), .CI(N2315));
ADDFX1 inst_cellmath__43_0_I1081 (.CO(N2363), .S(N2362), .A(N2317), .B(N2358), .CI(N2360));
ADDFX1 inst_cellmath__43_0_I1082 (.CO(N2365), .S(N2364), .A(N602), .B(N1738), .CI(N659));
ADDFX1 inst_cellmath__43_0_I1083 (.CO(N2367), .S(N2366), .A(N716), .B(N545), .CI(N773));
ADDFX1 inst_cellmath__43_0_I1084 (.CO(N2369), .S(N2368), .A(N887), .B(N830), .CI(N944));
ADDFX1 inst_cellmath__43_0_I1085 (.CO(N2371), .S(N2370), .A(N1058), .B(N1001), .CI(N1115));
ADDFX1 inst_cellmath__43_0_I1086 (.CO(N2373), .S(N2372), .A(N1229), .B(N1172), .CI(N1286));
ADDFX1 inst_cellmath__43_0_I1087 (.CO(N2375), .S(N2374), .A(N1400), .B(N1343), .CI(N1457));
ADDFX1 inst_cellmath__43_0_I1088 (.CO(N2377), .S(N2376), .A(N1571), .B(N1514), .CI(N1628));
ADDFX1 inst_cellmath__43_0_I1089 (.CO(N2379), .S(N2378), .A(N2321), .B(N1685), .CI(N2323));
ADDFX1 inst_cellmath__43_0_I1090 (.CO(N2381), .S(N2380), .A(N2327), .B(N2325), .CI(N2329));
ADDFX1 inst_cellmath__43_0_I1091 (.CO(N2383), .S(N2382), .A(N2333), .B(N2331), .CI(N2335));
ADDFX1 inst_cellmath__43_0_I1092 (.CO(N2385), .S(N2384), .A(N2366), .B(N2364), .CI(N2368));
ADDFX1 inst_cellmath__43_0_I1093 (.CO(N2387), .S(N2386), .A(N2372), .B(N2370), .CI(N2374));
ADDFX1 inst_cellmath__43_0_I1094 (.CO(N2389), .S(N2388), .A(N2337), .B(N2376), .CI(N2339));
ADDFX1 inst_cellmath__43_0_I1095 (.CO(N2391), .S(N2390), .A(N2378), .B(N2341), .CI(N2343));
ADDFX1 inst_cellmath__43_0_I1096 (.CO(N2393), .S(N2392), .A(N2380), .B(N2345), .CI(N2382));
ADDFX1 inst_cellmath__43_0_I1097 (.CO(N2395), .S(N2394), .A(N2384), .B(N2347), .CI(N2386));
ADDFX1 inst_cellmath__43_0_I1098 (.CO(N2397), .S(N2396), .A(N2388), .B(N2349), .CI(N2351));
ADDFX1 inst_cellmath__43_0_I1099 (.CO(N2399), .S(N2398), .A(N2392), .B(N2390), .CI(N2353));
ADDFX1 inst_cellmath__43_0_I1100 (.CO(N2401), .S(N2400), .A(N2394), .B(N2355), .CI(N2396));
ADDFX1 inst_cellmath__43_0_I1101 (.CO(N2403), .S(N2402), .A(N2398), .B(N2357), .CI(N2359));
ADDFX1 inst_cellmath__43_0_I1102 (.CO(N2405), .S(N2404), .A(N2361), .B(N2400), .CI(N2402));
ADDFX1 inst_cellmath__43_0_I1103 (.CO(N2407), .S(N2406), .A(N661), .B(N1740), .CI(N718));
ADDFX1 inst_cellmath__43_0_I1104 (.CO(N2409), .S(N2408), .A(N775), .B(N604), .CI(N832));
ADDFX1 inst_cellmath__43_0_I1105 (.CO(N2411), .S(N2410), .A(N946), .B(N889), .CI(N1003));
ADDFX1 inst_cellmath__43_0_I1106 (.CO(N2413), .S(N2412), .A(N1117), .B(N1060), .CI(N1174));
ADDFX1 inst_cellmath__43_0_I1107 (.CO(N2415), .S(N2414), .A(N1288), .B(N1231), .CI(N1345));
ADDFX1 inst_cellmath__43_0_I1108 (.CO(N2417), .S(N2416), .A(N1459), .B(N1402), .CI(N1516));
ADDFX1 inst_cellmath__43_0_I1109 (.CO(N2419), .S(N2418), .A(N1630), .B(N1573), .CI(N1687));
ADDFX1 inst_cellmath__43_0_I1110 (.CO(N2421), .S(N2420), .A(N2367), .B(N2365), .CI(N2369));
ADDFX1 inst_cellmath__43_0_I1111 (.CO(N2423), .S(N2422), .A(N2373), .B(N2371), .CI(N2375));
ADDFX1 inst_cellmath__43_0_I1112 (.CO(N2425), .S(N2424), .A(N2406), .B(N2377), .CI(N2408));
ADDFX1 inst_cellmath__43_0_I1113 (.CO(N2427), .S(N2426), .A(N2412), .B(N2410), .CI(N2414));
ADDFX1 inst_cellmath__43_0_I1114 (.CO(N2429), .S(N2428), .A(N2418), .B(N2416), .CI(N2379));
ADDFX1 inst_cellmath__43_0_I1115 (.CO(N2431), .S(N2430), .A(N2383), .B(N2381), .CI(N2385));
ADDFX1 inst_cellmath__43_0_I1116 (.CO(N2433), .S(N2432), .A(N2420), .B(N2387), .CI(N2422));
ADDFX1 inst_cellmath__43_0_I1117 (.CO(N2435), .S(N2434), .A(N2424), .B(N2389), .CI(N2426));
ADDFX1 inst_cellmath__43_0_I1118 (.CO(N2437), .S(N2436), .A(N2391), .B(N2428), .CI(N2393));
ADDFX1 inst_cellmath__43_0_I1119 (.CO(N2439), .S(N2438), .A(N2432), .B(N2430), .CI(N2395));
ADDFX1 inst_cellmath__43_0_I1120 (.CO(N2441), .S(N2440), .A(N2434), .B(N2397), .CI(N2436));
ADDFX1 inst_cellmath__43_0_I1121 (.CO(N2443), .S(N2442), .A(N2438), .B(N2399), .CI(N2401));
ADDFX1 inst_cellmath__43_0_I1122 (.CO(N2445), .S(N2444), .A(N2403), .B(N2440), .CI(N2442));
ADDFX1 inst_cellmath__43_0_I1123 (.CO(N2447), .S(N2446), .A(N720), .B(N1742), .CI(N777));
ADDFX1 inst_cellmath__43_0_I1124 (.CO(N2449), .S(N2448), .A(N834), .B(N663), .CI(N891));
ADDFX1 inst_cellmath__43_0_I1125 (.CO(N2451), .S(N2450), .A(N1005), .B(N948), .CI(N1062));
ADDFX1 inst_cellmath__43_0_I1126 (.CO(N2453), .S(N2452), .A(N1176), .B(N1119), .CI(N1233));
ADDFX1 inst_cellmath__43_0_I1127 (.CO(N2455), .S(N2454), .A(N1347), .B(N1290), .CI(N1404));
ADDFX1 inst_cellmath__43_0_I1128 (.CO(N2457), .S(N2456), .A(N1518), .B(N1461), .CI(N1575));
ADDFX1 inst_cellmath__43_0_I1129 (.CO(N2459), .S(N2458), .A(N1689), .B(N1632), .CI(N2407));
ADDFX1 inst_cellmath__43_0_I1130 (.CO(N2461), .S(N2460), .A(N2411), .B(N2409), .CI(N2413));
ADDFX1 inst_cellmath__43_0_I1131 (.CO(N2463), .S(N2462), .A(N2417), .B(N2415), .CI(N2419));
ADDFX1 inst_cellmath__43_0_I1132 (.CO(N2465), .S(N2464), .A(N2448), .B(N2446), .CI(N2450));
ADDFX1 inst_cellmath__43_0_I1133 (.CO(N2467), .S(N2466), .A(N2454), .B(N2452), .CI(N2456));
ADDFX1 inst_cellmath__43_0_I1134 (.CO(N2469), .S(N2468), .A(N2423), .B(N2421), .CI(N2458));
ADDFX1 inst_cellmath__43_0_I1135 (.CO(N2471), .S(N2470), .A(N2460), .B(N2425), .CI(N2462));
ADDFX1 inst_cellmath__43_0_I1136 (.CO(N2473), .S(N2472), .A(N2429), .B(N2427), .CI(N2464));
ADDFX1 inst_cellmath__43_0_I1137 (.CO(N2475), .S(N2474), .A(N2431), .B(N2466), .CI(N2433));
ADDFX1 inst_cellmath__43_0_I1138 (.CO(N2477), .S(N2476), .A(N2470), .B(N2468), .CI(N2435));
ADDFX1 inst_cellmath__43_0_I1139 (.CO(N2479), .S(N2478), .A(N2472), .B(N2437), .CI(N2474));
ADDFX1 inst_cellmath__43_0_I1140 (.CO(N2481), .S(N2480), .A(N2476), .B(N2439), .CI(N2441));
ADDFX1 inst_cellmath__43_0_I1141 (.CO(N2483), .S(N2482), .A(N2443), .B(N2478), .CI(N2480));
ADDFX1 inst_cellmath__43_0_I1142 (.CO(N2485), .S(N2484), .A(N779), .B(N1744), .CI(N836));
ADDFX1 inst_cellmath__43_0_I1143 (.CO(N2487), .S(N2486), .A(N893), .B(N722), .CI(N950));
ADDFX1 inst_cellmath__43_0_I1144 (.CO(N2489), .S(N2488), .A(N1064), .B(N1007), .CI(N1121));
ADDFX1 inst_cellmath__43_0_I1145 (.CO(N2491), .S(N2490), .A(N1235), .B(N1178), .CI(N1292));
ADDFX1 inst_cellmath__43_0_I1146 (.CO(N2493), .S(N2492), .A(N1406), .B(N1349), .CI(N1463));
ADDFX1 inst_cellmath__43_0_I1147 (.CO(N2495), .S(N2494), .A(N1577), .B(N1520), .CI(N1634));
ADDFX1 inst_cellmath__43_0_I1148 (.CO(N2497), .S(N2496), .A(N2447), .B(N1691), .CI(N2449));
ADDFX1 inst_cellmath__43_0_I1149 (.CO(N2499), .S(N2498), .A(N2453), .B(N2451), .CI(N2455));
ADDFX1 inst_cellmath__43_0_I1150 (.CO(N2501), .S(N2500), .A(N2484), .B(N2457), .CI(N2486));
ADDFX1 inst_cellmath__43_0_I1151 (.CO(N2503), .S(N2502), .A(N2490), .B(N2488), .CI(N2492));
ADDFX1 inst_cellmath__43_0_I1152 (.CO(N2505), .S(N2504), .A(N2459), .B(N2494), .CI(N2461));
ADDFX1 inst_cellmath__43_0_I1153 (.CO(N2507), .S(N2506), .A(N2465), .B(N2463), .CI(N2496));
ADDFX1 inst_cellmath__43_0_I1154 (.CO(N2509), .S(N2508), .A(N2498), .B(N2467), .CI(N2500));
ADDFX1 inst_cellmath__43_0_I1155 (.CO(N2511), .S(N2510), .A(N2469), .B(N2502), .CI(N2504));
ADDFX1 inst_cellmath__43_0_I1156 (.CO(N2513), .S(N2512), .A(N2473), .B(N2471), .CI(N2506));
ADDFX1 inst_cellmath__43_0_I1157 (.CO(N2515), .S(N2514), .A(N2508), .B(N2475), .CI(N2510));
ADDFX1 inst_cellmath__43_0_I1158 (.CO(N2517), .S(N2516), .A(N2512), .B(N2477), .CI(N2479));
ADDFX1 inst_cellmath__43_0_I1159 (.CO(N2519), .S(N2518), .A(N2481), .B(N2514), .CI(N2516));
ADDFX1 inst_cellmath__43_0_I1160 (.CO(N2521), .S(N2520), .A(N838), .B(N1746), .CI(N895));
ADDFX1 inst_cellmath__43_0_I1161 (.CO(N2523), .S(N2522), .A(N952), .B(N781), .CI(N1009));
ADDFX1 inst_cellmath__43_0_I1162 (.CO(N2525), .S(N2524), .A(N1123), .B(N1066), .CI(N1180));
ADDFX1 inst_cellmath__43_0_I1163 (.CO(N2527), .S(N2526), .A(N1294), .B(N1237), .CI(N1351));
ADDFX1 inst_cellmath__43_0_I1164 (.CO(N2529), .S(N2528), .A(N1465), .B(N1408), .CI(N1522));
ADDFX1 inst_cellmath__43_0_I1165 (.CO(N2531), .S(N2530), .A(N1636), .B(N1579), .CI(N1693));
ADDFX1 inst_cellmath__43_0_I1166 (.CO(N2533), .S(N2532), .A(N2487), .B(N2485), .CI(N2489));
ADDFX1 inst_cellmath__43_0_I1167 (.CO(N2535), .S(N2534), .A(N2493), .B(N2491), .CI(N2495));
ADDFX1 inst_cellmath__43_0_I1168 (.CO(N2537), .S(N2536), .A(N2522), .B(N2520), .CI(N2524));
ADDFX1 inst_cellmath__43_0_I1169 (.CO(N2539), .S(N2538), .A(N2528), .B(N2526), .CI(N2530));
ADDFX1 inst_cellmath__43_0_I1170 (.CO(N2541), .S(N2540), .A(N2499), .B(N2497), .CI(N2501));
ADDFX1 inst_cellmath__43_0_I1171 (.CO(N2543), .S(N2542), .A(N2532), .B(N2503), .CI(N2534));
ADDFX1 inst_cellmath__43_0_I1172 (.CO(N2545), .S(N2544), .A(N2536), .B(N2505), .CI(N2538));
ADDFX1 inst_cellmath__43_0_I1173 (.CO(N2547), .S(N2546), .A(N2509), .B(N2507), .CI(N2542));
ADDFX1 inst_cellmath__43_0_I1174 (.CO(N2549), .S(N2548), .A(N2511), .B(N2540), .CI(N2544));
ADDFX1 inst_cellmath__43_0_I1175 (.CO(N2551), .S(N2550), .A(N2546), .B(N2513), .CI(N2515));
ADDFX1 inst_cellmath__43_0_I1176 (.CO(N2553), .S(N2552), .A(N2517), .B(N2548), .CI(N2550));
ADDFX1 inst_cellmath__43_0_I1177 (.CO(N2555), .S(N2554), .A(N897), .B(N1748), .CI(N954));
ADDFX1 inst_cellmath__43_0_I1178 (.CO(N2557), .S(N2556), .A(N1011), .B(N840), .CI(N1068));
ADDFX1 inst_cellmath__43_0_I1179 (.CO(N2559), .S(N2558), .A(N1182), .B(N1125), .CI(N1239));
ADDFX1 inst_cellmath__43_0_I1180 (.CO(N2561), .S(N2560), .A(N1353), .B(N1296), .CI(N1410));
ADDFX1 inst_cellmath__43_0_I1181 (.CO(N2563), .S(N2562), .A(N1524), .B(N1467), .CI(N1581));
ADDFX1 inst_cellmath__43_0_I1182 (.CO(N2565), .S(N2564), .A(N1695), .B(N1638), .CI(N2521));
ADDFX1 inst_cellmath__43_0_I1183 (.CO(N2567), .S(N2566), .A(N2525), .B(N2523), .CI(N2527));
ADDFX1 inst_cellmath__43_0_I1184 (.CO(N2569), .S(N2568), .A(N2531), .B(N2529), .CI(N2554));
ADDFX1 inst_cellmath__43_0_I1185 (.CO(N2571), .S(N2570), .A(N2558), .B(N2556), .CI(N2560));
ADDFX1 inst_cellmath__43_0_I1186 (.CO(N2573), .S(N2572), .A(N2533), .B(N2562), .CI(N2535));
ADDFX1 inst_cellmath__43_0_I1187 (.CO(N2575), .S(N2574), .A(N2537), .B(N2564), .CI(N2566));
ADDFX1 inst_cellmath__43_0_I1188 (.CO(N2577), .S(N2576), .A(N2568), .B(N2539), .CI(N2570));
ADDFX1 inst_cellmath__43_0_I1189 (.CO(N2579), .S(N2578), .A(N2543), .B(N2541), .CI(N2572));
ADDFX1 inst_cellmath__43_0_I1190 (.CO(N2581), .S(N2580), .A(N2545), .B(N2574), .CI(N2576));
ADDFX1 inst_cellmath__43_0_I1191 (.CO(N2583), .S(N2582), .A(N2578), .B(N2547), .CI(N2549));
ADDFX1 inst_cellmath__43_0_I1192 (.CO(N2585), .S(N2584), .A(N2551), .B(N2580), .CI(N2582));
ADDFX1 inst_cellmath__43_0_I1193 (.CO(N2587), .S(N2586), .A(N956), .B(N1750), .CI(N1013));
ADDFX1 inst_cellmath__43_0_I1194 (.CO(N2589), .S(N2588), .A(N1070), .B(N899), .CI(N1127));
ADDFX1 inst_cellmath__43_0_I1195 (.CO(N2591), .S(N2590), .A(N1241), .B(N1184), .CI(N1298));
ADDFX1 inst_cellmath__43_0_I1196 (.CO(N2593), .S(N2592), .A(N1412), .B(N1355), .CI(N1469));
ADDFX1 inst_cellmath__43_0_I1197 (.CO(N2595), .S(N2594), .A(N1583), .B(N1526), .CI(N1640));
ADDFX1 inst_cellmath__43_0_I1198 (.CO(N2597), .S(N2596), .A(N2555), .B(N1697), .CI(N2557));
ADDFX1 inst_cellmath__43_0_I1199 (.CO(N2599), .S(N2598), .A(N2561), .B(N2559), .CI(N2563));
ADDFX1 inst_cellmath__43_0_I1200 (.CO(N2601), .S(N2600), .A(N2588), .B(N2586), .CI(N2590));
ADDFX1 inst_cellmath__43_0_I1201 (.CO(N2603), .S(N2602), .A(N2594), .B(N2592), .CI(N2565));
ADDFX1 inst_cellmath__43_0_I1202 (.CO(N2605), .S(N2604), .A(N2569), .B(N2567), .CI(N2571));
ADDFX1 inst_cellmath__43_0_I1203 (.CO(N2607), .S(N2606), .A(N2598), .B(N2596), .CI(N2573));
ADDFX1 inst_cellmath__43_0_I1204 (.CO(N2609), .S(N2608), .A(N2602), .B(N2600), .CI(N2575));
ADDFX1 inst_cellmath__43_0_I1205 (.CO(N2611), .S(N2610), .A(N2577), .B(N2604), .CI(N2606));
ADDFX1 inst_cellmath__43_0_I1206 (.CO(N2613), .S(N2612), .A(N2608), .B(N2579), .CI(N2581));
ADDFX1 inst_cellmath__43_0_I1207 (.CO(N2615), .S(N2614), .A(N2583), .B(N2610), .CI(N2612));
ADDFX1 inst_cellmath__43_0_I1208 (.CO(N2617), .S(N2616), .A(N1015), .B(N1752), .CI(N1072));
ADDFX1 inst_cellmath__43_0_I1209 (.CO(N2619), .S(N2618), .A(N1129), .B(N958), .CI(N1186));
ADDFX1 inst_cellmath__43_0_I1210 (.CO(N2621), .S(N2620), .A(N1300), .B(N1243), .CI(N1357));
ADDFX1 inst_cellmath__43_0_I1211 (.CO(N2623), .S(N2622), .A(N1471), .B(N1414), .CI(N1528));
ADDFX1 inst_cellmath__43_0_I1212 (.CO(N2625), .S(N2624), .A(N1642), .B(N1585), .CI(N1699));
ADDFX1 inst_cellmath__43_0_I1213 (.CO(N2627), .S(N2626), .A(N2589), .B(N2587), .CI(N2591));
ADDFX1 inst_cellmath__43_0_I1214 (.CO(N2629), .S(N2628), .A(N2595), .B(N2593), .CI(N2616));
ADDFX1 inst_cellmath__43_0_I1215 (.CO(N2631), .S(N2630), .A(N2620), .B(N2618), .CI(N2622));
ADDFX1 inst_cellmath__43_0_I1216 (.CO(N2633), .S(N2632), .A(N2597), .B(N2624), .CI(N2599));
ADDFX1 inst_cellmath__43_0_I1217 (.CO(N2635), .S(N2634), .A(N2626), .B(N2601), .CI(N2603));
ADDFX1 inst_cellmath__43_0_I1218 (.CO(N2637), .S(N2636), .A(N2630), .B(N2628), .CI(N2605));
ADDFX1 inst_cellmath__43_0_I1219 (.CO(N2639), .S(N2638), .A(N2607), .B(N2632), .CI(N2634));
ADDFX1 inst_cellmath__43_0_I1220 (.CO(N2641), .S(N2640), .A(N2636), .B(N2609), .CI(N2611));
ADDFX1 inst_cellmath__43_0_I1221 (.CO(N2643), .S(N2642), .A(N2613), .B(N2638), .CI(N2640));
ADDFX1 inst_cellmath__43_0_I1222 (.CO(N2645), .S(N2644), .A(N1074), .B(N1754), .CI(N1131));
ADDFX1 inst_cellmath__43_0_I1223 (.CO(N2647), .S(N2646), .A(N1188), .B(N1017), .CI(N1245));
ADDFX1 inst_cellmath__43_0_I1224 (.CO(N2649), .S(N2648), .A(N1359), .B(N1302), .CI(N1416));
ADDFX1 inst_cellmath__43_0_I1225 (.CO(N2651), .S(N2650), .A(N1530), .B(N1473), .CI(N1587));
ADDFX1 inst_cellmath__43_0_I1226 (.CO(N2653), .S(N2652), .A(N1701), .B(N1644), .CI(N2617));
ADDFX1 inst_cellmath__43_0_I1227 (.CO(N2655), .S(N2654), .A(N2621), .B(N2619), .CI(N2623));
ADDFX1 inst_cellmath__43_0_I1228 (.CO(N2657), .S(N2656), .A(N2644), .B(N2625), .CI(N2646));
ADDFX1 inst_cellmath__43_0_I1229 (.CO(N2659), .S(N2658), .A(N2650), .B(N2648), .CI(N2627));
ADDFX1 inst_cellmath__43_0_I1230 (.CO(N2661), .S(N2660), .A(N2629), .B(N2652), .CI(N2631));
ADDFX1 inst_cellmath__43_0_I1231 (.CO(N2663), .S(N2662), .A(N2656), .B(N2654), .CI(N2633));
ADDFX1 inst_cellmath__43_0_I1232 (.CO(N2665), .S(N2664), .A(N2635), .B(N2658), .CI(N2660));
ADDFX1 inst_cellmath__43_0_I1233 (.CO(N2667), .S(N2666), .A(N2662), .B(N2637), .CI(N2639));
ADDFX1 inst_cellmath__43_0_I1234 (.CO(N2669), .S(N2668), .A(N2641), .B(N2664), .CI(N2666));
ADDFX1 inst_cellmath__43_0_I1235 (.CO(N2671), .S(N2670), .A(N1133), .B(N1756), .CI(N1190));
ADDFX1 inst_cellmath__43_0_I1236 (.CO(N2673), .S(N2672), .A(N1247), .B(N1076), .CI(N1304));
ADDFX1 inst_cellmath__43_0_I1237 (.CO(N2675), .S(N2674), .A(N1418), .B(N1361), .CI(N1475));
ADDFX1 inst_cellmath__43_0_I1238 (.CO(N2677), .S(N2676), .A(N1589), .B(N1532), .CI(N1646));
ADDFX1 inst_cellmath__43_0_I1239 (.CO(N2679), .S(N2678), .A(N2645), .B(N1703), .CI(N2647));
ADDFX1 inst_cellmath__43_0_I1240 (.CO(N2681), .S(N2680), .A(N2651), .B(N2649), .CI(N2670));
ADDFX1 inst_cellmath__43_0_I1241 (.CO(N2683), .S(N2682), .A(N2674), .B(N2672), .CI(N2676));
ADDFX1 inst_cellmath__43_0_I1242 (.CO(N2685), .S(N2684), .A(N2655), .B(N2653), .CI(N2657));
ADDFX1 inst_cellmath__43_0_I1243 (.CO(N2687), .S(N2686), .A(N2659), .B(N2678), .CI(N2680));
ADDFX1 inst_cellmath__43_0_I1244 (.CO(N2689), .S(N2688), .A(N2661), .B(N2682), .CI(N2684));
ADDFX1 inst_cellmath__43_0_I1245 (.CO(N2691), .S(N2690), .A(N2686), .B(N2663), .CI(N2665));
ADDFX1 inst_cellmath__43_0_I1246 (.CO(N2693), .S(N2692), .A(N2667), .B(N2688), .CI(N2690));
ADDFX1 inst_cellmath__43_0_I1247 (.CO(N2695), .S(N2694), .A(N1192), .B(N1758), .CI(N1249));
ADDFX1 inst_cellmath__43_0_I1248 (.CO(N2697), .S(N2696), .A(N1306), .B(N1135), .CI(N1363));
ADDFX1 inst_cellmath__43_0_I1249 (.CO(N2699), .S(N2698), .A(N1477), .B(N1420), .CI(N1534));
ADDFX1 inst_cellmath__43_0_I1250 (.CO(N2701), .S(N2700), .A(N1648), .B(N1591), .CI(N1705));
ADDFX1 inst_cellmath__43_0_I1251 (.CO(N2703), .S(N2702), .A(N2673), .B(N2671), .CI(N2675));
ADDFX1 inst_cellmath__43_0_I1252 (.CO(N2705), .S(N2704), .A(N2694), .B(N2677), .CI(N2696));
ADDFX1 inst_cellmath__43_0_I1253 (.CO(N2707), .S(N2706), .A(N2700), .B(N2698), .CI(N2679));
ADDFX1 inst_cellmath__43_0_I1254 (.CO(N2709), .S(N2708), .A(N2683), .B(N2681), .CI(N2702));
ADDFX1 inst_cellmath__43_0_I1255 (.CO(N2711), .S(N2710), .A(N2685), .B(N2704), .CI(N2706));
ADDFX1 inst_cellmath__43_0_I1256 (.CO(N2713), .S(N2712), .A(N2708), .B(N2687), .CI(N2689));
ADDFX1 inst_cellmath__43_0_I1257 (.CO(N2715), .S(N2714), .A(N2691), .B(N2710), .CI(N2712));
ADDFX1 inst_cellmath__43_0_I1258 (.CO(N2717), .S(N2716), .A(N1251), .B(N1760), .CI(N1308));
ADDFX1 inst_cellmath__43_0_I1259 (.CO(N2719), .S(N2718), .A(N1365), .B(N1194), .CI(N1422));
ADDFX1 inst_cellmath__43_0_I1260 (.CO(N2721), .S(N2720), .A(N1536), .B(N1479), .CI(N1593));
ADDFX1 inst_cellmath__43_0_I1261 (.CO(N2723), .S(N2722), .A(N1707), .B(N1650), .CI(N2695));
ADDFX1 inst_cellmath__43_0_I1262 (.CO(N2725), .S(N2724), .A(N2699), .B(N2697), .CI(N2701));
ADDFX1 inst_cellmath__43_0_I1263 (.CO(N2727), .S(N2726), .A(N2718), .B(N2716), .CI(N2720));
ADDFX1 inst_cellmath__43_0_I1264 (.CO(N2729), .S(N2728), .A(N2722), .B(N2703), .CI(N2705));
ADDFX1 inst_cellmath__43_0_I1265 (.CO(N2731), .S(N2730), .A(N2707), .B(N2724), .CI(N2726));
ADDFX1 inst_cellmath__43_0_I1266 (.CO(N2733), .S(N2732), .A(N2728), .B(N2709), .CI(N2711));
ADDFX1 inst_cellmath__43_0_I1267 (.CO(N2735), .S(N2734), .A(N2713), .B(N2730), .CI(N2732));
ADDFX1 inst_cellmath__43_0_I1268 (.CO(N2737), .S(N2736), .A(N1310), .B(N1762), .CI(N1367));
ADDFX1 inst_cellmath__43_0_I1269 (.CO(N2739), .S(N2738), .A(N1424), .B(N1253), .CI(N1481));
ADDFX1 inst_cellmath__43_0_I1270 (.CO(N2741), .S(N2740), .A(N1595), .B(N1538), .CI(N1652));
ADDFX1 inst_cellmath__43_0_I1271 (.CO(N2743), .S(N2742), .A(N2717), .B(N1709), .CI(N2719));
ADDFX1 inst_cellmath__43_0_I1272 (.CO(N2745), .S(N2744), .A(N2736), .B(N2721), .CI(N2738));
ADDFX1 inst_cellmath__43_0_I1273 (.CO(N2747), .S(N2746), .A(N2723), .B(N2740), .CI(N2725));
ADDFX1 inst_cellmath__43_0_I1274 (.CO(N2749), .S(N2748), .A(N2742), .B(N2727), .CI(N2744));
ADDFX1 inst_cellmath__43_0_I1275 (.CO(N2751), .S(N2750), .A(N2746), .B(N2729), .CI(N2731));
ADDFX1 inst_cellmath__43_0_I1276 (.CO(N2753), .S(N2752), .A(N2733), .B(N2748), .CI(N2750));
ADDFX1 inst_cellmath__43_0_I1277 (.CO(N2755), .S(N2754), .A(N1369), .B(N1764), .CI(N1426));
ADDFX1 inst_cellmath__43_0_I1278 (.CO(N2757), .S(N2756), .A(N1483), .B(N1312), .CI(N1540));
ADDFX1 inst_cellmath__43_0_I1279 (.CO(N2759), .S(N2758), .A(N1654), .B(N1597), .CI(N1711));
ADDFX1 inst_cellmath__43_0_I1280 (.CO(N2761), .S(N2760), .A(N2739), .B(N2737), .CI(N2741));
ADDFX1 inst_cellmath__43_0_I1281 (.CO(N2763), .S(N2762), .A(N2756), .B(N2754), .CI(N2758));
ADDFX1 inst_cellmath__43_0_I1282 (.CO(N2765), .S(N2764), .A(N2745), .B(N2743), .CI(N2760));
ADDFX1 inst_cellmath__43_0_I1283 (.CO(N2767), .S(N2766), .A(N2762), .B(N2747), .CI(N2749));
ADDFX1 inst_cellmath__43_0_I1284 (.CO(N2769), .S(N2768), .A(N2751), .B(N2764), .CI(N2766));
ADDFX1 inst_cellmath__43_0_I1285 (.CO(N2771), .S(N2770), .A(N1428), .B(N1766), .CI(N1485));
ADDFX1 inst_cellmath__43_0_I1286 (.CO(N2773), .S(N2772), .A(N1542), .B(N1371), .CI(N1599));
ADDFX1 inst_cellmath__43_0_I1287 (.CO(N2775), .S(N2774), .A(N1713), .B(N1656), .CI(N2755));
ADDFX1 inst_cellmath__43_0_I1288 (.CO(N2777), .S(N2776), .A(N2759), .B(N2757), .CI(N2770));
ADDFX1 inst_cellmath__43_0_I1289 (.CO(N2779), .S(N2778), .A(N2761), .B(N2772), .CI(N2774));
ADDFX1 inst_cellmath__43_0_I1290 (.CO(N2781), .S(N2780), .A(N2776), .B(N2763), .CI(N2765));
ADDFX1 inst_cellmath__43_0_I1291 (.CO(N2783), .S(N2782), .A(N2767), .B(N2778), .CI(N2780));
ADDFX1 inst_cellmath__43_0_I1292 (.CO(N2785), .S(N2784), .A(N1487), .B(N1768), .CI(N1544));
ADDFX1 inst_cellmath__43_0_I1293 (.CO(N2787), .S(N2786), .A(N1601), .B(N1430), .CI(N1658));
ADDFX1 inst_cellmath__43_0_I1294 (.CO(N2789), .S(N2788), .A(N2771), .B(N1715), .CI(N2773));
ADDFX1 inst_cellmath__43_0_I1295 (.CO(N2791), .S(N2790), .A(N2786), .B(N2784), .CI(N2775));
ADDFX1 inst_cellmath__43_0_I1296 (.CO(N2793), .S(N2792), .A(N2788), .B(N2777), .CI(N2779));
ADDFX1 inst_cellmath__43_0_I1297 (.CO(N2795), .S(N2794), .A(N2781), .B(N2790), .CI(N2792));
ADDFX1 inst_cellmath__43_0_I1298 (.CO(N2797), .S(N2796), .A(N1546), .B(N1770), .CI(N1603));
ADDFX1 inst_cellmath__43_0_I1299 (.CO(N2799), .S(N2798), .A(N1660), .B(N1489), .CI(N1717));
ADDFX1 inst_cellmath__43_0_I1300 (.CO(N2801), .S(N2800), .A(N2787), .B(N2785), .CI(N2796));
ADDFX1 inst_cellmath__43_0_I1301 (.CO(N2803), .S(N2802), .A(N2789), .B(N2798), .CI(N2791));
ADDFX1 inst_cellmath__43_0_I1302 (.CO(N2805), .S(N2804), .A(N2793), .B(N2800), .CI(N2802));
ADDFX1 inst_cellmath__43_0_I1303 (.CO(N2807), .S(N2806), .A(N1605), .B(N1772), .CI(N1662));
ADDFX1 inst_cellmath__43_0_I1304 (.CO(N2809), .S(N2808), .A(N1719), .B(N1548), .CI(N2797));
ADDFX1 inst_cellmath__43_0_I1305 (.CO(N2811), .S(N2810), .A(N2806), .B(N2799), .CI(N2808));
ADDFX1 inst_cellmath__43_0_I1306 (.CO(N2813), .S(N2812), .A(N2803), .B(N2801), .CI(N2810));
ADDFX1 inst_cellmath__43_0_I1307 (.CO(N2815), .S(N2814), .A(N1664), .B(N1774), .CI(N1721));
ADDFX1 inst_cellmath__43_0_I1308 (.CO(N2817), .S(N2816), .A(N2807), .B(N1607), .CI(N2814));
ADDFX1 inst_cellmath__43_0_I1309 (.CO(N2819), .S(N2818), .A(N2816), .B(N2809), .CI(N2811));
ADDFX1 inst_cellmath__43_0_I1310 (.CO(N2821), .S(N2820), .A(N1723), .B(N1776), .CI(N1666));
ADDFX1 inst_cellmath__43_0_I1311 (.CO(N2823), .S(N2822), .A(N2820), .B(N2815), .CI(N2817));
ADDFX1 inst_cellmath__43_0_I1312 (.CO(N3376), .S(N2824), .A(N1725), .B(N1778), .CI(N2821));
NAND2XL inst_cellmath__43_0_I1313 (.Y(N2826), .A(N383), .B(N440));
NOR2XL inst_cellmath__43_0_I1314 (.Y(N2827), .A(N499), .B(N1812));
NAND2XL inst_cellmath__43_0_I1315 (.Y(N2828), .A(N499), .B(N1812));
NOR2XL inst_cellmath__43_0_I1316 (.Y(N2829), .A(N1814), .B(N1816));
NAND2XL inst_cellmath__43_0_I1317 (.Y(N2830), .A(N1814), .B(N1816));
NOR2XL inst_cellmath__43_0_I1318 (.Y(N2831), .A(N1820), .B(N1822));
NAND2XL inst_cellmath__43_0_I1319 (.Y(N2832), .A(N1820), .B(N1822));
NOR2XL inst_cellmath__43_0_I1320 (.Y(N2833), .A(N1823), .B(N1830));
AND2XL inst_cellmath__43_0_I2164 (.Y(N3636), .A(N1823), .B(N1830));
NOR2XL inst_cellmath__43_0_I1322 (.Y(N2835), .A(N1831), .B(N1840));
NAND2XL inst_cellmath__43_0_I1323 (.Y(N2836), .A(N1831), .B(N1840));
NOR2XL inst_cellmath__43_0_I1324 (.Y(N2837), .A(N1841), .B(N1852));
NAND2XL inst_cellmath__43_0_I1325 (.Y(N2838), .A(N1841), .B(N1852));
NOR2XL inst_cellmath__43_0_I1326 (.Y(N2839), .A(N1853), .B(N1866));
NAND2XL inst_cellmath__43_0_I1327 (.Y(N2840), .A(N1853), .B(N1866));
NOR2XL inst_cellmath__43_0_I1328 (.Y(N2841), .A(N1867), .B(N1882));
NAND2XL inst_cellmath__43_0_I1329 (.Y(N2842), .A(N1867), .B(N1882));
NOR2XL inst_cellmath__43_0_I1330 (.Y(N2843), .A(N1883), .B(N1900));
NAND2XL inst_cellmath__43_0_I1331 (.Y(N2844), .A(N1883), .B(N1900));
NOR2XL inst_cellmath__43_0_I1332 (.Y(N2845), .A(N1901), .B(N1920));
NAND2XL inst_cellmath__43_0_I1333 (.Y(N2846), .A(N1901), .B(N1920));
NOR2XL inst_cellmath__43_0_I1334 (.Y(N2847), .A(N1921), .B(N1942));
NAND2XL inst_cellmath__43_0_I1335 (.Y(N2848), .A(N1921), .B(N1942));
NOR2XL inst_cellmath__43_0_I1336 (.Y(N2849), .A(N1943), .B(N1966));
NAND2XL inst_cellmath__43_0_I1337 (.Y(N2850), .A(N1943), .B(N1966));
NOR2XL inst_cellmath__43_0_I1338 (.Y(N2851), .A(N1967), .B(N1992));
NAND2XL inst_cellmath__43_0_I1339 (.Y(N2852), .A(N1967), .B(N1992));
NOR2XL inst_cellmath__43_0_I1340 (.Y(N2853), .A(N1993), .B(N2020));
NAND2XL inst_cellmath__43_0_I1341 (.Y(N2854), .A(N1993), .B(N2020));
NOR2XL inst_cellmath__43_0_I1342 (.Y(N2855), .A(N2021), .B(N2050));
NAND2XL inst_cellmath__43_0_I1343 (.Y(N2856), .A(N2021), .B(N2050));
AOI21XL inst_cellmath__43_0_I1346 (.Y(N2859), .A0(N2828), .A1(N2826), .B0(N2827));
INVXL inst_cellmath__43_0_I2045 (.Y(N3639), .A(N2829));
INVXL inst_cellmath__43_0_I2046 (.Y(N3640), .A(N2830));
OAI21XL inst_cellmath__43_0_I1354 (.Y(N2867), .A0(N3640), .A1(N2859), .B0(N3639));
AOI21XL inst_cellmath__43_0_I1362 (.Y(N2875), .A0(N2832), .A1(N2867), .B0(N2831));
INVXL inst_cellmath__43_0_I2052 (.Y(N3646), .A(N2833));
OAI21XL inst_cellmath__43_0_I1374 (.Y(N2887), .A0(N3636), .A1(N2875), .B0(N3646));
AOI21XL inst_cellmath__43_0_I1386 (.Y(N2899), .A0(N2836), .A1(N2887), .B0(N2835));
INVXL inst_cellmath__43_0_I2063 (.Y(N3657), .A(N2837));
INVXL inst_cellmath__43_0_I2064 (.Y(N3658), .A(N2838));
OAI21XL inst_cellmath__43_0_I1402 (.Y(N2915), .A0(N3658), .A1(N2899), .B0(N3657));
AOI21XL inst_cellmath__43_0_I1418 (.Y(N2931), .A0(N2840), .A1(N2915), .B0(N2839));
AOI21XL inst_cellmath__43_0_I1422 (.Y(N2935), .A0(N2844), .A1(N2841), .B0(N2843));
NAND2XL inst_cellmath__43_0_I1423 (.Y(N2936), .A(N2844), .B(N2842));
OAI21XL inst_cellmath__43_0_I1442 (.Y(N2955), .A0(N2936), .A1(N2931), .B0(N2935));
AOI21XL inst_cellmath__43_0_I1446 (.Y(N2959), .A0(N2848), .A1(N2845), .B0(N2847));
INVXL inst_cellmath__43_0_I2096 (.Y(N3690), .A(N2959));
AOI21XL inst_cellmath__43_0_I1472 (.Y(N2985), .A0(N2846), .A1(N2955), .B0(N2845));
AOI31X1 inst_cellmath__43_0_I5053 (.Y(N2987), .A0(N2848), .A1(N2846), .A2(N2955), .B0(N3690));
AOI21XL inst_cellmath__43_0_I1478 (.Y(N2991), .A0(N2852), .A1(N2849), .B0(N2851));
NAND2XL inst_cellmath__43_0_I1479 (.Y(N2992), .A(N2852), .B(N2850));
OAI21XL inst_cellmath__43_0_I1506 (.Y(N3019), .A0(N2992), .A1(N2987), .B0(N2991));
AO21XL inst_cellmath__43_0_I2200 (.Y(N3724), .A0(N2856), .A1(N2853), .B0(N2855));
NOR2BX1 andori2bb1_A_I5054 (.Y(N3757), .AN(N2842), .B(N2931));
NOR2XL andori2bb1_A_I2222 (.Y(N3734), .A(N3757), .B(N2841));
NOR2BX1 andori2bb1_A_I5055 (.Y(N3764), .AN(N2850), .B(N2987));
NOR2XL andori2bb1_A_I2224 (.Y(N3738), .A(N3764), .B(N2849));
AOI21XL inst_cellmath__43_0_I1544 (.Y(N3057), .A0(N2854), .A1(N3019), .B0(N2853));
AOI31X1 inst_cellmath__43_0_I2173 (.Y(N3059), .A0(N2856), .A1(N2854), .A2(N3019), .B0(N3724));
NAND2BXL inst_cellmath__43_0_I1569 (.Y(N3082), .AN(N2827), .B(N2828));
NAND2BXL inst_cellmath__43_0_I1572 (.Y(N3085), .AN(N2829), .B(N2830));
NAND2BXL inst_cellmath__43_0_I1575 (.Y(N3088), .AN(N2831), .B(N2832));
OR2XL inst_cellmath__43_0_I2174 (.Y(N3091), .A(N3636), .B(N2833));
NAND2BXL inst_cellmath__43_0_I1581 (.Y(N3094), .AN(N2835), .B(N2836));
NAND2BXL inst_cellmath__43_0_I1584 (.Y(N3097), .AN(N2837), .B(N2838));
NAND2BXL inst_cellmath__43_0_I1587 (.Y(N3100), .AN(N2839), .B(N2840));
NAND2BXL inst_cellmath__43_0_I1590 (.Y(N3103), .AN(N2841), .B(N2842));
NAND2BXL inst_cellmath__43_0_I1593 (.Y(N3106), .AN(N2843), .B(N2844));
NAND2BXL inst_cellmath__43_0_I1596 (.Y(N3109), .AN(N2845), .B(N2846));
NAND2BXL inst_cellmath__43_0_I1599 (.Y(N3112), .AN(N2847), .B(N2848));
NAND2BXL inst_cellmath__43_0_I1602 (.Y(N3115), .AN(N2849), .B(N2850));
NAND2BXL inst_cellmath__43_0_I1605 (.Y(N3118), .AN(N2851), .B(N2852));
NAND2BXL inst_cellmath__43_0_I1608 (.Y(N3121), .AN(N2853), .B(N2854));
NAND2BXL inst_cellmath__43_0_I1611 (.Y(N3124), .AN(N2855), .B(N2856));
XOR2XL inst_cellmath__43_0_I1612 (.Y(inst_cellmath__43_0_out0[1]), .A(N383), .B(N440));
XOR2XL inst_cellmath__43_0_I2175 (.Y(inst_cellmath__43_0_out0[2]), .A(N2826), .B(N3082));
XNOR2X1 inst_cellmath__43_0_I2176 (.Y(inst_cellmath__43_0_out0[3]), .A(N2859), .B(N3085));
XOR2XL inst_cellmath__43_0_I2203 (.Y(inst_cellmath__43_0_out0[4]), .A(N2867), .B(N3088));
XNOR2X1 inst_cellmath__43_0_I2178 (.Y(inst_cellmath__43_0_out0[5]), .A(N2875), .B(N3091));
XOR2XL inst_cellmath__43_0_I2204 (.Y(inst_cellmath__43_0_out0[6]), .A(N2887), .B(N3094));
XNOR2X1 inst_cellmath__43_0_I2180 (.Y(inst_cellmath__43_0_out0[7]), .A(N2899), .B(N3097));
XOR2XL inst_cellmath__43_0_I2205 (.Y(inst_cellmath__43_0_out0[8]), .A(N2915), .B(N3100));
XNOR2X1 inst_cellmath__43_0_I2182 (.Y(inst_cellmath__43_0_out0[9]), .A(N2931), .B(N3103));
XNOR2X1 inst_cellmath__43_0_I2183 (.Y(inst_cellmath__43_0_out0[10]), .A(N3734), .B(N3106));
XOR2XL inst_cellmath__43_0_I2206 (.Y(inst_cellmath__43_0_out0[11]), .A(N2955), .B(N3109));
XNOR2X1 inst_cellmath__43_0_I2185 (.Y(inst_cellmath__43_0_out0[12]), .A(N2985), .B(N3112));
XNOR2X1 inst_cellmath__43_0_I2186 (.Y(inst_cellmath__43_0_out0[13]), .A(N2987), .B(N3115));
XNOR2X1 inst_cellmath__43_0_I1625 (.Y(inst_cellmath__43_0_out0[14]), .A(N3738), .B(N3118));
XOR2XL inst_cellmath__43_0_I2187 (.Y(inst_cellmath__43_0_out0[15]), .A(N3019), .B(N3121));
XNOR2X1 inst_cellmath__43_0_I1627 (.Y(inst_cellmath__43_0_out0[16]), .A(N3057), .B(N3124));
INVXL inst_cellmath__43_0_I1628 (.Y(N3141), .A(N3059));
NOR2XL inst_cellmath__43_0_I1629 (.Y(N3143), .A(N2051), .B(N2082));
XOR2XL inst_cellmath__43_0_I1630 (.Y(N3144), .A(N2051), .B(N2082));
NOR2XL inst_cellmath__43_0_I1631 (.Y(N3145), .A(N2083), .B(N2116));
XOR2XL inst_cellmath__43_0_I1632 (.Y(N3146), .A(N2083), .B(N2116));
NOR2XL inst_cellmath__43_0_I1633 (.Y(N3147), .A(N2117), .B(N2152));
XOR2XL inst_cellmath__43_0_I1634 (.Y(N3148), .A(N2117), .B(N2152));
NOR2XL inst_cellmath__43_0_I1635 (.Y(N3149), .A(N2153), .B(N2190));
XOR2XL inst_cellmath__43_0_I1636 (.Y(N3150), .A(N2153), .B(N2190));
NOR2XL inst_cellmath__43_0_I1637 (.Y(N3151), .A(N2191), .B(N2230));
XOR2XL inst_cellmath__43_0_I1638 (.Y(N3152), .A(N2191), .B(N2230));
NOR2XL inst_cellmath__43_0_I1639 (.Y(N3153), .A(N2231), .B(N2274));
XOR2XL inst_cellmath__43_0_I1640 (.Y(N3154), .A(N2231), .B(N2274));
NOR2XL inst_cellmath__43_0_I1641 (.Y(N3155), .A(N2275), .B(N2318));
XOR2XL inst_cellmath__43_0_I1642 (.Y(N3156), .A(N2275), .B(N2318));
NOR2XL inst_cellmath__43_0_I1643 (.Y(N3157), .A(N2319), .B(N2362));
XOR2XL inst_cellmath__43_0_I1644 (.Y(N3158), .A(N2319), .B(N2362));
NOR2XL inst_cellmath__43_0_I1645 (.Y(N3159), .A(N2363), .B(N2404));
XOR2XL inst_cellmath__43_0_I1646 (.Y(N3160), .A(N2363), .B(N2404));
NOR2XL inst_cellmath__43_0_I1647 (.Y(N3161), .A(N2405), .B(N2444));
XOR2XL inst_cellmath__43_0_I1648 (.Y(N3162), .A(N2405), .B(N2444));
NOR2XL inst_cellmath__43_0_I1649 (.Y(N3163), .A(N2445), .B(N2482));
XOR2XL inst_cellmath__43_0_I1650 (.Y(N3164), .A(N2445), .B(N2482));
NOR2XL inst_cellmath__43_0_I1651 (.Y(N3165), .A(N2483), .B(N2518));
XOR2XL inst_cellmath__43_0_I1652 (.Y(N3166), .A(N2483), .B(N2518));
NOR2XL inst_cellmath__43_0_I1653 (.Y(N3167), .A(N2519), .B(N2552));
XOR2XL inst_cellmath__43_0_I1654 (.Y(N3168), .A(N2519), .B(N2552));
NOR2XL inst_cellmath__43_0_I1655 (.Y(N3169), .A(N2553), .B(N2584));
XOR2XL inst_cellmath__43_0_I1656 (.Y(N3170), .A(N2553), .B(N2584));
NOR2XL inst_cellmath__43_0_I1657 (.Y(N3171), .A(N2585), .B(N2614));
XOR2XL inst_cellmath__43_0_I1658 (.Y(N3172), .A(N2585), .B(N2614));
NOR2XL inst_cellmath__43_0_I1659 (.Y(N3173), .A(N2615), .B(N2642));
XOR2XL inst_cellmath__43_0_I1660 (.Y(N3174), .A(N2615), .B(N2642));
NOR2XL inst_cellmath__43_0_I1661 (.Y(N3175), .A(N2643), .B(N2668));
XOR2XL inst_cellmath__43_0_I1662 (.Y(N3176), .A(N2643), .B(N2668));
NOR2XL inst_cellmath__43_0_I1663 (.Y(N3177), .A(N2669), .B(N2692));
XOR2XL inst_cellmath__43_0_I1664 (.Y(N3178), .A(N2669), .B(N2692));
NOR2XL inst_cellmath__43_0_I1665 (.Y(N3179), .A(N2693), .B(N2714));
XOR2XL inst_cellmath__43_0_I1666 (.Y(N3180), .A(N2693), .B(N2714));
NOR2XL inst_cellmath__43_0_I1667 (.Y(N3181), .A(N2715), .B(N2734));
XOR2XL inst_cellmath__43_0_I1668 (.Y(N3182), .A(N2715), .B(N2734));
NOR2XL inst_cellmath__43_0_I1669 (.Y(N3183), .A(N2735), .B(N2752));
XOR2XL inst_cellmath__43_0_I1670 (.Y(N3184), .A(N2735), .B(N2752));
NOR2XL inst_cellmath__43_0_I1671 (.Y(N3185), .A(N2753), .B(N2768));
XOR2XL inst_cellmath__43_0_I1672 (.Y(N3186), .A(N2753), .B(N2768));
NOR2XL inst_cellmath__43_0_I1673 (.Y(N3187), .A(N2769), .B(N2782));
XOR2XL inst_cellmath__43_0_I1674 (.Y(N3188), .A(N2769), .B(N2782));
NOR2XL inst_cellmath__43_0_I1675 (.Y(N3189), .A(N2783), .B(N2794));
XOR2XL inst_cellmath__43_0_I1676 (.Y(N3190), .A(N2783), .B(N2794));
NOR2XL inst_cellmath__43_0_I1677 (.Y(N3191), .A(N2795), .B(N2804));
XOR2XL inst_cellmath__43_0_I1678 (.Y(N3192), .A(N2795), .B(N2804));
NOR2XL inst_cellmath__43_0_I1679 (.Y(N3193), .A(N2805), .B(N2812));
XOR2XL inst_cellmath__43_0_I1680 (.Y(N3194), .A(N2805), .B(N2812));
NOR2XL inst_cellmath__43_0_I1681 (.Y(N3195), .A(N2818), .B(N2813));
XOR2XL inst_cellmath__43_0_I1682 (.Y(N3196), .A(N2818), .B(N2813));
NOR2XL inst_cellmath__43_0_I1683 (.Y(N3197), .A(N2822), .B(N2819));
XOR2XL inst_cellmath__43_0_I1684 (.Y(N3198), .A(N2822), .B(N2819));
NOR2XL inst_cellmath__43_0_I1685 (.Y(N3199), .A(N2824), .B(N2823));
XOR2XL inst_cellmath__43_0_I1686 (.Y(N3200), .A(N2824), .B(N2823));
AOI21XL inst_cellmath__43_0_I1688 (.Y(N3202), .A0(N3144), .A1(N3141), .B0(N3143));
AOI21XL inst_cellmath__43_0_I1690 (.Y(N3204), .A0(N3148), .A1(N3145), .B0(N3147));
NAND2XL inst_cellmath__43_0_I1691 (.Y(N3205), .A(N3148), .B(N3146));
AOI21XL inst_cellmath__43_0_I1692 (.Y(N3206), .A0(N3152), .A1(N3149), .B0(N3151));
NAND2XL inst_cellmath__43_0_I1693 (.Y(N3207), .A(N3152), .B(N3150));
AOI21XL inst_cellmath__43_0_I1694 (.Y(N3208), .A0(N3156), .A1(N3153), .B0(N3155));
NAND2XL inst_cellmath__43_0_I1695 (.Y(N3209), .A(N3156), .B(N3154));
AOI21XL inst_cellmath__43_0_I1696 (.Y(N3210), .A0(N3160), .A1(N3157), .B0(N3159));
NAND2XL inst_cellmath__43_0_I1697 (.Y(N3211), .A(N3160), .B(N3158));
AOI21XL inst_cellmath__43_0_I1698 (.Y(N3212), .A0(N3164), .A1(N3161), .B0(N3163));
NAND2XL inst_cellmath__43_0_I1699 (.Y(N3213), .A(N3164), .B(N3162));
AOI21XL inst_cellmath__43_0_I1700 (.Y(N3214), .A0(N3168), .A1(N3165), .B0(N3167));
NAND2XL inst_cellmath__43_0_I1701 (.Y(N3215), .A(N3168), .B(N3166));
AOI21XL inst_cellmath__43_0_I1702 (.Y(N3216), .A0(N3172), .A1(N3169), .B0(N3171));
NAND2XL inst_cellmath__43_0_I1703 (.Y(N3217), .A(N3172), .B(N3170));
AOI21XL inst_cellmath__43_0_I1704 (.Y(N3218), .A0(N3176), .A1(N3173), .B0(N3175));
NAND2XL inst_cellmath__43_0_I1705 (.Y(N3219), .A(N3176), .B(N3174));
AOI21XL inst_cellmath__43_0_I1706 (.Y(N3220), .A0(N3180), .A1(N3177), .B0(N3179));
NAND2XL inst_cellmath__43_0_I1707 (.Y(N3221), .A(N3180), .B(N3178));
AOI21XL inst_cellmath__43_0_I1708 (.Y(N3222), .A0(N3184), .A1(N3181), .B0(N3183));
NAND2XL inst_cellmath__43_0_I1709 (.Y(N3223), .A(N3184), .B(N3182));
AOI21XL inst_cellmath__43_0_I1710 (.Y(N3224), .A0(N3188), .A1(N3185), .B0(N3187));
NAND2XL inst_cellmath__43_0_I1711 (.Y(N3225), .A(N3188), .B(N3186));
AOI21XL inst_cellmath__43_0_I1712 (.Y(N3226), .A0(N3192), .A1(N3189), .B0(N3191));
NAND2XL inst_cellmath__43_0_I1713 (.Y(N3227), .A(N3192), .B(N3190));
AOI21XL inst_cellmath__43_0_I1714 (.Y(N3228), .A0(N3196), .A1(N3193), .B0(N3195));
NAND2XL inst_cellmath__43_0_I1715 (.Y(N3229), .A(N3196), .B(N3194));
AOI21XL inst_cellmath__43_0_I1716 (.Y(N3230), .A0(N3200), .A1(N3197), .B0(N3199));
OAI21XL inst_cellmath__43_0_I1718 (.Y(N3232), .A0(N3205), .A1(N3202), .B0(N3204));
OAI21XL inst_cellmath__43_0_I1720 (.Y(N3234), .A0(N3209), .A1(N3206), .B0(N3208));
NOR2XL inst_cellmath__43_0_I1721 (.Y(N3235), .A(N3209), .B(N3207));
OAI21XL inst_cellmath__43_0_I1722 (.Y(N3236), .A0(N3213), .A1(N3210), .B0(N3212));
NOR2XL inst_cellmath__43_0_I1723 (.Y(N3237), .A(N3213), .B(N3211));
OAI21XL inst_cellmath__43_0_I1724 (.Y(N3238), .A0(N3217), .A1(N3214), .B0(N3216));
NOR2XL inst_cellmath__43_0_I1725 (.Y(N3239), .A(N3217), .B(N3215));
OAI21XL inst_cellmath__43_0_I1726 (.Y(N3240), .A0(N3221), .A1(N3218), .B0(N3220));
NOR2XL inst_cellmath__43_0_I1727 (.Y(N3241), .A(N3221), .B(N3219));
OAI21XL inst_cellmath__43_0_I1728 (.Y(N3242), .A0(N3225), .A1(N3222), .B0(N3224));
NOR2XL inst_cellmath__43_0_I1729 (.Y(N3243), .A(N3225), .B(N3223));
AOI21XL inst_cellmath__43_0_I1732 (.Y(N3246), .A0(N3235), .A1(N3232), .B0(N3234));
AOI21XL inst_cellmath__43_0_I1734 (.Y(N3248), .A0(N3239), .A1(N3236), .B0(N3238));
NAND2XL inst_cellmath__43_0_I1735 (.Y(N3249), .A(N3239), .B(N3237));
AOI21XL inst_cellmath__43_0_I1736 (.Y(N3250), .A0(N3243), .A1(N3240), .B0(N3242));
OAI21XL inst_cellmath__43_0_I1738 (.Y(N3252), .A0(N3249), .A1(N3246), .B0(N3248));
INVXL inst_cellmath__43_0_I1741 (.Y(N3255), .A(N3250));
AOI31X1 inst_cellmath__43_0_I2217 (.Y(N3256), .A0(N3243), .A1(N3241), .A2(N3252), .B0(N3255));
INVXL inst_cellmath__43_0_I1744 (.Y(N3258), .A(N3237));
INVXL inst_cellmath__43_0_I1745 (.Y(N3259), .A(N3236));
OAI21XL inst_cellmath__43_0_I1746 (.Y(N3260), .A0(N3258), .A1(N3246), .B0(N3259));
INVXL inst_cellmath__43_0_I2148 (.Y(N3742), .A(N3252));
AOI21XL inst_cellmath__43_0_I1750 (.Y(N3264), .A0(N3241), .A1(N3252), .B0(N3240));
INVXL inst_cellmath__43_0_I2149 (.Y(N3743), .A(N3256));
OA21X1 inst_cellmath__43_0_I1972 (.Y(N3269), .A0(N3229), .A1(N3226), .B0(N3228));
OAI31X1 inst_cellmath__43_0_I2218 (.Y(N3270), .A0(N3229), .A1(N3227), .A2(N3256), .B0(N3269));
INVXL inst_cellmath__43_0_I1758 (.Y(N3272), .A(N3207));
INVXL inst_cellmath__43_0_I1759 (.Y(N3273), .A(N3206));
AOI21XL inst_cellmath__43_0_I1760 (.Y(N3274), .A0(N3272), .A1(N3232), .B0(N3273));
INVXL inst_cellmath__43_0_I2150 (.Y(N3744), .A(N3246));
OAI21XL inst_cellmath__43_0_I1764 (.Y(N3278), .A0(N3211), .A1(N3246), .B0(N3210));
INVXL inst_cellmath__43_0_I2151 (.Y(N3745), .A(N3260));
INVXL inst_cellmath__43_0_I1768 (.Y(N3282), .A(N3215));
INVXL inst_cellmath__43_0_I1769 (.Y(N3283), .A(N3214));
AOI21XL inst_cellmath__43_0_I1770 (.Y(N3284), .A0(N3282), .A1(N3260), .B0(N3283));
INVXL inst_cellmath__43_0_I2152 (.Y(N3746), .A(N3742));
OAI21XL inst_cellmath__43_0_I1774 (.Y(N3288), .A0(N3219), .A1(N3742), .B0(N3218));
INVXL inst_cellmath__43_0_I2153 (.Y(N3747), .A(N3264));
OAI21XL inst_cellmath__43_0_I1778 (.Y(N3292), .A0(N3223), .A1(N3264), .B0(N3222));
INVXL inst_cellmath__43_0_I2154 (.Y(N3748), .A(N3743));
INVXL inst_cellmath__43_0_I1782 (.Y(N3296), .A(N3227));
INVXL inst_cellmath__43_0_I1783 (.Y(N3297), .A(N3226));
AOI21XL inst_cellmath__43_0_I1784 (.Y(N3298), .A0(N3296), .A1(N3743), .B0(N3297));
INVXL inst_cellmath__43_0_I2155 (.Y(N3749), .A(N3270));
INVXL inst_cellmath__43_0_I1789 (.Y(N3303), .A(N3230));
AOI31X1 inst_cellmath__43_0_I2191 (.Y(N3304), .A0(N3200), .A1(N3198), .A2(N3270), .B0(N3303));
INVXL inst_cellmath__43_0_I1792 (.Y(N3306), .A(N3146));
INVXL inst_cellmath__43_0_I1793 (.Y(N3307), .A(N3145));
OAI21XL inst_cellmath__43_0_I1794 (.Y(N3308), .A0(N3306), .A1(N3202), .B0(N3307));
AOI21XL inst_cellmath__43_0_I1798 (.Y(N3312), .A0(N3150), .A1(N3232), .B0(N3149));
INVXL inst_cellmath__43_0_I1802 (.Y(N3316), .A(N3154));
INVXL inst_cellmath__43_0_I1803 (.Y(N3317), .A(N3153));
OAI21XL inst_cellmath__43_0_I1804 (.Y(N3318), .A0(N3316), .A1(N3274), .B0(N3317));
AOI21XL inst_cellmath__43_0_I1808 (.Y(N3322), .A0(N3158), .A1(N3744), .B0(N3157));
AOI21XL inst_cellmath__43_0_I1812 (.Y(N3326), .A0(N3162), .A1(N3278), .B0(N3161));
INVXL inst_cellmath__43_0_I1816 (.Y(N3330), .A(N3166));
INVXL inst_cellmath__43_0_I1817 (.Y(N3331), .A(N3165));
OAI21XL inst_cellmath__43_0_I1818 (.Y(N3332), .A0(N3330), .A1(N3745), .B0(N3331));
INVXL inst_cellmath__43_0_I1822 (.Y(N3336), .A(N3170));
INVXL inst_cellmath__43_0_I1823 (.Y(N3337), .A(N3169));
OAI21XL inst_cellmath__43_0_I1824 (.Y(N3338), .A0(N3336), .A1(N3284), .B0(N3337));
AOI21XL inst_cellmath__43_0_I1828 (.Y(N3342), .A0(N3174), .A1(N3746), .B0(N3173));
AOI21XL inst_cellmath__43_0_I1832 (.Y(N3346), .A0(N3178), .A1(N3288), .B0(N3177));
AOI21XL inst_cellmath__43_0_I1836 (.Y(N3350), .A0(N3182), .A1(N3747), .B0(N3181));
AOI21XL inst_cellmath__43_0_I1840 (.Y(N3354), .A0(N3186), .A1(N3292), .B0(N3185));
INVXL inst_cellmath__43_0_I1844 (.Y(N3358), .A(N3190));
INVXL inst_cellmath__43_0_I1845 (.Y(N3359), .A(N3189));
OAI21XL inst_cellmath__43_0_I1846 (.Y(N3360), .A0(N3358), .A1(N3748), .B0(N3359));
INVXL inst_cellmath__43_0_I1850 (.Y(N3364), .A(N3194));
INVXL inst_cellmath__43_0_I1851 (.Y(N3365), .A(N3193));
OAI21XL inst_cellmath__43_0_I1852 (.Y(N3366), .A0(N3364), .A1(N3298), .B0(N3365));
INVXL inst_cellmath__43_0_I1856 (.Y(N3370), .A(N3198));
INVXL inst_cellmath__43_0_I1857 (.Y(N3371), .A(N3197));
OAI21XL inst_cellmath__43_0_I1858 (.Y(N3372), .A0(N3370), .A1(N3749), .B0(N3371));
OR2XL inst_cellmath__43_0_I1864 (.Y(inst_cellmath__43_0_out0[47]), .A(N3376), .B(N3304));
XNOR2X1 inst_cellmath__43_0_I1870 (.Y(inst_cellmath__43_0_out0[17]), .A(N3141), .B(N3144));
XOR2XL inst_cellmath__43_0_I1871 (.Y(inst_cellmath__43_0_out0[18]), .A(N3202), .B(N3146));
XNOR2X1 inst_cellmath__43_0_I1872 (.Y(inst_cellmath__43_0_out0[19]), .A(N3308), .B(N3148));
XNOR2X1 inst_cellmath__43_0_I1873 (.Y(inst_cellmath__43_0_out0[20]), .A(N3232), .B(N3150));
XOR2XL inst_cellmath__43_0_I1874 (.Y(inst_cellmath__43_0_out0[21]), .A(N3312), .B(N3152));
XOR2XL inst_cellmath__43_0_I2192 (.Y(inst_cellmath__43_0_out0[22]), .A(N3274), .B(N3154));
XNOR2X1 inst_cellmath__43_0_I1876 (.Y(inst_cellmath__43_0_out0[23]), .A(N3318), .B(N3156));
XNOR2X1 inst_cellmath__43_0_I1877 (.Y(inst_cellmath__43_0_out0[24]), .A(N3744), .B(N3158));
XOR2XL inst_cellmath__43_0_I1878 (.Y(inst_cellmath__43_0_out0[25]), .A(N3322), .B(N3160));
XNOR2X1 inst_cellmath__43_0_I1879 (.Y(inst_cellmath__43_0_out0[26]), .A(N3278), .B(N3162));
XOR2XL inst_cellmath__43_0_I1880 (.Y(inst_cellmath__43_0_out0[27]), .A(N3326), .B(N3164));
XOR2XL inst_cellmath__43_0_I2193 (.Y(inst_cellmath__43_0_out0[28]), .A(N3745), .B(N3166));
XNOR2X1 inst_cellmath__43_0_I1882 (.Y(inst_cellmath__43_0_out0[29]), .A(N3332), .B(N3168));
XOR2XL inst_cellmath__43_0_I2194 (.Y(inst_cellmath__43_0_out0[30]), .A(N3284), .B(N3170));
XNOR2X1 inst_cellmath__43_0_I1884 (.Y(inst_cellmath__43_0_out0[31]), .A(N3338), .B(N3172));
XNOR2X1 inst_cellmath__43_0_I1885 (.Y(inst_cellmath__43_0_out0[32]), .A(N3746), .B(N3174));
XOR2XL inst_cellmath__43_0_I1886 (.Y(inst_cellmath__43_0_out0[33]), .A(N3342), .B(N3176));
XNOR2X1 inst_cellmath__43_0_I1887 (.Y(inst_cellmath__43_0_out0[34]), .A(N3288), .B(N3178));
XOR2XL inst_cellmath__43_0_I1888 (.Y(inst_cellmath__43_0_out0[35]), .A(N3346), .B(N3180));
XNOR2X1 inst_cellmath__43_0_I1889 (.Y(inst_cellmath__43_0_out0[36]), .A(N3747), .B(N3182));
XOR2XL inst_cellmath__43_0_I1890 (.Y(inst_cellmath__43_0_out0[37]), .A(N3350), .B(N3184));
XNOR2X1 inst_cellmath__43_0_I1891 (.Y(inst_cellmath__43_0_out0[38]), .A(N3292), .B(N3186));
XOR2XL inst_cellmath__43_0_I1892 (.Y(inst_cellmath__43_0_out0[39]), .A(N3354), .B(N3188));
XOR2XL inst_cellmath__43_0_I2195 (.Y(inst_cellmath__43_0_out0[40]), .A(N3748), .B(N3190));
XNOR2X1 inst_cellmath__43_0_I1894 (.Y(inst_cellmath__43_0_out0[41]), .A(N3360), .B(N3192));
XOR2XL inst_cellmath__43_0_I2196 (.Y(inst_cellmath__43_0_out0[42]), .A(N3298), .B(N3194));
XNOR2X1 inst_cellmath__43_0_I1896 (.Y(inst_cellmath__43_0_out0[43]), .A(N3366), .B(N3196));
XOR2XL inst_cellmath__43_0_I2197 (.Y(inst_cellmath__43_0_out0[44]), .A(N3749), .B(N3198));
XNOR2X1 inst_cellmath__43_0_I1898 (.Y(inst_cellmath__43_0_out0[45]), .A(N3372), .B(N3200));
XNOR2X1 inst_cellmath__43_0_I1899 (.Y(inst_cellmath__43_0_out0[46]), .A(N3304), .B(N3376));
endmodule

module cynw_cm_float_mul_inst_cellmath__30__13__bdw3636473930_bdw (
	inst_cellmath__30__13__out0,
	inst_cellmath__30__13__in0,
	inst_cellmath__30__13__in1,
	inst_cellmath__30__13__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__30__13__out0;
input  inst_cellmath__30__13__in0,
	inst_cellmath__30__13__in1,
	inst_cellmath__30__13__in2;
wire N6;
NOR2XL inst_cellmath__30__13__I0 (.Y(N6), .A(inst_cellmath__30__13__in0), .B(inst_cellmath__30__13__in2));
AND2XL inst_cellmath__30__13__I1 (.Y(inst_cellmath__30__13__out0[0]), .A(N6), .B(inst_cellmath__30__13__in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__30__14__bdw3636473930_bdw (
	inst_cellmath__30__14__out0,
	inst_cellmath__30__14__in0,
	inst_cellmath__30__14__in1,
	inst_cellmath__30__14__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__30__14__out0;
input  inst_cellmath__30__14__in0,
	inst_cellmath__30__14__in1,
	inst_cellmath__30__14__in2;
wire N6;
NOR2XL inst_cellmath__30__14__I0 (.Y(N6), .A(inst_cellmath__30__14__in0), .B(inst_cellmath__30__14__in2));
AND2XL inst_cellmath__30__14__I1 (.Y(inst_cellmath__30__14__out0[0]), .A(N6), .B(inst_cellmath__30__14__in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__30_0_bdw3636473930_bdw (
	inst_cellmath__30_0_out0,
	inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__30_0_out0;
input [0:0] inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1;
OR2XL inst_cellmath__30_0_I0 (.Y(inst_cellmath__30_0_out0), .A(inst_cellmath__30_0_in1[0]), .B(inst_cellmath__30_0_in0[0]));
endmodule

module cynw_cm_float_mul_inst_cellmath__34_0_bdw3636473930_bdw (
	inst_cellmath__34_0_out0,
	inst_cellmath__34_0_in0,
	inst_cellmath__34_0_in1
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__34_0_out0;
input [7:0] inst_cellmath__34_0_in0,
	inst_cellmath__34_0_in1;
wire N106,N111,N115,N117,N119,N121,N123 
	,N125,N127;
INVXL inst_cellmath__34_0_I40 (.Y(N106), .A(inst_cellmath__34_0_in1[7]));
XNOR2X1 hap1_A_I54 (.Y(inst_cellmath__34_0_out0[0]), .A(inst_cellmath__34_0_in0[0]), .B(inst_cellmath__34_0_in1[0]));
OR2XL hap1_A_I55 (.Y(N111), .A(inst_cellmath__34_0_in0[0]), .B(inst_cellmath__34_0_in1[0]));
ADDFX1 inst_cellmath__34_0_I42 (.CO(N115), .S(inst_cellmath__34_0_out0[1]), .A(inst_cellmath__34_0_in0[1]), .B(inst_cellmath__34_0_in1[1]), .CI(N111));
ADDFX1 inst_cellmath__34_0_I43 (.CO(N117), .S(inst_cellmath__34_0_out0[2]), .A(inst_cellmath__34_0_in0[2]), .B(inst_cellmath__34_0_in1[2]), .CI(N115));
ADDFX1 inst_cellmath__34_0_I44 (.CO(N119), .S(inst_cellmath__34_0_out0[3]), .A(inst_cellmath__34_0_in0[3]), .B(inst_cellmath__34_0_in1[3]), .CI(N117));
ADDFX1 inst_cellmath__34_0_I45 (.CO(N121), .S(inst_cellmath__34_0_out0[4]), .A(inst_cellmath__34_0_in0[4]), .B(inst_cellmath__34_0_in1[4]), .CI(N119));
ADDFX1 inst_cellmath__34_0_I46 (.CO(N123), .S(inst_cellmath__34_0_out0[5]), .A(inst_cellmath__34_0_in0[5]), .B(inst_cellmath__34_0_in1[5]), .CI(N121));
ADDFX1 inst_cellmath__34_0_I47 (.CO(N125), .S(inst_cellmath__34_0_out0[6]), .A(inst_cellmath__34_0_in0[6]), .B(inst_cellmath__34_0_in1[6]), .CI(N123));
ADDFX1 inst_cellmath__34_0_I48 (.CO(N127), .S(inst_cellmath__34_0_out0[7]), .A(N106), .B(inst_cellmath__34_0_in0[7]), .CI(N125));
XNOR2X1 hap1_A_I56 (.Y(inst_cellmath__34_0_out0[8]), .A(inst_cellmath__34_0_in1[7]), .B(N127));
NOR2XL hap1_A_I57 (.Y(inst_cellmath__34_0_out0[9]), .A(inst_cellmath__34_0_in1[7]), .B(N127));
endmodule

module cynw_cm_float_mul_inst_cellmath__41__24__bdw3636473930_bdw (
	inst_cellmath__41__24__out0,
	inst_cellmath__41__24__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__41__24__out0;
input [7:0] inst_cellmath__41__24__in0;
wire N15,N20,N46;
AND4XL inst_cellmath__41__24__I14 (.Y(N15), .A(inst_cellmath__41__24__in0[0]), .B(inst_cellmath__41__24__in0[1]), .C(inst_cellmath__41__24__in0[2]), .D(inst_cellmath__41__24__in0[3]));
NAND3XL inst_cellmath__41__24__I15 (.Y(N20), .A(inst_cellmath__41__24__in0[4]), .B(inst_cellmath__41__24__in0[7]), .C(inst_cellmath__41__24__in0[5]));
NAND2XL hyperpropagate_3_1_A_I17 (.Y(N46), .A(inst_cellmath__41__24__in0[6]), .B(N15));
NOR2XL hyperpropagate_3_1_A_I18 (.Y(inst_cellmath__41__24__out0[0]), .A(N20), .B(N46));
endmodule

module cynw_cm_float_mul_inst_cellmath__41__23__bdw3636473930_bdw (
	inst_cellmath__41__23__out0,
	inst_cellmath__41__23__in0,
	inst_cellmath__41__23__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__41__23__out0;
input [0:0] inst_cellmath__41__23__in0;
input [8:8] inst_cellmath__41__23__in1;
OR2XL inst_cellmath__41__23__I0 (.Y(inst_cellmath__41__23__out0[0]), .A(inst_cellmath__41__23__in1[8]), .B(inst_cellmath__41__23__in0[0]));
endmodule

module cynw_cm_float_mul_inst_cellmath__41_0_bdw3636473930_bdw (
	inst_cellmath__41_0_out0,
	inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__41_0_out0;
input [0:0] inst_cellmath__41_0_in0;
input [9:9] inst_cellmath__41_0_in1;
NOR2BX1 inst_cellmath__41_0_I3 (.Y(inst_cellmath__41_0_out0), .AN(inst_cellmath__41_0_in0[0]), .B(inst_cellmath__41_0_in1[9]));
endmodule

module cynw_cm_float_mul_inst_cellmath__37_0_bdw3636473930_bdw (
	inst_cellmath__37_0_out0,
	inst_cellmath__37_0_in0,
	inst_cellmath__37_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__37_0_out0;
input  inst_cellmath__37_0_in0,
	inst_cellmath__37_0_in1;
OR2XL inst_cellmath__37_0_I0 (.Y(inst_cellmath__37_0_out0), .A(inst_cellmath__37_0_in1), .B(inst_cellmath__37_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__35__16__bdw3636473930_bdw (
	inst_cellmath__35__16__out0,
	inst_cellmath__35__16__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__35__16__out0;
input [9:0] inst_cellmath__35__16__in0;
wire N14,N20,N21,N23;
NOR2XL inst_cellmath__35__16__I0 (.Y(N14), .A(inst_cellmath__35__16__in0[0]), .B(inst_cellmath__35__16__in0[9]));
NOR4BX1 inst_cellmath__35__16__I79 (.Y(N20), .AN(N14), .B(inst_cellmath__35__16__in0[1]), .C(inst_cellmath__35__16__in0[8]), .D(inst_cellmath__35__16__in0[2]));
NOR2XL inst_cellmath__35__16__I8 (.Y(N21), .A(inst_cellmath__35__16__in0[7]), .B(inst_cellmath__35__16__in0[6]));
OR3XL inst_cellmath__35__16__I78 (.Y(N23), .A(inst_cellmath__35__16__in0[3]), .B(inst_cellmath__35__16__in0[4]), .C(inst_cellmath__35__16__in0[5]));
NAND3BXL inst_cellmath__35__16__I76 (.Y(inst_cellmath__35__16__out0[0]), .AN(N23), .B(N21), .C(N20));
endmodule

module cynw_cm_float_mul_inst_cellmath__32__11__bdw3636473930_bdw (
	inst_cellmath__32__11__out0,
	inst_cellmath__32__11__in0,
	inst_cellmath__32__11__in1,
	inst_cellmath__32__11__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__32__11__out0;
input  inst_cellmath__32__11__in0,
	inst_cellmath__32__11__in1,
	inst_cellmath__32__11__in2;
NOR3BXL inst_cellmath__32__11__I5 (.Y(inst_cellmath__32__11__out0[0]), .AN(inst_cellmath__32__11__in0), .B(inst_cellmath__32__11__in2), .C(inst_cellmath__32__11__in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__32__12__bdw3636473930_bdw (
	inst_cellmath__32__12__out0,
	inst_cellmath__32__12__in0,
	inst_cellmath__32__12__in1,
	inst_cellmath__32__12__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__32__12__out0;
input  inst_cellmath__32__12__in0,
	inst_cellmath__32__12__in1,
	inst_cellmath__32__12__in2;
NOR3BXL inst_cellmath__32__12__I5 (.Y(inst_cellmath__32__12__out0[0]), .AN(inst_cellmath__32__12__in0), .B(inst_cellmath__32__12__in2), .C(inst_cellmath__32__12__in1));
endmodule

module cynw_cm_float_mul_inst_cellmath__32_0_bdw3636473930_bdw (
	inst_cellmath__32_0_out0,
	inst_cellmath__32_0_in0,
	inst_cellmath__32_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__32_0_out0;
input [0:0] inst_cellmath__32_0_in0,
	inst_cellmath__32_0_in1;
OR2XL inst_cellmath__32_0_I0 (.Y(inst_cellmath__32_0_out0), .A(inst_cellmath__32_0_in1[0]), .B(inst_cellmath__32_0_in0[0]));
endmodule

module cynw_cm_float_mul_inst_cellmath__60_0_bdw3636473930_bdw (
	inst_cellmath__60_0_out0,
	inst_cellmath__60_0_in0,
	inst_cellmath__60_0_in1,
	inst_cellmath__60_0_in2,
	inst_cellmath__60_0_in3,
	inst_cellmath__60_0_in4
	); /* architecture "gate_level" */ 
output  inst_cellmath__60_0_out0;
input  inst_cellmath__60_0_in0;
input [0:0] inst_cellmath__60_0_in1;
input [9:9] inst_cellmath__60_0_in2;
input  inst_cellmath__60_0_in3,
	inst_cellmath__60_0_in4;
wire N10,N11;
NOR3XL inst_cellmath__60_0_I6 (.Y(N10), .A(inst_cellmath__60_0_in3), .B(inst_cellmath__60_0_in4), .C(inst_cellmath__60_0_in2[9]));
NAND2XL inst_cellmath__60_0_I3 (.Y(N11), .A(N10), .B(inst_cellmath__60_0_in1[0]));
OR2XL inst_cellmath__60_0_I4 (.Y(inst_cellmath__60_0_out0), .A(N11), .B(inst_cellmath__60_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__42__22__bdw3636473930_bdw (
	inst_cellmath__42__22__out0,
	inst_cellmath__42__22__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__42__22__out0;
input [7:1] inst_cellmath__42__22__in0;
wire N11,N12,N13,N15,N16,N43;
NAND2XL inst_cellmath__42__22__I0 (.Y(N13), .A(inst_cellmath__42__22__in0[1]), .B(inst_cellmath__42__22__in0[2]));
NAND2XL inst_cellmath__42__22__I1 (.Y(N11), .A(inst_cellmath__42__22__in0[3]), .B(inst_cellmath__42__22__in0[4]));
NAND2XL inst_cellmath__42__22__I2 (.Y(N12), .A(inst_cellmath__42__22__in0[7]), .B(inst_cellmath__42__22__in0[6]));
INVXL inst_cellmath__42__22__I16 (.Y(N43), .A(inst_cellmath__42__22__in0[5]));
NOR2XL inst_cellmath__42__22__I4 (.Y(N16), .A(N13), .B(N43));
NOR2XL inst_cellmath__42__22__I5 (.Y(N15), .A(N11), .B(N12));
AND2XL inst_cellmath__42__22__I7 (.Y(inst_cellmath__42__22__out0[0]), .A(N16), .B(N15));
endmodule

module cynw_cm_float_mul_inst_cellmath__42__21__bdw3636473930_bdw (
	inst_cellmath__42__21__out0,
	inst_cellmath__42__21__in0,
	inst_cellmath__42__21__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__42__21__out0;
input [0:0] inst_cellmath__42__21__in0;
input [8:8] inst_cellmath__42__21__in1;
OR2XL inst_cellmath__42__21__I0 (.Y(inst_cellmath__42__21__out0[0]), .A(inst_cellmath__42__21__in1[8]), .B(inst_cellmath__42__21__in0[0]));
endmodule

module cynw_cm_float_mul_inst_cellmath__42_0_bdw3636473930_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__42_0_out0;
input [0:0] inst_cellmath__42_0_in0;
input [9:9] inst_cellmath__42_0_in1;
NOR2BX1 inst_cellmath__42_0_I3 (.Y(inst_cellmath__42_0_out0), .AN(inst_cellmath__42_0_in0[0]), .B(inst_cellmath__42_0_in1[9]));
endmodule

module cynw_cm_float_mul_inst_cellmath__38_0_bdw3636473930_bdw (
	inst_cellmath__38_0_out0,
	inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__38_0_out0;
input  inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1;
OR2XL inst_cellmath__38_0_I0 (.Y(inst_cellmath__38_0_out0), .A(inst_cellmath__38_0_in1), .B(inst_cellmath__38_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__61_0_bdw3636473930_bdw (
	inst_cellmath__61_0_out0,
	inst_cellmath__61_0_in0,
	inst_cellmath__61_0_in1,
	inst_cellmath__61_0_in2,
	inst_cellmath__61_0_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__61_0_out0;
input  inst_cellmath__61_0_in0;
input [9:9] inst_cellmath__61_0_in1;
input  inst_cellmath__61_0_in2,
	inst_cellmath__61_0_in3;
OR4X1 inst_cellmath__61_0_I7 (.Y(inst_cellmath__61_0_out0), .A(inst_cellmath__61_0_in2), .B(inst_cellmath__61_0_in3), .C(inst_cellmath__61_0_in1[9]), .D(inst_cellmath__61_0_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__56_1_bdw3636473930_bdw (
	inst_cellmath__56_1_out0,
	inst_cellmath__56_1_in0,
	inst_cellmath__56_1_in1,
	inst_cellmath__56_1_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__56_1_out0;
input  inst_cellmath__56_1_in0,
	inst_cellmath__56_1_in1;
input [47:47] inst_cellmath__56_1_in2;
MX2XL inst_cellmath__56_1_I2 (.Y(inst_cellmath__56_1_out0), .A(inst_cellmath__56_1_in1), .B(inst_cellmath__56_1_in0), .S0(inst_cellmath__56_1_in2[47]));
endmodule

module cynw_cm_float_mul_inst_cellmath__50_0_bdw3636473930_bdw (
	inst_cellmath__50_0_out0,
	inst_cellmath__50_0_in0
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__50_0_out0;
input [7:0] inst_cellmath__50_0_in0;
wire N87,N90,N97,N102,N112,N173,N175 
	,N179;
INVXL inst_cellmath__50_0_I91 (.Y(inst_cellmath__50_0_out0[0]), .A(inst_cellmath__50_0_in0[0]));
NOR2BX1 inst_cellmath__50_0_I153 (.Y(N87), .AN(inst_cellmath__50_0_in0[1]), .B(inst_cellmath__50_0_out0[0]));
XNOR2X1 inst_cellmath__50_0_I40 (.Y(inst_cellmath__50_0_out0[1]), .A(inst_cellmath__50_0_out0[0]), .B(inst_cellmath__50_0_in0[1]));
NAND2XL inst_cellmath__50_0_I43 (.Y(N90), .A(inst_cellmath__50_0_in0[2]), .B(N87));
INVXL inst_cellmath__50_0_I92 (.Y(N175), .A(inst_cellmath__50_0_in0[4]));
INVXL inst_cellmath__50_0_I90 (.Y(N173), .A(inst_cellmath__50_0_in0[3]));
NOR3XL inst_cellmath__50_0_I96 (.Y(N97), .A(N175), .B(N173), .C(N90));
NAND3XL inst_cellmath__50_0_I154 (.Y(N102), .A(inst_cellmath__50_0_in0[5]), .B(N97), .C(inst_cellmath__50_0_in0[6]));
NAND2XL inst_cellmath__50_0_I61 (.Y(N112), .A(inst_cellmath__50_0_in0[5]), .B(N97));
XOR2XL inst_cellmath__50_0_I73 (.Y(inst_cellmath__50_0_out0[2]), .A(N87), .B(inst_cellmath__50_0_in0[2]));
XOR2XL inst_cellmath__50_0_I74 (.Y(inst_cellmath__50_0_out0[3]), .A(N90), .B(N173));
NOR2XL node_cs_const1_cs_A_I109 (.Y(N179), .A(N173), .B(N90));
XNOR2X1 node_cs_const1_cs_A_I110 (.Y(inst_cellmath__50_0_out0[4]), .A(N175), .B(N179));
XOR2XL inst_cellmath__50_0_I155 (.Y(inst_cellmath__50_0_out0[5]), .A(N97), .B(inst_cellmath__50_0_in0[5]));
XNOR2X1 inst_cellmath__50_0_I77 (.Y(inst_cellmath__50_0_out0[6]), .A(N112), .B(inst_cellmath__50_0_in0[6]));
XNOR2X1 inst_cellmath__50_0_I78 (.Y(inst_cellmath__50_0_out0[7]), .A(N102), .B(inst_cellmath__50_0_in0[7]));
endmodule

module cynw_cm_float_mul_inst_cellmath__54_7_bdw3636473930_bdw (
	inst_cellmath__54_7_out0,
	inst_cellmath__54_7_in0,
	inst_cellmath__54_7_in1,
	inst_cellmath__54_7_in2
	); /* architecture "gate_level" */ 
output [7:7] inst_cellmath__54_7_out0;
input  inst_cellmath__54_7_in0,
	inst_cellmath__54_7_in1,
	inst_cellmath__54_7_in2;
OR3XL inst_cellmath__54_7_I6 (.Y(inst_cellmath__54_7_out0[7]), .A(inst_cellmath__54_7_in2), .B(inst_cellmath__54_7_in1), .C(inst_cellmath__54_7_in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__54__30__bdw3636473930_bdw (
	inst_cellmath__54__30__out0,
	inst_cellmath__54__30__in0,
	inst_cellmath__54__30__in1,
	inst_cellmath__54__30__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__54__30__out0;
input  inst_cellmath__54__30__in0,
	inst_cellmath__54__30__in1,
	inst_cellmath__54__30__in2;
OR3XL inst_cellmath__54__30__I6 (.Y(inst_cellmath__54__30__out0[0]), .A(inst_cellmath__54__30__in2), .B(inst_cellmath__54__30__in1), .C(inst_cellmath__54__30__in0));
endmodule

module cynw_cm_float_mul_inst_cellmath__64_2WWMM_bdw3636473930_bdw (
	inst_cellmath__64_2WWMM_out0,
	inst_cellmath__64_2WWMM_in0,
	inst_cellmath__64_2WWMM_in1,
	inst_cellmath__64_2WWMM_in2,
	inst_cellmath__64_2WWMM_in3,
	inst_cellmath__64_2WWMM_in4,
	inst_cellmath__64_2WWMM_in5,
	inst_cellmath__64_2WWMM_in6
	); /* architecture "gate_level" */ 
output [30:0] inst_cellmath__64_2WWMM_out0;
input  inst_cellmath__64_2WWMM_in0;
input [0:0] inst_cellmath__64_2WWMM_in1;
input [7:7] inst_cellmath__64_2WWMM_in2;
input [7:0] inst_cellmath__64_2WWMM_in3;
input [47:23] inst_cellmath__64_2WWMM_in4;
input [7:0] inst_cellmath__64_2WWMM_in5;
input  inst_cellmath__64_2WWMM_in6;
wire N157,N159,N161,N163,N165,N167,N169 
	,N171,N173,N175,N177,N179,N181,N183,N185 
	,N187,N189,N191,N193,N195,N197,N199,N201 
	,N203,N205,N207,N209,N211,N213,N215,N217 
	,N317,N348,N359,N367;
NOR2X1 inst_cellmath__64_2WWMM_I146 (.Y(N348), .A(inst_cellmath__64_2WWMM_in4[47]), .B(inst_cellmath__64_2WWMM_in0));
NOR2BX1 inst_cellmath__64_2WWMM_I147 (.Y(N317), .AN(inst_cellmath__64_2WWMM_in4[47]), .B(inst_cellmath__64_2WWMM_in0));
AOI22XL inst_cellmath__64_2WWMM_I6 (.Y(N157), .A0(inst_cellmath__64_2WWMM_in3[0]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[0]));
AOI22XL inst_cellmath__64_2WWMM_I7 (.Y(N159), .A0(inst_cellmath__64_2WWMM_in3[1]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[1]));
AOI22XL inst_cellmath__64_2WWMM_I8 (.Y(N161), .A0(inst_cellmath__64_2WWMM_in3[2]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[2]));
AOI22XL inst_cellmath__64_2WWMM_I9 (.Y(N163), .A0(inst_cellmath__64_2WWMM_in3[3]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[3]));
AOI22XL inst_cellmath__64_2WWMM_I10 (.Y(N165), .A0(inst_cellmath__64_2WWMM_in3[4]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[4]));
AOI22XL inst_cellmath__64_2WWMM_I11 (.Y(N167), .A0(inst_cellmath__64_2WWMM_in3[5]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[5]));
AOI22XL inst_cellmath__64_2WWMM_I12 (.Y(N169), .A0(inst_cellmath__64_2WWMM_in3[6]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[6]));
AOI22XL inst_cellmath__64_2WWMM_I13 (.Y(N171), .A0(inst_cellmath__64_2WWMM_in3[7]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in5[7]));
AOI22XL inst_cellmath__64_2WWMM_I14 (.Y(N173), .A0(inst_cellmath__64_2WWMM_in4[24]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[23]));
AOI22XL inst_cellmath__64_2WWMM_I15 (.Y(N175), .A0(inst_cellmath__64_2WWMM_in4[25]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[24]));
AOI22XL inst_cellmath__64_2WWMM_I16 (.Y(N177), .A0(inst_cellmath__64_2WWMM_in4[26]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[25]));
AOI22XL inst_cellmath__64_2WWMM_I17 (.Y(N179), .A0(inst_cellmath__64_2WWMM_in4[27]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[26]));
AOI22XL inst_cellmath__64_2WWMM_I18 (.Y(N181), .A0(inst_cellmath__64_2WWMM_in4[28]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[27]));
AOI22XL inst_cellmath__64_2WWMM_I19 (.Y(N183), .A0(inst_cellmath__64_2WWMM_in4[29]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[28]));
AOI22XL inst_cellmath__64_2WWMM_I20 (.Y(N185), .A0(inst_cellmath__64_2WWMM_in4[30]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[29]));
AOI22XL inst_cellmath__64_2WWMM_I21 (.Y(N187), .A0(inst_cellmath__64_2WWMM_in4[31]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[30]));
AOI22XL inst_cellmath__64_2WWMM_I22 (.Y(N189), .A0(inst_cellmath__64_2WWMM_in4[32]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[31]));
AOI22XL inst_cellmath__64_2WWMM_I23 (.Y(N191), .A0(inst_cellmath__64_2WWMM_in4[33]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[32]));
AOI22XL inst_cellmath__64_2WWMM_I24 (.Y(N193), .A0(inst_cellmath__64_2WWMM_in4[34]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[33]));
AOI22XL inst_cellmath__64_2WWMM_I25 (.Y(N195), .A0(inst_cellmath__64_2WWMM_in4[35]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[34]));
AOI22XL inst_cellmath__64_2WWMM_I26 (.Y(N197), .A0(inst_cellmath__64_2WWMM_in4[36]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[35]));
AOI22XL inst_cellmath__64_2WWMM_I27 (.Y(N199), .A0(inst_cellmath__64_2WWMM_in4[37]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[36]));
AOI22XL inst_cellmath__64_2WWMM_I28 (.Y(N201), .A0(inst_cellmath__64_2WWMM_in4[38]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[37]));
AOI22XL inst_cellmath__64_2WWMM_I29 (.Y(N203), .A0(inst_cellmath__64_2WWMM_in4[39]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[38]));
AOI22XL inst_cellmath__64_2WWMM_I30 (.Y(N205), .A0(inst_cellmath__64_2WWMM_in4[40]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[39]));
AOI22XL inst_cellmath__64_2WWMM_I31 (.Y(N207), .A0(inst_cellmath__64_2WWMM_in4[41]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[40]));
AOI22XL inst_cellmath__64_2WWMM_I32 (.Y(N209), .A0(inst_cellmath__64_2WWMM_in4[42]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[41]));
AOI22XL inst_cellmath__64_2WWMM_I33 (.Y(N211), .A0(inst_cellmath__64_2WWMM_in4[43]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[42]));
AOI22XL inst_cellmath__64_2WWMM_I34 (.Y(N213), .A0(inst_cellmath__64_2WWMM_in4[44]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[43]));
AOI22XL inst_cellmath__64_2WWMM_I35 (.Y(N215), .A0(inst_cellmath__64_2WWMM_in4[45]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[44]));
AOI22XL inst_cellmath__64_2WWMM_I36 (.Y(N217), .A0(inst_cellmath__64_2WWMM_in4[46]), .A1(N317), .B0(N348), .B1(inst_cellmath__64_2WWMM_in4[45]));
NAND2XL inst_cellmath__64_2WWMM_I149 (.Y(N359), .A(inst_cellmath__64_2WWMM_in0), .B(inst_cellmath__64_2WWMM_in1[0]));
NAND2X1 inst_cellmath__64_2WWMM_I155 (.Y(N367), .A(inst_cellmath__64_2WWMM_in0), .B(inst_cellmath__64_2WWMM_in6));
NAND2XL inst_cellmath__64_2WWMM_I71 (.Y(inst_cellmath__64_2WWMM_out0[0]), .A(N359), .B(N157));
NAND2XL inst_cellmath__64_2WWMM_I72 (.Y(inst_cellmath__64_2WWMM_out0[1]), .A(N359), .B(N159));
NAND2XL inst_cellmath__64_2WWMM_I73 (.Y(inst_cellmath__64_2WWMM_out0[2]), .A(N359), .B(N161));
NAND2XL inst_cellmath__64_2WWMM_I74 (.Y(inst_cellmath__64_2WWMM_out0[3]), .A(N359), .B(N163));
NAND2XL inst_cellmath__64_2WWMM_I75 (.Y(inst_cellmath__64_2WWMM_out0[4]), .A(N359), .B(N165));
NAND2XL inst_cellmath__64_2WWMM_I76 (.Y(inst_cellmath__64_2WWMM_out0[5]), .A(N359), .B(N167));
NAND2XL inst_cellmath__64_2WWMM_I77 (.Y(inst_cellmath__64_2WWMM_out0[6]), .A(N359), .B(N169));
OAI2BB1X1 inst_cellmath__64_2WWMM_I152 (.Y(inst_cellmath__64_2WWMM_out0[7]), .A0N(inst_cellmath__64_2WWMM_in0), .A1N(inst_cellmath__64_2WWMM_in2[7]), .B0(N171));
NAND2XL inst_cellmath__64_2WWMM_I79 (.Y(inst_cellmath__64_2WWMM_out0[8]), .A(N367), .B(N173));
NAND2XL inst_cellmath__64_2WWMM_I80 (.Y(inst_cellmath__64_2WWMM_out0[9]), .A(N367), .B(N175));
NAND2XL inst_cellmath__64_2WWMM_I81 (.Y(inst_cellmath__64_2WWMM_out0[10]), .A(N367), .B(N177));
NAND2XL inst_cellmath__64_2WWMM_I82 (.Y(inst_cellmath__64_2WWMM_out0[11]), .A(N367), .B(N179));
NAND2XL inst_cellmath__64_2WWMM_I83 (.Y(inst_cellmath__64_2WWMM_out0[12]), .A(N367), .B(N181));
NAND2XL inst_cellmath__64_2WWMM_I84 (.Y(inst_cellmath__64_2WWMM_out0[13]), .A(N367), .B(N183));
NAND2XL inst_cellmath__64_2WWMM_I85 (.Y(inst_cellmath__64_2WWMM_out0[14]), .A(N367), .B(N185));
NAND2XL inst_cellmath__64_2WWMM_I86 (.Y(inst_cellmath__64_2WWMM_out0[15]), .A(N367), .B(N187));
NAND2XL inst_cellmath__64_2WWMM_I87 (.Y(inst_cellmath__64_2WWMM_out0[16]), .A(N367), .B(N189));
NAND2XL inst_cellmath__64_2WWMM_I88 (.Y(inst_cellmath__64_2WWMM_out0[17]), .A(N367), .B(N191));
NAND2XL inst_cellmath__64_2WWMM_I89 (.Y(inst_cellmath__64_2WWMM_out0[18]), .A(N367), .B(N193));
NAND2XL inst_cellmath__64_2WWMM_I90 (.Y(inst_cellmath__64_2WWMM_out0[19]), .A(N367), .B(N195));
NAND2XL inst_cellmath__64_2WWMM_I91 (.Y(inst_cellmath__64_2WWMM_out0[20]), .A(N367), .B(N197));
NAND2XL inst_cellmath__64_2WWMM_I92 (.Y(inst_cellmath__64_2WWMM_out0[21]), .A(N367), .B(N199));
NAND2XL inst_cellmath__64_2WWMM_I93 (.Y(inst_cellmath__64_2WWMM_out0[22]), .A(N367), .B(N201));
NAND2XL inst_cellmath__64_2WWMM_I94 (.Y(inst_cellmath__64_2WWMM_out0[23]), .A(N367), .B(N203));
NAND2XL inst_cellmath__64_2WWMM_I95 (.Y(inst_cellmath__64_2WWMM_out0[24]), .A(N367), .B(N205));
NAND2XL inst_cellmath__64_2WWMM_I96 (.Y(inst_cellmath__64_2WWMM_out0[25]), .A(N367), .B(N207));
NAND2XL inst_cellmath__64_2WWMM_I97 (.Y(inst_cellmath__64_2WWMM_out0[26]), .A(N367), .B(N209));
NAND2XL inst_cellmath__64_2WWMM_I98 (.Y(inst_cellmath__64_2WWMM_out0[27]), .A(N367), .B(N211));
NAND2XL inst_cellmath__64_2WWMM_I99 (.Y(inst_cellmath__64_2WWMM_out0[28]), .A(N367), .B(N213));
NAND2XL inst_cellmath__64_2WWMM_I100 (.Y(inst_cellmath__64_2WWMM_out0[29]), .A(N367), .B(N215));
NAND2XL inst_cellmath__64_2WWMM_I101 (.Y(inst_cellmath__64_2WWMM_out0[30]), .A(N367), .B(N217));
endmodule

/* CADENCE  urn2Qw/arRs= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




module DFT_compute_cynw_cm_float_mul_E8_M23_2( a_sign, a_exp, a_man, b_sign, b_exp, b_man, x, aclk, astall );
input a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
wire[31:0] x_wire;
input aclk;
input astall;
cynw_cm_float_mul_inst_cellmath__64_2WWMM_bdw3636473930_bdw cynw_cm_float_mul_inst_cellmath__64_2WWMM_bdw1103716848_bdw_inst( .a_sign(a_sign), .a_exp(a_exp), .a_man(a_man), .b_sign(b_sign), .b_exp(b_exp), .b_man(b_man), .x(x_wire));
reg [31:0] x_reg_0;
/* $A : movable_reg */
always @(posedge aclk) begin
    if ( !astall) x_reg_0 <= x_wire;
end
/* $A : movable_reg = reset */
assign x = x_reg_0;
endmodule


