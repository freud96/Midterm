/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:24:31 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__21,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__46;
wire [22:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82;
wire [0:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195;
wire [20:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197;
wire [32:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N677,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N679,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N683,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N684,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N700,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N702,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N703,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N709,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N711,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N713,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N718,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N720,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N724,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N729,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N731,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N732,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N737,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N738,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N743,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N750,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N755,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N758,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N759,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N761,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3946,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3968,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4006,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4009,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4018,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4029,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4070,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4088,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4095,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4109,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4118,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4127,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4154,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4157,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4167,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4170,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4211,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4219,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4236,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4247,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4249,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4252,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4257,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4258,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4260,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4261,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4264,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4266,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4271,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4279,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4282,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4284,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4338,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4351,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4382,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4384,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4395,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4397,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4420,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4457,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4468,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4488,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4506,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4524,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4614,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4618,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4621,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4649,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4653,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5461,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5558,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5583,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5951,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5964,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5968,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5981,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5991,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6003,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6006,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6009,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6013,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6020,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6036,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6053,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6061,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6069,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6088,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6094,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6095,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6125,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6140,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6153,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6154,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6159,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6164,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6189,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6219,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6240,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6248,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6251,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6252,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6256,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6258,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6264,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6265,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6266,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6267,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6269,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6274,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6279,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6282,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6357,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6361,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6362,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6382,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6395,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6401,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6412,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6420,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6461,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6475,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6477,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6488,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6506,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6517,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6558,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6570,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7319,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7328,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7354,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7375,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7395,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7457,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7488,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7517,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7524,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7572,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7620,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7633,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7661,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7663,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7665,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7666,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7667,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7669,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7670,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7674,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7676,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7679,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7684,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7702,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7709,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7713,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7715,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7716,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7720,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7731,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7738,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7759,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7761,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7764,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7765,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7766,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7768,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7769,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7773,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7775,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7776,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7777,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7780,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7781,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7782,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7785,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7787,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7788,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7791,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7792,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7795,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7798,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7800,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7801,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7804,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7805,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7806,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7807,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7808,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7812,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7813,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7814,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7816,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7819,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7822,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7825,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7826,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7828,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7835,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7841,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7843,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7849,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7851,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7855,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7857,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7860,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7861,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7866,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7867,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7875,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7902,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7916,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8583,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8589,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8603,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8618,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8620,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8621,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8642,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8651,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8653,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8656,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8659,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8661,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8662,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8663,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8665,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8666,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8667,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8668,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8670,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8671,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8672,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8673,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8674,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8675,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8676,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8679,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8703,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8713,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8714,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8715,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8716,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8731,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8732,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8740,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8743,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8750,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8758,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8765,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8766,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8768,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8769,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8770,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8771,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8773,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8774,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8775,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8777,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8778,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8780,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8782,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8783,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8785,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8787,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8788,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8789,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8790,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8791,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8793,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8796,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8797,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8798,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8800,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8802,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8803,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8804,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8806,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8808,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8809,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8810,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8812,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8813,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8814,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8816,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8818,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8820,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8822,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8823,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8825,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8826,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8831,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8834,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8835,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8839,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8841,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8846,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8849,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8851,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8855,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8857,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8858,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8860,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8862,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8866,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8868,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8870,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8873,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8875,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8898,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8916,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8930,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8943,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8946,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8972,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8981,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8982,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9003,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9006,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9013,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9060,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9094,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9109,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9140,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9143,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9157,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9159,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9164,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9180,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9189,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9196,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9236,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9240,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9247,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9248,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9257,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9258,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9259,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9263,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9264,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9265,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9266,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9267,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9269,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9273,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9274,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9357,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9361,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9362,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9389,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9397,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9401,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9461,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9468,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9475,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9517,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9524,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9570,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9572,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9589,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9593,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9614,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9620,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9621,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9633,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9642,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9653,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9659,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9661,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9662,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9663,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9665,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9666,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9667,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9668,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9670,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9674,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9676,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9683,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9702,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9709,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9715,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9720,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9724,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9743,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9755,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9759,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9761,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9764,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9766,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9768,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9770,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9771,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9772,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9774,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9779,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9780,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9781,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9784,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9786,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9787,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9788,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9790,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9791,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9792,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9793,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9794,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9797,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9798,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9800,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9801,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9805,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9806,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9807,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9809,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9810,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9812,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9813,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9814,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9815,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9818,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9819,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9821,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9824,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9825,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9831,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9841,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9842,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9848,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9849,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9851,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9855,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9856,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9857,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9862,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9870,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9871,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9873,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9898,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9930,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9946,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9956,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9964,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9968,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9981,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9991,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10003,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10009,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10018,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10020,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10029,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10053,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10060,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10061,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10088,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10094,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10118,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10140,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10143,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10153,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10164,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10170,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10180,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10211,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10233,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10236,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11846,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11866,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11916,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11930,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12061,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12196,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12219,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12259,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12269,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12327,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13477,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18828,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18861,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18874,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N37297;
wire N18241,N18245,N18402,N18406,N19158,N19431,N19751 
	,N19755,N20260,N20265,N20270,N20275,N20280,N20285,N20290 
	,N20295,N20355,N20370,N20382,N20609,N20613,N20621,N20625 
	,N20628,N20632,N20654,N20872,N20876,N20886,N20890,N20899 
	,N20903,N20912,N20916,N21060,N21064,N21306,N21310,N21559 
	,N21570,N21574,N21818,N21831,N21833,N21853,N21863,N21873 
	,N21883,N21893,N21903,N21913,N21923,N21933,N21943,N21953 
	,N21963,N21973,N21983,N21993,N21997,N22003,N22005,N22007 
	,N22034,N22040,N22048,N22056,N22064,N22066,N22072,N22080 
	,N22082,N22091,N22097,N22101,N22105,N22109,N22113,N22117 
	,N22121,N22123,N22125,N22129,N22131,N22133,N22137,N22139 
	,N22141,N22145,N22147,N22149,N22153,N22155,N22157,N22194 
	,N22199,N22201,N22203,N22205,N22209,N22211,N22213,N22217 
	,N22219,N22221,N22225,N22227,N22229,N22233,N22235,N22237 
	,N22241,N22243,N22245,N22249,N22251,N22253,N22258,N22260 
	,N22268,N22270,N22278,N22286,N22288,N22290,N22294,N22296 
	,N22306,N22310,N22314,N22316,N22318,N22322,N22324,N22326 
	,N22678,N22680,N22961,N22962,N22963,N22964,N22965,N22966 
	,N22968,N22969,N22971;
EDFFHQX1 x_reg_22__retimed_I12950 (.Q(N22680), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12949 (.Q(N22678), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12809 (.Q(N22326), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9253), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12808 (.Q(N22324), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10035), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12807 (.Q(N22322), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10214), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12806 (.Q(N22318), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8673), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12805 (.Q(N22316), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10176), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12804 (.Q(N22314), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9633), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12803 (.Q(N22310), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9017), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12801 (.Q(N22306), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9999), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12798 (.Q(N22296), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12797 (.Q(N22294), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12796 (.Q(N22290), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9642), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12795 (.Q(N22288), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8873), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12794 (.Q(N22286), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9829), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12792 (.Q(N22278), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12790 (.Q(N22270), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10005), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12789 (.Q(N22268), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9052), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12787 (.Q(N22260), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9402), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12786 (.Q(N22258), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9205), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12785 (.Q(N22253), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9143), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12784 (.Q(N22251), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9720), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12783 (.Q(N22249), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10117), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12782 (.Q(N22245), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9597), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12781 (.Q(N22243), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10140), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12780 (.Q(N22241), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8835), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12779 (.Q(N22237), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9098), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12778 (.Q(N22235), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10073), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12777 (.Q(N22233), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8592), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12776 (.Q(N22229), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9559), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12775 (.Q(N22227), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9130), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12774 (.Q(N22225), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8800), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12773 (.Q(N22221), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9257), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12772 (.Q(N22219), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9827), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12771 (.Q(N22217), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10217), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12770 (.Q(N22213), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8588), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12769 (.Q(N22211), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9862), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12768 (.Q(N22209), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9521), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12767 (.Q(N22205), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12391), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12766 (.Q(N22203), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12765 (.Q(N22201), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12764 (.Q(N22199), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12134), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12762 (.Q(N22194), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11893), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12748 (.Q(N22157), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8629), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12747 (.Q(N22155), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9320), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12746 (.Q(N22153), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9578), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12745 (.Q(N22149), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8845), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12744 (.Q(N22147), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10061), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12743 (.Q(N22145), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9627), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12742 (.Q(N22141), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8967), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12741 (.Q(N22139), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10185), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12740 (.Q(N22137), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9946), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12739 (.Q(N22133), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8942), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12738 (.Q(N22131), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9681), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12737 (.Q(N22129), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9919), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12736 (.Q(N22125), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9532), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12735 (.Q(N22123), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9942), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12734 (.Q(N22121), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8777), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12733 (.Q(N22117), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9688), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12731 (.Q(N22113), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8918), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12730 (.Q(N22109), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9289), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12728 (.Q(N22105), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8587), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12727 (.Q(N22101), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9571), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12725 (.Q(N22097), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8813), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12723 (.Q(N22091), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12028), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12719 (.Q(N22082), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9909), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12718 (.Q(N22080), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8745), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12715 (.Q(N22072), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8846), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12713 (.Q(N22066), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10049), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12712 (.Q(N22064), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9296), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12709 (.Q(N22056), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9169), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12706 (.Q(N22048), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9899), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12703 (.Q(N22040), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8877), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12701 (.Q(N22034), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12690 (.Q(N22007), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[34]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12689 (.Q(N22005), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[34]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12688 (.Q(N22003), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12687 (.Q(N21997), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[33]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12685 (.Q(N21993), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12682 (.Q(N21983), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12679 (.Q(N21973), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12676 (.Q(N21963), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12673 (.Q(N21953), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12670 (.Q(N21943), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12667 (.Q(N21933), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12664 (.Q(N21923), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12661 (.Q(N21913), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12658 (.Q(N21903), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12655 (.Q(N21893), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12652 (.Q(N21883), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12649 (.Q(N21873), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12646 (.Q(N21863), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12643 (.Q(N21853), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12636 (.Q(N21833), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12635 (.Q(N21831), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12632 (.Q(N21818), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12171), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12562 (.Q(N21574), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12560 (.Q(N21570), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12557 (.Q(N21559), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12327), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12474 (.Q(N21310), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12472 (.Q(N21306), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12391 (.Q(N21064), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12389 (.Q(N21060), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12340 (.Q(N20916), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12338 (.Q(N20912), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12335 (.Q(N20903), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12333 (.Q(N20899), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12330 (.Q(N20890), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12328 (.Q(N20886), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12325 (.Q(N20876), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12323 (.Q(N20872), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12241 (.Q(N20654), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12004), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12232 (.Q(N20632), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12086), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12230 (.Q(N20628), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12222), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12229 (.Q(N20625), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12444), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12227 (.Q(N20621), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11950), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12224 (.Q(N20613), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12168), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12222 (.Q(N20609), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12306), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12129 (.Q(N20382), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12309), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12124 (.Q(N20370), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11895), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12118 (.Q(N20355), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12089), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12103 (.Q(N20295), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11872), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12101 (.Q(N20290), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11829), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12099 (.Q(N20285), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12040), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12097 (.Q(N20280), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12063), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12095 (.Q(N20275), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12259), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12093 (.Q(N20270), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12285), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12091 (.Q(N20265), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12234), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12089 (.Q(N20260), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11852), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I11924 (.Q(N19755), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12367), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I11922 (.Q(N19751), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11869), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I11834 (.Q(N19431), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I11739 (.Q(N19158), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_26__retimed_I11459 (.Q(N18406), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_26__retimed_I11457 (.Q(N18402), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I11390 (.Q(N18245), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I11388 (.Q(N18241), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I13091 (.Y(N22961), .A(N18241));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13096 (.Y(N22966), .A(N22961));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13095 (.Y(N22965), .A(N22961));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13094 (.Y(N22964), .A(N22961));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13093 (.Y(N22963), .A(N22961));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13092 (.Y(N22962), .A(N22961));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_3_I0 (.Y(bdw_enable), .A(astall));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13161), .A(a_exp[7]), .B(a_exp[0]));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13163), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18854), .A(a_exp[6]), .B(a_exp[5]), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13163));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I4 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13161), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18854));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I5 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18861), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I6 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18861));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I7 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13197), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I8 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13201), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13197));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I9 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13184), .A(a_man[10]), .B(a_man[9]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I10 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13203), .A(a_man[6]), .B(a_man[5]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I11 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13192), .A(a_man[8]), .B(a_man[7]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I12 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13212), .A(a_man[4]), .B(a_man[3]));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13195), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13203), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13192), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13212));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I14 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13206), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I15 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13216), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I16 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__24), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13201), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13195), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13206), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13216));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I17 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__24));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I18 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I19 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13110), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I20 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13114), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I21 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__17), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13110), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13114));
AOI211XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I22 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13141), .A0(a_exp[2]), .A1(a_exp[1]), .B0(a_exp[3]), .C0(a_exp[4]));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I23 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13138), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13141), .B(a_exp[5]), .C(a_exp[6]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I24 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__21), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13138), .B(a_exp[7]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I25 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385), .A(a_exp[3]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I26 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364), .A(a_exp[1]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I27 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364), .B(a_exp[2]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I28 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I29 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371), .A(a_exp[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I30 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379), .A(a_exp[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I31 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376), .A(a_exp[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I32 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376), .B(a_exp[7]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I33 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379), .B(a_exp[6]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I34 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18845), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[6]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I35 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[8]), .AN(a_exp[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I36 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__46), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18845), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[8]));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I37 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__17), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__21), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__46));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I38 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I39 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13910), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I40 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13910));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I41 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[29]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I42 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .A(a_man[21]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I43 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270), .A(a_man[22]), .B(a_man[20]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I44 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I45 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957), .A(a_man[21]), .B(a_man[19]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I46 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I47 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4204), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4042), .A(a_man[19]), .B(a_man[22]), .CI(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I48 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361), .A(a_man[18]), .B(a_man[20]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4204));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I49 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I50 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4545), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4391), .A(a_man[16]), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I51 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622), .A(a_man[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4545), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4042));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I52 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I53 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I54 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4506), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .B(a_man[19]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I55 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4229), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4185), .A(a_man[15]), .B(a_man[17]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4506));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I56 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198), .A(a_man[22]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I57 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4170), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198), .B(a_man[20]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I58 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4229), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4170), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4391));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I59 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I60 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198), .B(a_man[20]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I61 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .A(a_man[20]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I62 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .B(a_man[18]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I63 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4571), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4081), .A(a_man[14]), .B(a_man[16]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4130));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I64 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4571), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4185));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I65 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I66 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I67 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I68 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .B(a_man[19]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I69 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975), .A(a_man[19]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I70 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4466), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975), .B(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I71 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4193), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3976), .A(a_man[13]), .B(a_man[15]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4466));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I72 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4348), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4193), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4081));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I73 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I74 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .B(a_man[18]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I75 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385), .A(a_man[18]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I76 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4404), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4246), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385), .B(a_man[16]), .CI(a_man[13]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I77 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4533), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4594), .A(a_man[12]), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4404));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I78 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4533), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3976));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I79 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I80 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I81 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975), .B(a_man[17]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I82 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069), .A(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I83 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4336), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4183), .A(a_man[10]), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I84 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4029), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4588), .A(a_man[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I85 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4158), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4488), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4336), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4029));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I86 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4311), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4158), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4594));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I87 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I88 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471), .A(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I89 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3960), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4126), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I90 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4092), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4617), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3960), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4588), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4183));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I91 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4246), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4092), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4488));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I92 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I93 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I94 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I95 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4435), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I96 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565), .A(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I97 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4577), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4420), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975), .B(a_man[21]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I98 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162), .A(a_man[15]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I99 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I100 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4455), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4359), .A(a_man[13]), .B(a_man[22]), .CI(a_man[10]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I101 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4300), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4577), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4232), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4359));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I102 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4428), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4006), .A(a_man[9]), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4300));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4395), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I104 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4521), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4365), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4455), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4126));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I105 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4428), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4521), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4617));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I107 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4324), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4377), .A(a_man[9]), .B(a_man[12]), .CI(a_man[7]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I108 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4314), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4161), .A(a_man[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I109 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4510), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4625), .A(a_man[6]), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4314));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I110 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4173), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4018), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4420), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4510), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4377));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I111 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4207), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4241), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4324), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4173));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I112 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4207), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4006));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253), .A(a_man[13]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I116 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4043), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I117 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4444), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4288), .A(a_man[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I118 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4186), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4031), .A(a_man[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I119 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4383), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4135), .A(a_man[5]), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4186));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I120 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4351), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4197), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4383), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4625));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I121 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4078), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4260), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4444), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4351));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I122 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4078), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4241));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939), .A(a_man[12]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I125 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4640), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I126 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4058), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4630), .A(a_man[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I127 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4252), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4368), .A(a_man[4]), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4058));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I128 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4221), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4470), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4252), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4135));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I129 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4264), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4495), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4640), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4288), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4221));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I130 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4018), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4264), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4260));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339), .A(a_man[11]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I135 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4500), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471), .B(a_man[9]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I136 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4120), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4613), .A(a_man[3]), .B(a_man[5]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4630));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I137 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4093), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4338), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4120), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4368));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I138 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4137), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4500), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4161), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4093));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I139 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4197), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4137), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4495));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032), .A(a_man[10]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I142 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4369), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4210), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I143 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4236), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4237), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385), .B(a_man[16]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I144 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3963), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4524), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4236), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4210), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4613));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I145 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4002), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4249), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4031), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3963));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I146 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4067), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4002), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4016));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I149 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4023), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4474), .A(a_man[3]), .B(a_man[6]), .CI(a_man[1]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121), .A(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I151 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4266), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4601), .A(a_man[15]), .B(a_man[22]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I152 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4082), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4653), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4023), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4266), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4237));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I153 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432), .A(a_man[9]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I154 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3987), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4123), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432), .B(a_man[7]), .CI(a_man[4]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4200), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I156 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4549), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4397), .A(a_man[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4200), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4123));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I157 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4591), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4485), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4082), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3987), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4549));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I158 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3936), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4591), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4249));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525), .A(a_man[7]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I161 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4386), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4012), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I163 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4107), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3952), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4386), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4046), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4601));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I164 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4641), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4473), .A(a_man[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I165 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4138), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4621), .A(a_man[2]), .B(a_man[5]), .CI(a_man[0]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I166 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4581), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4421), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4641), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4138), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4474));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I167 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4457), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4004), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4107), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4581), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4653));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I168 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4524), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4485));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I169 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097), .A(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I173 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4096), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3940), .A(a_man[4]), .B(a_man[13]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I174 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4187), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I175 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4224), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4096), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4187), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4012));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I176 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3977), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4541), .A(a_man[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4473), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4621));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I177 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4486), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4224), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3977), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4421));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I178 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4397), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4486), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4004));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631), .A(a_man[5]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I181 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4372), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4211), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I182 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4566), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4247), .A(a_man[19]), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4372));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I183 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4614), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4541), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4566), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4070));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I184 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3952), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4614), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4355));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I187 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4655), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4175), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I188 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4124), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4511), .A(a_man[0]), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4655));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I189 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4409), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4033), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4124), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4247));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I190 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4458), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I191 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3965), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4211), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4306), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4511));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I192 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4317), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4458), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3965));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I193 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4409), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4317), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4493));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I195 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445), .A(a_man[3]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I196 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3955), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4516), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I197 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4049), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I198 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4489), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3955), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4049), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4175));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304), .A(a_man[4]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I200 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4400), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4056), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I201 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4238), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4086), .A(a_man[17]), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4056));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I202 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4597), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4489), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4400), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4238));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I203 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4597), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4255), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4132));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I206 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I207 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4227), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975), .B(a_man[9]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I208 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4423), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4410), .A(a_man[16]), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4227));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I209 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4151), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3937), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4331), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4423), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4086));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I210 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4151), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4527), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4394));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I211 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398), .A(a_man[2]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4505), .A(a_man[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I214 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3980), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4505));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I215 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4268), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4110), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3980), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4410));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I216 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4320), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4166), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I217 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4543), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4388), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4166), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3953));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I218 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4179), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4516), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4320), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4543));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I219 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4268), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4179), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3937));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I221 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I222 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4284), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4574), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I223 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4214), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I224 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4333), .A(a_man[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I225 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4346), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4191), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4284), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4214), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4333));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I226 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4258), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .A(a_man[1]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I228 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4100), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4215));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I229 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4449), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4346), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4258), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4100));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I230 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4449), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4110), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4293));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I232 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4403), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4244), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121), .B(a_man[13]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I233 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4156), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I234 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4129), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4403), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4156), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4574));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I235 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4009), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4129), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4191));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I236 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4388), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4009), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4550));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966), .A(a_man[0]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I242 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4335), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162), .B(a_man[5]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I243 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3993), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4335), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4116), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4244));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I244 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4037), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3993));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I245 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3944), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4037), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4101));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I247 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4586), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I248 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4519), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069), .B(a_man[4]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I249 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4182), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4027), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4519), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4427), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4353));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I250 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4636), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4000), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4586), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4182));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I251 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3969), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4454));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I254 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4052), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4624), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I255 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3984), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4109), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I256 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4364), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3984), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4624), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4592));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I257 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4090), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4364));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I258 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4556), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4090), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4000));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I260 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4230), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4076), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I261 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4172), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I262 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4546), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4393), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4172), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4076), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4109));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I263 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4271), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4230), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4546));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I264 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4271), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4235));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I266 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4638));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4178), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4104), .A(a_man[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3948), .A(a_man[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I270 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4649), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4225), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3948));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I271 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4453), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3988), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4649));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I272 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4453), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4206), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4472));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I274 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4507), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4242), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I275 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4041), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4360), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I276 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4014), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4041), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4343));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I277 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4014), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4393), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3988));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I278 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4001), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4602), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4001));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I280 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4219), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4066), .A(a_man[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I281 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4536), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4382), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I282 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4608), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4219), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4536), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4360));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I283 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4480), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4573), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4608), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4225));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4480));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4145));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4498), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I288 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4639), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4604), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4498));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I289 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4160), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3999), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I290 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4287), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4066), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4160));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I291 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4382), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4639), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4478));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I292 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4442), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4287), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4242));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I293 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I294 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4529), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I295 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4560), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I296 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4560), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3999), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4604));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I298 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4184), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253), .B(a_man[4]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4337), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I300 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4337), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3995));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4567), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I302 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3962), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I303 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4429), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4015), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I304 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4015));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I305 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4429), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4626));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I308 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4456), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4367), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I309 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4208), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4250), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I310 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4456), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4250));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I311 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4208), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4136));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I312 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4576), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I314 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4396), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I315 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4396), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4367));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I317 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4484), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I318 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4234));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I320 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4325));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I321 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4530), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I322 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445), .CI(a_man[6]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I323 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I324 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I325 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I326 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3978), .A(a_man[1]), .B(a_man[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I333 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4088), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I334 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4243), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4047), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4088), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4243));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4329), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4201), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3978), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4047));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4154), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I339 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4514), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4554), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4154));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4595), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3992), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4329), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4514));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I341 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4222), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4634), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4595), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4580), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4213), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4222), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4062));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4118), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4530), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4580), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3968), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4282), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4563), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3968), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4282));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4508), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4127), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4118), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4563));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4283), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4576), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4508));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I350 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I351 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I352 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4418), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4599), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4190));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I353 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4098), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4323), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4503), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4098));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4600), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4418), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4323));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4347), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4283), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4600));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I359 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3961), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4413), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4007));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4460), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4567), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4347), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3961));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I363 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I364 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4373), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4318), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4643));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I365 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3935), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4529), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4460), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4373));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I366 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4128), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18828), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3935), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I367 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4559), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I368 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4439), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4559), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I369 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4602), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4128), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4439));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I370 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4468), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4468), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4345), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I374 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4025), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4345));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13097 (.Y(N22968), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4025));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13098 (.Y(N22971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13099 (.Y(N22969), .A(N22968), .B(N22971));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I13100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059), .A(N22969));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I377 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I378 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I379 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4257), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4257));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I381 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I382 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I383 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I384 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4167), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I385 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4654), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4167));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I386 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4371), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4654));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I387 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4526), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4371));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I388 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I389 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I390 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4072), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I392 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4072));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3979), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4551), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3979));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I398 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4341), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4551));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I399 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4341));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I400 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4619), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I404 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4619));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I406 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I407 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4515), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4459), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4515));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4279), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4459));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4435), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4279));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270));
OAI2BB2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4499), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I414 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4499));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169), .A(a_man[22]), .B(a_man[21]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4102), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I420 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4261), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3946), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4102));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I421 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4261), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I422 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649), .S0(a_exp[0]));
OA22X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938), .B0(a_man[22]), .B1(a_man[21]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651), .S0(a_exp[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N37297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[1]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I428 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N37297));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I429 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4223), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4387), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4223), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4387));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I434 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4119), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4275));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I437 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4217), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I438 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4380), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4532), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4217), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4380));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I442 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645), .S0(a_exp[0]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I445 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4607), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I446 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4038), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4440), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4607));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4038), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I450 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[1]), .B(a_exp[2]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371), .B(a_exp[5]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5483), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372), .B(a_exp[4]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650), .S0(a_exp[0]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652), .B(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5578), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5578), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N706), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4629), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4629), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4057));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4310), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3998), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4157));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I482 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I483 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I486 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I487 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5606), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_3_I489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N704));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_3_I490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I493 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4091), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4497), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3933));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5513), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I503 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N702), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I504 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N702), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I514 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5465), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5465), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I519 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N701), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I520 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5558), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5558), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_3_I528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N703));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I529 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5436), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I535 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N705));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6280), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6280));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6209), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_3_I541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I542 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I543 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I544 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6125), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6209), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I547 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6355));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[28]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6125), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5921), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178), .A(1'B0), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I554 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I555 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6057), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I557 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6478), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I558 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5965), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6057), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6478), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6254), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I562 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6254));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I563 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[27]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5965), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6172), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I564 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399), .A(1'B1), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[27]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6003), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5890), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6003), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I570 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I571 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6332), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I572 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6519), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5890), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6332), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I573 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6103), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6251), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I576 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6022), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6103), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6251), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[26]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6519), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6022), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I578 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122), .A(1'B1), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[26]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I581 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979));
AOI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6446), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I588 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I589 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6066), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6175), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6066), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I592 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6369), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6446), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6175), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I595 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5940), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5952), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5952));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6564), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5940), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5936), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[25]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6369), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6564), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I600 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853), .A(1'B1), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[25]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I603 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I604 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4587), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I605 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4587), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I610 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5586), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I611 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5586), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I612 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5580), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I613 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N699), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I614 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3959), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3959), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5539), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5485), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I623 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5485), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I624 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N698), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I625 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5417), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5417), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I630 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N700), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8912), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8912));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I635 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9401), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9401), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I638 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N763), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6042), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N763));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I642 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[42]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I643 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I644 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I645 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6299), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I646 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I647 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6024), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6217), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6299), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6024), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6493), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I653 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I654 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6507), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I655 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I656 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6488), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6507), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6412), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6493), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6488), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[24]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6217), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6412), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I659 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[24]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I663 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6144), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I664 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6567), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6067), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6144), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6567), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6189), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6341), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6265), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6189), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6341), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[23]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6067), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6265), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[41]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[42]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5490), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I679 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5608), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5490), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5604), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5604), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4054), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I687 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5515), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5444), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5616), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5509), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5616), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N696), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5515), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5509), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8946), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8946));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9435), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I703 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5970), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6431), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6491), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6566), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6431), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6491), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N762), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5970), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6566), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I710 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N762));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9092), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I713 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[41]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[40]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9092));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I714 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[23]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[41]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[41]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6539), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I717 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I719 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6415), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I720 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5897), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6539), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6415), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I721 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6494), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6185), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6134), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6110), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6580), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6185), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[22]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5897), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6110), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I729 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6523), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6285), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I732 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6342), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6414), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6285), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6342), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N761), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6523), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6414), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N761));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I738 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8732), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9236), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I744 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I745 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I746 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5613), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5613), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5523), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N695), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5419), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5414), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N695), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4146), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4146), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I755 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I757 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5566), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5537), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5428), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5537), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8982), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I765 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8982));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I766 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I767 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I768 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6178), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I769 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6376), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6178), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I770 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I771 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6131), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I772 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I773 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6188), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6267), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6131), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6188), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N760), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6376), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6267), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I777 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N760));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I778 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I779 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10066), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I780 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9847), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9128), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10066));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I781 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[40]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[39]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8732), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9236), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9847));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I782 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[40]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[22]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[40]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I783 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I786 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144), .A(N22678), .B(N22680));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I787 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6088), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I789 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I790 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6268), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I791 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6453), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6088), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6268), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I794 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6427), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I795 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I796 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6036), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5948), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6427), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6036), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[21]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6453), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5948), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9468), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I800 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I801 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I802 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I803 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I804 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I805 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I806 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I807 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5520), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I810 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I811 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5550), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5447), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5440), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N693), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4650), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4582), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I816 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4095), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I817 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I818 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4095), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4254));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I819 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4582), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4022));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I822 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4231), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4650), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4079));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I823 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4231), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I827 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5472), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9013), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I834 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9013));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8766), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I838 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9302), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9555), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8766));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10100), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I841 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I842 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9166), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I843 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9163), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I844 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8986), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10100), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9166), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9163));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I845 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6090), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I846 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I847 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6028), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I848 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6223), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6090), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6028), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I849 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I850 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5971), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I851 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6168), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6038), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6168), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6112), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5971), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6038), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I855 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N759), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6223), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6112), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I858 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I859 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10055), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9691), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8986), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9707), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8924));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I860 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[39]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[38]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9302), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10055));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I861 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[39]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[21]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[39]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I862 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I863 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5920), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I864 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I865 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6113), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6308), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5920), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6113), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I870 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6282), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I871 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I872 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6577), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I873 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6502), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6282), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6577), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I874 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[20]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6308), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6502), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I875 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9497), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I879 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I881 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I882 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I883 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5461), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I884 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5424), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5461), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5476), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5424), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N691), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5476), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N691), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4579), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4017), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4419), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4579));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I892 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4017), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I893 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I894 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5413), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5599), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I899 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N690), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I900 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9050), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I901 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9050));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I902 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I903 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6212), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I904 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5922), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6212), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6207), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6571), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6207), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6072), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5922), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6571), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I908 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6525), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I910 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6579), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I912 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5950), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6525), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6579), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I913 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N758), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6072), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5950), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I914 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N758));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I915 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6061), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I916 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6475), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6061), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I917 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I918 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I919 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6417), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I920 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5903), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6475), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6417), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I921 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6426), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6505), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6074), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6426), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N757), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5903), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6505), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I927 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N757));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I928 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I929 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I930 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8699), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8940));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I931 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I932 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9321), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I933 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8774), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10114), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8699), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9321), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8648));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I934 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I935 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9742), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I936 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I937 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8797), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I938 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I939 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6329), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6270), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6456), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6329), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6270), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5904), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I947 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6279), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I949 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6360), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5904), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6279), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N756), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6456), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6360), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I951 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N756));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I952 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I953 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I955 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9200), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I956 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9228), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I957 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8624), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9200), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9228));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I958 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9438), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9742), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8797), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8624));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I959 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I960 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I962 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10135), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I963 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9528), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I965 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I966 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I967 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I968 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I969 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I970 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I971 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5583), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5583), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5505), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5547), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5505), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I975 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I976 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I977 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4509), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4509), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5535), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5501), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5535), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I983 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5501), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I984 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I985 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N688), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I986 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9086), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I987 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9086));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I989 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I990 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I991 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10210), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8974));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I992 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10088), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9358), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10135), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10210));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I993 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10178), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9818), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10088), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10032), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9045));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I994 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9529), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9140), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10114), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9438), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10178));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I995 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[38]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[37]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9691), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8774), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9529));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I996 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[38]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[20]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[38]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I997 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I998 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I999 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1000 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6474), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1002 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5951), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6153), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6474), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5951), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1005 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6126), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1006 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6424), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6356), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6126), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6424), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[19]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6153), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6356), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8834), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1013 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6173), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1014 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1015 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6116), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6312), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6173), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6116), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1017 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1018 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1019 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6458), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1020 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6124), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1021 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6202), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6458), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6124), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1022 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N755), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6312), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6202), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1023 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N755));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1025 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9920), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1027 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1028 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9247), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8870), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8834), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9920), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9781));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1029 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9109), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8751), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9247), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9724));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1030 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1031 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9956), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1033 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6023), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6304), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5955), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6159), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6023), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5955), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1038 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6182), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6314), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6182), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5964), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1044 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6049), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6314), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5964), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1045 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N754), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6159), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6049), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1046 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N754));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1047 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1048 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6565), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1049 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1050 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6509), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1051 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6000), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6565), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6509), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6160), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1055 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6518), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1058 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5882), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6160), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6518), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N753), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6000), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5882), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N753));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1061 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1062 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9158), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1063 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8866), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1065 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9510), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9158), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8866));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1066 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1067 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1069 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5403), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1074 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5487), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5403), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1075 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5452), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5487), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1076 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5532), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5452), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1077 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1078 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N687), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1079 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1080 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4611), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1081 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1082 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1083 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5571), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1084 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5571), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1085 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5404), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5441), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1086 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5435), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5404), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1087 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1088 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N686), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9124), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9124));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1091 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1092 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1093 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1094 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8758), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10094), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9668), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9005));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1095 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1096 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9546), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9242), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9294), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1100 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8656), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9546), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9242), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9294));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1101 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9149), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8782), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9510), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8758), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10173), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1105 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1107 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1108 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10123), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10173), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8638), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9392));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1109 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10002), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8656), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9854));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1110 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9019), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8674), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9149), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8870), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9637));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1111 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9883), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9502), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9019), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10002), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8751));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1112 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9208), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8839), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9109), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9883));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7459), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1118 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7328), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1120 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1121 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7459), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7328), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7293));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1122 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7316), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1128 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7375), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7709), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1130 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7896), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7751), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7375), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7709));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1131 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7316), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7344), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7896));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1135 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7887), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1136 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1137 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1138 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7616), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7473), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7887), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7682));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1139 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7753), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1140 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7616), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7753), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7751));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1142 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7543), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1144 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7787), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7608), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1146 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7872), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7731), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7543), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7787), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7608));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7837), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1149 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7300), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7455), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1152 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7592), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7452), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7300), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7322), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7455));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1153 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7330), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7835), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7734), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7837), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7592));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1154 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7471), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7872), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7330));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1158 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7926), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1162 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7676), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7535), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7909), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7926), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7687));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7395), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1165 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7665), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7878), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1168 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7308), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7814), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7665), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7878));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1169 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7697), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7676), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7395), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7308));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1170 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7731), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7835));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1173 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7379), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1175 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7754), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7620), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7379), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7538));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1176 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7411), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7535), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7754), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7814));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1177 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7556), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7452), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7411));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1178 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7761), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1183 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7765), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1187 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7337), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7765), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7745));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1188 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7388), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7900), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7761), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7599), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7337));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7314), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1192 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7838), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7903), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7893), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7314));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1193 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7613), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7465), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1195 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1196 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7702), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7613), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7465), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7924));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1197 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7545), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1198 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7476), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7702), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7545), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7841));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1199 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7775), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7620), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7838), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7476));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1200 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7925), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7388), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7775));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1206 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7927), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7777), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7680), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7483));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1207 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1208 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1209 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1210 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7417), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7931), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7639), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7325), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7394));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1211 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7341), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7336), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1215 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7780), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7341), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7336), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7828));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1216 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7557), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7417), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7780), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7560));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1217 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7499), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7699), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7927), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7557));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1218 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7499), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7900), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7640));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1219 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1221 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7365), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1224 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1225 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7354), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1226 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7826), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1228 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7865), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7726), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7354), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7694), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7826));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1229 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7356), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7861), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7628), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7865));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1230 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7342), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7759), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1232 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7730), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1233 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7503), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7359), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7759), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7730));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1234 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7641), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7500), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7643), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7503), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7931));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1235 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7859), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7777), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7356), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7641));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1236 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7333), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7355));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5486), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5526), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5610), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5573), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5556), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[1]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1247 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7918), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1249 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1250 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7667), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7706), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7918), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7407));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1251 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7843), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1254 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7480), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1256 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7301), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7806), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7720), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7480));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1257 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7440), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7667), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7843), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7301));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1258 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1261 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7586), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7451), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7707), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7358));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1262 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7723), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7582), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7586), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7359));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1263 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7581), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7438), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7861), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7440), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7723));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1264 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7581), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7414), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7722));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1266 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7437), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4384), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4615), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1272 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4045), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4446), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4615));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4537), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1274 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3973), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4384), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4045), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4537));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1275 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N623), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1276 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5438), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N623), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1277 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5438), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1278 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5478), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5463), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5528), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N684), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1283 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7565), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1284 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7746), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7611), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7915), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7437), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7565));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7830), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7813), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7421), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7725), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1291 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7380), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7813), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7421), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7725));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1292 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7524), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7378), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7830), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7380));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1293 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7804), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7663), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7806), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7526), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7444));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1294 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7296), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7297), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7524), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7804));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1295 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7296), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7500), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7438));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1300 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7552), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7534));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1302 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7520), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1303 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1304 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7635), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7520), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7494));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1305 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7609), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7552), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7635));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7631), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7800), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1309 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7920), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7769), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7631), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7800), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7625));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1310 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7888), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7744), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7920), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7891));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1311 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7661), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7609), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7888));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1312 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7661), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7582), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7801));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1318 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7349), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7852), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7882), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7507));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1320 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1321 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7339), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1322 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7346), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1323 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7716), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7574), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7522), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7339), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7346));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1324 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7688), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7442), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7716));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1325 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7323), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7492), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7405), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7769));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1326 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7377), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7886), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7688), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7323));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1327 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7377), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7663), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7523));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7604), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7885), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1332 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7795), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7657), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7604), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7576), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7885));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1333 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7402), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7916), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7852), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7795), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7574));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1334 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7805), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1338 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7431), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7705));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1339 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7766), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7633), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7805), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7899), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7431));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1340 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7742), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7607), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7402), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7766), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7550));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1341 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7742), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7744), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7886));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7619), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7869), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1347 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7849), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7619), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7869), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7525));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1350 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7517), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7419), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7606));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1351 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7488), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7347), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7517), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7657));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1352 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7463), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7321), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7633), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7849), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7488));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1353 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7827), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7607));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7320), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1357 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7880), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7684), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7320));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7889), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1359 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7572), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7880), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7889), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7372));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7332), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1363 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7286), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7319), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7426), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7332));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1364 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7825), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7286), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7713));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1365 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7916), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7825), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7321));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1366 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1367 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1368 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1369 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1370 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7791), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7782), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1374 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7370), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7791), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7306), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7782));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1375 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1377 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7655), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7514), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7610), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7698), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7739));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1378 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7547), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7792), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7370), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7655));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1379 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7347), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7547), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7686));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1381 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1382 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7505), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1383 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7398), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1384 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7457), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7312), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7513), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7505), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7398));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1385 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1386 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1387 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7736), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7597), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7413), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7324));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1388 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7914), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7764), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7736), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7877));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1389 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7428), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7400));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1390 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1392 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1395 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7540), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7399), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1398 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7819), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7776));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1399 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7630), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7486), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7540), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7819), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7597));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1400 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7514), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7630), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7764));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7588), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7596), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1404 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7906), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7588), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7596));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1406 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7345), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7906), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7690), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7679));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1407 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7345), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7312), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7486));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7860), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7768), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1414 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7424), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7938), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7860), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7304), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7768));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7404), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7845), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1419 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7623), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7845), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7311));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1420 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7710), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7404), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7484), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7623));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1421 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7424), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7757), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7569));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1422 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7392), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7710), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7847));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7632), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7670), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1427 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7788), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7650), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7670), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7568));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1428 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7788), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7938));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1429 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7935), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7391), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1432 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7509), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7366), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7935), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7391));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7490), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1434 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7509), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7490), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7650));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7851), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1437 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7383), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1438 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7851), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7383), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7366));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7866), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1442 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7749), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7648));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7587), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7364), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1445 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7469), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1446 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7364), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7469));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1450 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7482), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7600), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7669), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7482), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7430), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7303), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7600), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7808));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7829), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7587), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7430), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7585), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7866), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7829), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7727));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7905), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7504), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7585), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7571), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7781), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7905), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7645));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7563), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7487), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7933), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7563));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7632), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7571), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7487));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1482 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1483 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1486 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1487 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1493 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7807), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7551), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7807));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7939), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7551));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7674), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7939));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1503 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7409), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7812), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7674));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1504 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7443), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[32]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7409), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7443));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1514 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1519 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1520 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1529 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1535 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7528), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7917), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7528));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7652), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7917));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7387), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7652));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7773), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7533), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7387));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7666), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1542 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7773), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7666));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1543 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10143), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9397), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[32]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1544 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10143));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9397));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10121), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1547 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[37]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[36]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9140), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10121));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1548 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[37]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[19]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[37]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6187), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6326), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6187), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6506), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1554 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5995), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6326), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6506), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1555 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6264), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1557 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5967), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6264), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1558 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6277), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6199), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5967), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6277), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[18]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5995), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6199), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1562 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1563 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[19]), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6115), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1564 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[19]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9620), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9588), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1570 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9362), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1571 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9091), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8731), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9588), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9276), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9362));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1572 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1573 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9813), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1576 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1578 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1580 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8875), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8668), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9432));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1581 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8579), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9889), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9813), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8875));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9596), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9596), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9702), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1588 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1589 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9455), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9063), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9702), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9040));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6413), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1592 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5986), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6363), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5986), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6550), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6413), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6363), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1595 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6274), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6002), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6274), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6368), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6438), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6002), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6368), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1600 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N752), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6550), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6438), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N752));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1603 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1604 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1605 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9988), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9195), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8901), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1610 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10192), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9832), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9988), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9195), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8901));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1611 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9644), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9455), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8789), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10192));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1612 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9283), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10094), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9644));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1613 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9912), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9539), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8579), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9763), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9283));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1614 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6266), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6205), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6398), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6266), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6205), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6120), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6552), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6120), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6370), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6216), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6370), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1623 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6291), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6552), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6216), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1624 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N751), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6398), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6291), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1625 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N751));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9851), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051));
NAND2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1630 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[1]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1635 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1638 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9269), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9350));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9315), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1642 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10018), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9654), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9841), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9315), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1643 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9223), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8849), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10128), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9851), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10018));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1644 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8678), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8731), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9223), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10216));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1645 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10038), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9674), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9889), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8678), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8907));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1646 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8934), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8601), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8782), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10038));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1647 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9790), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8674), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9912), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8934));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6020), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6020), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5975), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5975));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1653 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[18]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5981), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1654 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[18]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1655 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8855), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1656 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8897), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10233), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9790), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9502), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8855));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1657 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[36]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[35]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9620), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8839), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8897));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1658 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[36]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[36]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1663 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1664 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7634), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7368), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7634));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7752), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7368));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7496), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7897), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7752));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7890), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1679 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7496), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7890));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7617), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1687 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7348), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7733), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7348));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7472), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7733));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7855), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7617), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7472));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7466), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7855), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7466));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9524), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9524), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6495), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6536), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6495), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[17]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6536), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[17]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1703 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9837), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6111), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6054), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6248), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6111), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6054), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1710 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6399), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6065), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1714 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6137), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6399), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6065), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N750), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6248), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6137), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N750));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1717 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9772), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1719 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1720 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8826), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1721 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8825), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10163), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9470), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9772), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8826));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9621), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10237), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1728 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9805), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9621), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10237));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1729 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9979), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9615), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8825), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9805), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9063));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1732 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9459), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5949), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5885), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6472), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6096), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5949), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5885), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1738 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6513), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6098), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6513), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6377), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5896), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6377), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5979), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6098), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5896), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1744 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N749), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6096), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5979), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1745 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N749));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1746 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1748 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9623), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9230), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9459), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9386));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10027), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9231), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8937), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1755 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8667), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9987), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9231), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8937));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1756 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9587), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9194), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9623), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9654), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8667));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1757 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9002), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8661), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9587), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9832), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8849));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1758 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9415), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9027), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9255), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9979), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9002));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10164), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9884), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9661), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1765 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1766 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8723), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1767 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8694), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9661), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9269), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8723));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1768 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9391), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10164), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9884), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8694));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1769 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8640), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9955), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9391), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9425), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10163));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1770 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9771), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9385), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8640), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9615), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8661));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1771 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10158), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9797), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9771), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10008), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9027));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1772 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9056), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9674), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9415), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10158));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1773 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6316), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6345), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6385), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6316), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6345), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6053), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1777 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6123), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6053));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1778 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[16]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6385), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6123), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1779 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[16]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1780 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9066), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1781 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9699), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8601), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9066));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1782 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8810), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9407), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9699));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1783 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[35]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[34]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10233), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8810));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1786 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6171), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1787 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6361), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6547), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6171), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6361), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1789 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1790 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6520), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1791 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6461), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6122), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6461), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6046), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6520), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6122), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1794 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[17]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6547), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6046), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1795 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12171), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[35]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[17]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[35]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1796 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838), .A(N21831), .B(N21833));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6017), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5957), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1800 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1801 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6479), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1802 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6203), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6479), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1803 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6395), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6017), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6203), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1804 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6371), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1805 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1806 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5961), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1807 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5879), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6371), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5961), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[16]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6395), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5879), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10180), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1810 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10180));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1811 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9996), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1816 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6161), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1817 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6192), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1818 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6232), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6161), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6192), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1819 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5884), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5963), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5884), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[15]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6232), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5963), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1822 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[15]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1823 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10047), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9806), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1827 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8603), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6503), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6443), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5933), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6503), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6443), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5934), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1834 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6452), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6533), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5934), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6452), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N748), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5933), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6533), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1838 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N748));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9000), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1841 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9431), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9039), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9806), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8603), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9000));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1842 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10137), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9230), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9431), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9987));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1843 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9357), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10137), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9194), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9955));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1844 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1845 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1846 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6357), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1847 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1848 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6296), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1849 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6481), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6357), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6296), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1850 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6210), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1851 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6483), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6210), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6075), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6307), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6075), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6382), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6483), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6307), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1855 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N747), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6481), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6382), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N747));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1858 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8662), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1859 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1860 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1861 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1862 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10197), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1863 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9241), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8865), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8662), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9915), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10197));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1864 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1865 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10058), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1870 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10208), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9850), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10058), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9267), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8970));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1871 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9203), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9241), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10208), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10026));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1872 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1873 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8857), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1874 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1875 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9114), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9305), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1879 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1881 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9469), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9078), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9114), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9305), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9422));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1882 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10172), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9814), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8857), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9504), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9469));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1883 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9165), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8796), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10172), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9008));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1884 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6200), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6142), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6339), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6200), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6142), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6058), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6058));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5907), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1892 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6154), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1893 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6152), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5907), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6154), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1894 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6229), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6033), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6152), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N746), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6339), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6229), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N746));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1899 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1900 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8753), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1901 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1902 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9541), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1903 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9503), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9113), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8753), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9541));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1904 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1908 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9727), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9693), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10145));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1910 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9842), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1912 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8632), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1913 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1914 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9031), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1915 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10236), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9885), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9842), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8632), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9031));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1916 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9997), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9631), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9503), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9727), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10236));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1917 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9964), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9594), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9039), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9814));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1918 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9928), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9964), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9780), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8796));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1919 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10099), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9744), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9165), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9928));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1920 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8788), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9385), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9357), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10099));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1921 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7537), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7352), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7537));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7491), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7352), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7491));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1927 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7902), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1928 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7857), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7902));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1929 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7715), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1930 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7857), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7715));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1931 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1932 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1933 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7816), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1934 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7498), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7816));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1935 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7919), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1936 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7498), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7919));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1937 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9325), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1938 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9186), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8788), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9797), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1939 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9824), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10047), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8706), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9186));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7454), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7836), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7454));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7578), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7331), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7836));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1947 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7691), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7691));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1949 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9424), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9424), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1951 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8726), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10061), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9824), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9311));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1952 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[34]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[33]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10150), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9996), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8726));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1953 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897), .A(N22005), .B(N22003), .CI(N22007));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032), .B(N21818));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1955 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1956 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1957 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9627), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1958 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1959 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9238), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1960 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9248), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9248));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1962 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1963 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1965 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9047), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1966 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8845), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10185), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9238), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9047), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9447));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1967 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[33]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[32]), .A(N22147), .B(N22145), .CI(N22149));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1968 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6562), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1969 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6025), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1970 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6050), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6025), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1971 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6245), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6562), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6050), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6521), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6219), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6521), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6515), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1975 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6435), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6219), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6515), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1976 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[15]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6245), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6435), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I1977 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[33]), .B(N21993), .CI(N21997));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6517), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6410), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6517), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1983 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5883), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1984 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6093), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6410), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5883), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1985 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6068), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1986 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1987 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6366), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6288), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6068), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6366), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1989 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[14]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6093), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6288), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1990 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1991 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6006), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1992 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6039), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1993 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6085), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6006), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6039), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1994 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6442), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1995 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6201), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1996 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6516), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6442), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6201), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1997 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[14]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6085), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6516), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1998 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[14]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I1999 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9292), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2000 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2002 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9946), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9578), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9292), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8698));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8863), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2005 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6582), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2006 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5917), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6582), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6295), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6048), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6367), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6295), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6048), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[13]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5917), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6367), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[13]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2013 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8590), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2014 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9015), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9850), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9078), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8865));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2015 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2017 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2018 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2019 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2020 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10230), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2021 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8602), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9914), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8686), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9947), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10230));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2022 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10034), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9667), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9343), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8602), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9113));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2023 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2025 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9151), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2027 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10205), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2028 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9766), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9379), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9306), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9151), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10205));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2029 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2030 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2031 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9460), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2033 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10090), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6047), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5984), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2038 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6181), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6047), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5984), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6574), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5994), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6082), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6574), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5994), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2044 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N745), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6181), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6082), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2045 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N745));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2046 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2047 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9613), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2048 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9540), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9152), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9460), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10090), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9613));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2049 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9277), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8900), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9766), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8891), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9540));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2050 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9788), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9398), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9277), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9631));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2051 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8981), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8644), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8833), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9015), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9788));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5880), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6141), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6538), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2055 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6031), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5880), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6538), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2058 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6421), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6546), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5913), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6421), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6546), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2061 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N744), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6031), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5913), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2062 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N744));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2063 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9224), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2065 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2066 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2067 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2069 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8820), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10160), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9224), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8785), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2074 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9800), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9226), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9728));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2075 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2076 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2077 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2078 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2079 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2080 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8928), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2081 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9581), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9189), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9067), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9877), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8928));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2082 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9314), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8820), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9800), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9581));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2083 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9049), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9314), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9885), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8900));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2084 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8803), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9049), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8672), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9398));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2085 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9751), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8644), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9594), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8803));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2086 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8949), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8613), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9557), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8981), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9751));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2087 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7721), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2088 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7289), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7289));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7579), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2091 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7516), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2092 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7579), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7516));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2093 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2094 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2095 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9129), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8765), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8949), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9744), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2096 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9548), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8590), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10130), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9129));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10031), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10039), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10039));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2101 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9856), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2105 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10203), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2107 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8608), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10031), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9856), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10203));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2108 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8967), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8629), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8863), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9548), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8608));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2109 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[32]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[31]), .A(N22139), .B(N22137), .CI(N22141));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2110 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[32]), .B(N21973), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[32]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2111 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2112 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839), .A(N20872), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12199), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6250), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6428), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2118 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6467), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6250), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6428), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6140), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2120 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2121 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5881), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2122 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6215), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6140), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5881), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[12]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6467), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6215), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[12]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9523), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9475), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2128 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9896), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8765), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9523), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9475));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6100), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2130 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6283), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6324), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6100), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6283), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5983), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2135 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6179), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2136 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6359), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2137 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6437), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6179), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6359), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2138 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6063), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5983), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6437), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2139 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[11]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6324), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6063), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[11]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8769), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2142 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10063), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9152), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9379), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9914));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2144 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9655), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2146 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10124), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2149 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9617), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9225), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10124), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8717));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2150 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9352), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9617), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10160));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2152 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2153 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10193), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2155 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9064), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9190), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10193), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9582), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2158 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9342), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6436), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6388), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2165 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6573), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6436), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6388), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6301), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6272), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6301), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2168 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6094), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2169 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6394), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6094), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6464), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6394), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N743), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6573), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6464), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N743));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2173 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8850), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2175 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8852), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10194), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9496), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9342), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8850));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2176 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8631), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9950), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9582), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8852));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2177 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9085), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9352), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8631), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8936));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2178 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9819), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9667), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10063), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9085));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9262), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2183 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6289), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6235), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6420), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6289), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6235), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6146), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2187 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6119), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6146), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2188 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6244), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6320), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6119), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6244), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N742), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6420), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6320), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N742));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2193 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2195 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10075), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9262), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10190), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2196 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2197 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8597), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2198 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8818), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2200 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9764), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10050), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2204 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9873), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9764), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10050));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2205 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8663), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10075), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8597), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9873));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2206 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10096), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8663), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9189), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9950));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2207 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9857), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10096), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9701), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8728));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2208 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8841), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10181), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8701), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9440));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2209 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9564), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9173), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9819), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8841));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2210 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7435), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2211 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7738), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7738));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7295), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7315), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7295), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7315));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2216 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9121), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2217 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9121), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2218 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8770), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10108), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9564), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9363), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2219 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9715), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9329), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8613), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8769), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8770));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2221 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9666), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9849), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2224 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8911), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8587), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9715), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9666), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9849));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2225 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9320), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9157), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8911));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2226 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[31]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[30]), .A(N22155), .B(N22153), .CI(N22157));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6262), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2229 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6439), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2230 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5927), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6262), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6439), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5899), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2232 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6466), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2233 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2234 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6213), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6466), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6101), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6135), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5899), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6213), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2236 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[13]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5927), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6135), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2237 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[31]), .B(N21953), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[31]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9090), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9090));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8906), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9083), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2247 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9274), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2249 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8740), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8906), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9083), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9274));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2250 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2251 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9466), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5935), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5988), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2254 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6128), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5988), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6166), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5935), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6128), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2256 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2257 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6537), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2258 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6290), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5895), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6537), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6290), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[10]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6166), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2261 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[10]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2262 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9749), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2263 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2264 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2265 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9525), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10108), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9749), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8727));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2266 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9491), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9098), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9466), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9525));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2267 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9681), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9289), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9519), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8740), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9491));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2268 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[30]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[29]), .A(N22131), .B(N22129), .CI(N22133));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6108), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6292), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2272 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6480), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6108), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6292), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2274 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6454), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2275 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6062), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2276 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5976), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6454), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6062), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2277 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[12]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6480), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5976), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2278 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[30]), .B(N21983), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[30]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8896), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2283 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6009), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6486), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6009), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5968), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6013), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6486), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5968), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6386), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2291 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6136), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2292 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6451), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6386), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6136), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2293 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[9]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6013), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6451), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2294 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[9]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2295 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8979), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9910), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2300 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8962), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2302 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8885), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10225), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9910), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8962));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2303 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9389), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9003), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8885), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10194));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2304 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2305 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9380), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2309 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2310 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9135), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8771), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9533), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9380), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8881));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2311 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8714), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2312 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2314 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10111), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9752), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8714), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9833));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2318 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10161), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2320 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8744), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2321 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9906), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9686), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10161), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8744));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2322 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9657), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9264), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9135), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10111), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9906));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2323 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10131), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9657), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9225), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9983));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2324 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9123), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8760), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8969), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9389), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10131));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2325 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8688), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9493), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9717), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10225));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2326 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9941), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9870), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2333 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9971), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9602), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8915), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9870));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2334 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8957), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8622), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8998), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9941), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9971));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2335 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9689), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9299), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9752), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8771));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10224), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2339 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2341 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9175), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8806), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10224), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9683), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9297));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10083), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2350 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9937), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10083), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9801), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9141));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2351 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8921), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8594), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8626), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9937));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2352 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9426), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8921), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9264));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2353 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9159), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8791), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9003), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8688), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9426));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2354 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9891), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9159), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9735), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8760));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2355 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8872), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10212), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9123), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9891));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7798), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7542), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7798), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7542));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2359 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7760), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7760));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9021), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2363 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9600), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9209), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8872), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10181), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2364 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8619), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9935), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9173), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8979), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9600));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2365 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8592), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8580), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8619));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2366 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10223), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9869), .A(N22235), .B(N22233), .CI(N22237));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2367 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[29]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10223), .B(N22105), .CI(N22109));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2368 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5947), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2369 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5905), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2370 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6138), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5905), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6333), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5947), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6138), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6309), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2374 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6012), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2375 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5893), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6012), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6530), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6309), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5893), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2377 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[11]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6333), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6530), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2378 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[29]), .B(N21963), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[29]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2379 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2381 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2382 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2383 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2384 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10082), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8722), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9888), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9935));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2385 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2386 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2387 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6184), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2388 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6237), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2389 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6373), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6237), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2390 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6407), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6184), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6373), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6541), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2392 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6086), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6541), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6531), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6151), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6086), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6531), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[7]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6407), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6151), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[7]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6340), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2398 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6391), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2399 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6071), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2400 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6522), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6391), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6071), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6558), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6340), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6522), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6234), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5977), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2404 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6306), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6234), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5977), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[8]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6558), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6306), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2406 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[8]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2407 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9199), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8778), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9721), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8657), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2414 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9759), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9373), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8778), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9721), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8657));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9572), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9417), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2420 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2421 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8992), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8653), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9417), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8919));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2422 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9722), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9337), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9759), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8992), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8806));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2423 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8719), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10053), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9722), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9526), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8594));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2424 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10166), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8719), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10021), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9034));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2425 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9923), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9551), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9774), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8791));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7340), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7340));
NAND2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2428 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[18]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2429 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8908), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8581), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9513), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9923), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2430 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9639), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9250), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9199), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10212), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9509), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2433 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9370), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8989), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9882), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9639), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9509));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2434 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9960), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2437 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8651), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9209), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9960), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9697));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2438 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9895), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9895));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2442 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2445 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10060), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2446 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2448 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9336), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10060), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10235));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2449 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9103), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9370), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8651), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8954));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2450 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10049), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9903), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10082), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9103));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2453 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9296), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8918), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9336), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9074), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9133));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2454 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[28]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[27]), .A(N22066), .B(N22064), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9869));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6499), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5980), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6176), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6499), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5980), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6155), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6449), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6379), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6155), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6449), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[10]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6176), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6379), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2464 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[28]), .B(N21913), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[28]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8947), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8947));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9312), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8941), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2482 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8675), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10004), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9312), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8941));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2483 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10117), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10057), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9322), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8675));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9500), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2486 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2487 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2490 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9409), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9500), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9120), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9690));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2491 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9143), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8777), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9409), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9969), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8989));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2492 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9879), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9495), .A(N22251), .B(N22249), .CI(N22253));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2493 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[27]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9879), .B(N22113), .CI(N22117));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6352), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6145), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6534), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6026), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6352), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6534), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5997), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6305), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6226), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5997), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6305), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[9]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6026), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6226), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2503 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[27]), .B(N21893), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[27]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2504 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10118), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9181), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2511 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8814), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10118), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9333), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9181));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9131), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2513 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9611), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9221), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9131));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2514 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9898), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2517 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9794), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9898), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8591));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2518 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8780), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8814), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9794), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9602));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2519 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8746), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10085), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9566), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8780));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2520 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9462), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9072), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9299), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10053));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7564), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7564));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2523 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9197), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9462), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9809));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6576), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6069), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6106), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6576), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6069), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6240), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6469), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6240), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2529 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6511), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6511), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6545), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6469), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[5]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6106), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6545), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[5]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6035), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2535 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6220), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6256), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6035), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6220), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5918), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6380), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5993), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5918), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6380), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2542 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[6]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6256), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5993), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2543 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[6]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2544 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9427), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2545 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8943), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9197), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9427));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10170), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2547 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9676), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9285), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10170), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8581));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2554 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8708), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8933), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8606));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2555 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10152), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9676), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9250), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8708));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2557 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9111), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2558 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2562 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9449), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9058), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9111), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8757), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9304));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2563 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9180), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8813), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10004), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9449), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9022));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2564 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9909), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9532), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10152), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9180));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2565 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[26]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[25]), .A(N22082), .B(N22080), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9495));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6197), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6004), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6294), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6383), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6004), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6294), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2570 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6569), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6197), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6383), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2571 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2572 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6548), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2573 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6150), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6078), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6548), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6150), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[8]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6569), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6078), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2576 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[26]), .B(N21923), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[26]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2578 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2581 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9977), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9904), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8955), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2587 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8658), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9221), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9904), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8955));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2588 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9575), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9028), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9977), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8658));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2589 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9535), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9575), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8653), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9373));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2590 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9499), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9107), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9337), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9535), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10085));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9963), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2592 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10201), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9845), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9499), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9963), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9072));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6423), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5901), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2595 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5944), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6423), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5901), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6325), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6079), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6393), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6325), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6079), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2600 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[4]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5944), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6393), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[4]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8691), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2603 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9958), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8829), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10201), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8691));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2604 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2605 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[18]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8600), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2610 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9709), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9958), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9556), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8600));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2611 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2612 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2613 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2614 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9743), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2617 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8733), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9743), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8750));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2618 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10186), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9285), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9709), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8733));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10093), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8926), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2623 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9486), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9093), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8610), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10093), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8926));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2624 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9217), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8846), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10040), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9486), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9058));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2625 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9942), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9571), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9792), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10186), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9217));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2626 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[25]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[24]), .A(N22123), .B(N22121), .CI(N22125));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6045), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6230), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6416), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6045), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6230), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2630 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5908), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5998), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6396), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5908), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5998), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6346), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5991), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6346), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2635 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5909), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6396), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5991), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[7]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6416), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5909), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2637 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[25]), .B(N21903), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[25]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2638 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2642 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9356), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2643 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2644 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10087), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2645 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9746), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9360), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9547), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9356), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10087));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2646 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2647 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2653 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9383), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8999), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9756), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9609), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8812));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2654 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8627), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9411), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9383), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10155));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2655 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8598), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8627), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9145));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2656 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10231), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9880), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9201), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8598), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9107));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6276), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6455), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6496), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6276), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6455), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6559), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6228), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5910), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6228), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2663 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6243), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6559), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5910), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2664 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[3]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6496), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6243), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[3]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9659), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2667 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9234), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8860), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9845), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10231), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9659));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9164), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2672 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8977), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8641), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9234), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9164), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9913));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2673 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10217), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9862), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8977), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9324));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9733), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8596), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2678 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8768), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9591), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9733), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8596));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2679 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9257), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10068), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8768), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9093));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2680 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9976), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9608), .A(N22219), .B(N22217), .CI(N22221));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2681 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[24]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[23]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9976), .B(N22097), .CI(N22101));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5876), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6401), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6083), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6401), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6269), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5876), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6083), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2687 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6246), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6193), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6543), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6193), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6462), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6246), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6543), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[6]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6269), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6462), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2692 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[24]), .B(N21943), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[24]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9156), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8975), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9726), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2703 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9011), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8670), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9156), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8975), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9726));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10174), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8620), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9371), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2710 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9192), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8620), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10104), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9371));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2714 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10153), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2717 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2719 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9952), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10153), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9216));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2720 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10126), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9768), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8680), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9952));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2721 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9346), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8965), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9183), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10126), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9944));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2722 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9308), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8930), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10174), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9346), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6121), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6311), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6348), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6121), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6311), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6081), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6463), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6081), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6092), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6463), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2729 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[2]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6348), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6092), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[2]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8887), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2732 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9270), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9880), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9308), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8887));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8798), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9537), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2737 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9991), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9270), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8798), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9537));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2738 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9521), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9991), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8641));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2743 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9784), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8860), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9348), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9908));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2744 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8588), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9360), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9784), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10103));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2745 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10011), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9646), .A(N22211), .B(N22209), .CI(N22213));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2746 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[23]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10011), .B(N22072), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9608));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6434), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5914), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6114), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6434), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5914), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6095), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6392), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6317), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6095), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6392), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[5]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6114), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6317), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2755 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[23]), .B(N21933), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[23]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2757 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8790), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9340), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2763 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9042), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8695), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8790), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8639), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9340));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2765 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2766 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2767 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2768 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9647), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2769 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2770 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2771 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2772 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9793), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2773 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9553), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9162), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8990), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9793));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9359), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2777 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8793), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9359), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9936));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2778 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8972), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9553), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8793), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8822));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2779 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9155), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8787), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8999), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9978), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8972));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2780 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10092), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9730), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9430), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9155), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8965));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2781 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2782 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8650), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2783 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8642), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2786 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9901), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8650), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8642), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9408));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2787 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2789 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8611), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9901), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8847), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10132));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2790 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9739), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9585), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8635));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2791 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9917), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9543), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8787), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9768), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9739));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2794 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9258), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2795 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2796 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10187), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2800 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9266), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9970));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2801 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8916), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8589), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9258), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10187), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9266));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2802 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9326), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9162), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8916), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9925));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2803 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9662), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2804 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8762), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10098), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9355), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9326), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9662));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2805 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8938), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9543), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8693), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8762));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2806 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9116), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9730), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9917), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8938));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2807 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10059), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9695), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8930), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10092), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9116));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2810 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10029), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9663), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10059), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9148));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2811 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8800), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10140), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10029), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9625));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8966), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2816 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9815), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9434), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8966), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9531));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2817 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9559), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9169), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8670), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9815), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9394));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2818 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9291), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8914), .A(N22227), .B(N22225), .CI(N22229));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2819 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[22]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9291), .B(N22040), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9646));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6287), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6465), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2822 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5953), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6287), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6465), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2823 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5929), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6242), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6162), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5929), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6242), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[4]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5953), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6162), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2827 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[22]), .B(N21883), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[22]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2834 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9852), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9695), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9954), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8959));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9779), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5960), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2838 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6156), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6195), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5960), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6156), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6258), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2841 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5887), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2842 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5912), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2843 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6318), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5887), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5912), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2844 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5926), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6258), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6318), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2845 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[1]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6195), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5926), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2846 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[1]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2847 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9876), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2848 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2849 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8783), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2850 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9080), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8725), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9779), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9876), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8783));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2851 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8835), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10176), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9852), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9080), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9663));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2855 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10129), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2858 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8868), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10209), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10129), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9138));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2859 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9597), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9205), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8695), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8868), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9434));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2860 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8615), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9930), .A(N22243), .B(N22241), .CI(N22245));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2861 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[21]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8615), .B(N22048), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8914));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2862 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6133), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2863 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2864 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6321), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2865 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6508), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6133), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6321), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6334), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6091), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6008), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6334), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6091), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2870 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[3]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6508), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6008), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2871 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[21]), .B(N21853), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[21]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2872 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2873 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2874 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9589), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2875 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10122), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9770), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2879 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8904), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10238), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9589), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10122), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9770));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2881 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6514), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6372), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2882 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5999), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2883 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6040), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6514), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5999), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2884 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6174), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6107), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6174), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6163), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6477), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6107), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6163), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[0]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6040), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6477), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[0]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9101), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2892 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9393), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2893 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9887), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8756), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9101), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9393));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2894 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9633), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9244), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8904), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9887), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8725));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2899 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2900 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8773), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2901 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9670), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9280), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8625), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9945), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8773));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2902 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8673), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9999), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9472), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9670), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10209));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2903 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8645), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9966), .A(N22316), .B(N22314), .CI(N22318));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2904 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[20]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8645), .B(N22056), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9930));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5973), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6164), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6322), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2908 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6362), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5973), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6164), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6177), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2910 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6450), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5925), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6450), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2912 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6555), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6177), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5925), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2913 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[2]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6362), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6555), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2914 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[20]), .B(N21873), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[20]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2915 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2916 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2917 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2918 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10078), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2919 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2920 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9006), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2921 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9704), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10078), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8605), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9006));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9196), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9761), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2927 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9387), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2928 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8730), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9196), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9761), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9387));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2929 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8703), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9704), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8730));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2930 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2931 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9939), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2932 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2933 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2934 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2935 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2936 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9480), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9089), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9939), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9577), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10116));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2937 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9443), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9052), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10238), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9480), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9280));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2938 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9402), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9244), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8703), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9443));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2939 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[19]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[18]), .A(N22260), .B(N22258), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9966));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6528), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6010), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6204), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6528), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6010), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6027), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6476), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6403), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6027), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6476), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[1]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6204), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6403), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2947 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[19]), .B(N21863), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[19]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2949 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6378), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6556), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2951 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6052), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6378), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6556), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2952 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6570), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2953 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6331), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6252), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6570), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6331), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2955 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[0]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6052), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6252), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2956 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2957 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9825), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2958 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2959 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2960 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2962 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10024), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9658), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9023), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2963 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9685), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9522), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10024), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8589));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8890), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2965 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10072), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8945), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9685), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8890));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2966 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2967 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8666), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2968 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9517), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9126), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10098), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10072), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8666));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2969 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2970 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2971 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9377), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9001), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2975 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8583), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8823), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9377), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9001));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2976 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10214), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9859), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9318), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9517), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8583));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2977 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9187), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9755), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2983 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9288), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8910), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9568), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9187), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9755));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2984 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9253), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8873), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9288), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9089));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2985 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10182), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9821), .A(N22324), .B(N22322), .CI(N22326));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2986 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[18]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10182), .B(N22306), .CI(N22310));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2987 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910), .A(N22278), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[18]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2989 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2990 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8676), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2991 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2992 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2993 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9450), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2994 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10144), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9786), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8676), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8827), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9450));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2995 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9037), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8888), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10144), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9658));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2996 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9878), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I2997 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8715), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9293), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9037), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9878));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2998 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I2999 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9989), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3000 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9096), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8736), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8715), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9989));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3002 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8996), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9178), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3005 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9865), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9490), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8996), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9178));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3006 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10043), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9678), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9126), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9096), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9865));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8659), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10165), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8816), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3013 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8880), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10165), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8816));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3014 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9810), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3015 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10003), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3017 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9303), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10003));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3018 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3019 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3020 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9171), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9303), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10218), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9786));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3021 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3022 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9812), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8690), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9171), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9105));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3023 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9622), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3025 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9458), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9065), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10046), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9812), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9622));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3027 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9367), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3028 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9650), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9259), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9458), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9367), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8736));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3029 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9060), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8880), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9650));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3030 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10005), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9642), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10043), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9060));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3031 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[17]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[16]), .A(N22270), .B(N22268), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9821));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3033 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[17]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[17]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9975), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9423), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3038 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9593), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9975), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9423));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10149), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9614), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3044 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9798), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3045 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8643), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9961), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10149), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9614), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9798));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3046 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9985), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9619), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9593), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9065), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8643));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3047 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9421), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9030), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10220), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9259));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3048 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3049 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3050 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3051 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10156), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9863), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3055 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9059), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3058 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9485), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3061 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9968), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8707), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9035), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9485));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3062 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10056), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9863), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9059), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9968));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3063 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10020), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3065 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10041), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3066 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8898), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10020), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10041));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3067 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9094), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3069 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9265), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3074 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3075 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9791), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10226), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10067));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3076 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9339), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8960), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8734), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9265), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9791));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3077 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9665), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10234), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9094), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9339));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3078 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8987), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8647), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8898), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9665));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3079 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9076), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8721), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8925), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8987));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3080 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9934), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8802), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10056), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9076));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3081 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3082 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9229), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3083 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8831), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10169), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9428), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9934), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9229));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3084 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9227), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10156), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8831));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3085 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3086 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9807), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3087 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3088 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8655), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3091 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10195), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9838), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8655), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9981));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3092 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8682), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9227), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10195), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9490));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3093 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9829), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9453), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8910), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8682));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3094 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[15]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8710), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9453));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3095 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[16]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[15]), .A(N22288), .B(N22286), .CI(N22290));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3096 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[16]));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12443), .A0N(N22034), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[15]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10081), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3101 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8952), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9561), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10081), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8858));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3105 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3107 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9222), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3108 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9719), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9332), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9032), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9606), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9222));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3109 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9361), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10169), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8952), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9719));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3110 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9004), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8665), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9838), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9361));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3111 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[14]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10014), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9004), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9030));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3112 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307), .A(N22294), .B(N22296));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9334), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3114 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9848), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9465), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9334), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3117 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8743), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9848), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9414), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8618));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3118 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10106), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9748), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8743), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9198), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9961));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3119 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[13]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10106), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9619), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8665));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3120 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[13]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3121 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3122 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8851), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8621), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3128 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9754), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9369), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8621), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8647), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9840));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3129 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9629), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9237), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9026), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8851), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9754));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3130 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9214), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3135 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3136 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8862), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9214), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10198), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8687));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3137 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9494), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9100), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9629), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8862), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9332));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3138 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[12]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8978), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9748));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3139 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12391), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[12]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10191), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3142 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3144 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3146 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8775), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10191), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10017), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8679));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3147 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8671), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8775), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9465), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10204));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3148 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[11]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8671), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10079), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9100));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3149 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[11]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9563), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3152 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9461), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3153 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8697), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9563), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9273), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9461));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9653), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9831), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3158 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9439), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9653), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9831));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3159 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9530), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9137), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8697), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9439));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3160 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[10]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9530), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9237), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9995));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[10]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3165 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10089), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9725), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8960), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9068));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3168 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10179), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10089), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10007), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10033));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3169 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[9]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10115), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10179), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9137));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12191), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[9]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3173 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9263), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3175 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9787), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3176 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3177 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8716), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3178 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8808), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10151), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9787), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9405), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8716));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3179 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9110), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9263), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8808));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3180 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[8]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9046), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9110), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9817));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11916), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[8]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3183 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3186 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9570), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9177), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8882), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9062));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3187 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[7]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9725), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8749));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3188 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12272), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[7]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3193 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10001), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9014), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9492), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10051));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3194 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[6]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10151), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10001), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9177));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3195 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11993), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[6]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3196 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3197 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10211), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9855), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9998), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3198 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10222), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3200 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[5]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10211), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10222), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9638));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[5]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9871), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3206 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[4]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9871), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9687), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9855));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3207 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12075), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[4]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3208 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9240), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3209 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3210 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9295), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3211 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[3]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9295));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[3]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10207), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3214 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[2]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[2]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3216 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3217 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3218 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[1]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3219 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12037), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12155), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12201), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[2]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[2]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12295), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[3]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3221 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11879), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12433), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12037), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12295));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12269), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12075), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11879), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[4]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[4]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[5]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3224 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12025), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12353), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12269), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12213));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3225 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12340), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11993), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12025), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[6]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[6]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3226 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[7]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12011), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12272), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12340), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12130));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12241), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11916), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12011), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[8]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[8]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3229 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[9]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3230 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11847), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12191), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12241), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12051));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11986), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11840), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11847), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[10]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[10]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3232 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[11]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3233 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12134), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12112), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11986), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11974));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3234 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12203), .A0(N22205), .A1(N22199), .B0(N22201), .B1(N22203));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[13]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3236 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12169), .A(N22294), .B(N22296));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12425), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307), .A1(N22194), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12169));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12388), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307), .A1(N22091), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12203), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12425));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12443), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12388));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12445), .A(N22034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[15]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12087), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[16]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12305), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12445), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12087));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12368), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[17]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12221), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12368), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12005));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11900), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12305), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12221));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3247 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12082), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12254), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11900));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12283), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3249 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12419), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12082), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12283));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3250 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3251 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3254 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3256 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3257 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3258 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3261 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3262 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3263 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3264 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3266 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3272 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3274 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3275 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3276 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3277 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3278 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032), .B(N21818));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12327), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049), .B0(N21559));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3283 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329), .A0(N20872), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436), .B0(N20876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3291 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3292 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3293 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3294 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3295 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3300 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928));
AO22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3302 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11954), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3303 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12004), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11954));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3304 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12057), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329), .B0(N20654));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3305 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12199), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12057));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3309 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3310 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3311 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3312 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11869), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023), .A(N21570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136), .A(N21060), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3318 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3320 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11926), .A(N19751), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3321 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3322 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3323 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3324 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3325 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3326 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3333 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3334 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3339 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3341 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888), .A0(N21570), .A1(N21559), .B0(N21574));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997), .A0(N21060), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888), .B0(N21064));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3350 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3351 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3352 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3353 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12117), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12310), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12117));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12367), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12310));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12417), .A0(N19751), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050), .B0(N19755));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11846), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11926), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12417));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3359 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[48]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11846), .B(N19431));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18865), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[48]), .B(N19158));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18865));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3363 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3364 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12222), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3365 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863), .A(N21306), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3366 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3367 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3368 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12280), .A(N20628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3369 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3370 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3374 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3375 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3377 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3378 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357), .A0(N21306), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243), .B0(N21310));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3379 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3381 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12031), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3382 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12086), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12031));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3383 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12141), .A0(N20628), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410), .B0(N20632));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3384 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12196), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12280), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12141));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3385 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12234), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3386 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[47]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12196), .B(N20265));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3387 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[47]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3388 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3389 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3390 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11950), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3392 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12001), .A(N20621), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3398 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3399 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3400 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3404 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3406 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3407 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12394), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12444), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12394));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11866), .A0(N20621), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129), .B0(N20625));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11922), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12001), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11866));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11829), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[46]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11922), .B(N20290));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[46]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3414 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12363), .A(N20609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3420 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3421 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3422 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12168), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12219), .A0(N20609), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859), .B0(N20613));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12277), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12363), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12219));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12040), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[45]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12277), .B(N20285));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[45]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3428 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027), .A(N20912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3429 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12083), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3434 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11892), .A0(N20912), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997), .B0(N20916));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11947), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11892));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3437 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11999), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12083), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11947));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3438 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12259), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[44]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11999), .B(N20275));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[44]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3442 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390), .A(N20899), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3445 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3446 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12246), .A0(N20899), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357), .B0(N20903));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12301), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12246));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3450 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12359), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12440), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12301));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11852), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[43]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12359), .B(N20260));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[43]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111), .A(N20886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12165), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11973), .A0(N20886), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078), .B0(N20890));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12024), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11973));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12080), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12165), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12024));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12063), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[42]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12080), .B(N20280));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11889), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12386), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12438), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11889), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12386));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12285), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[41]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12438), .B(N20270));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[41]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12244), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12106), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12161), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12244), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12106));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11872), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[40]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12161), .B(N20295));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[40]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3482 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11837), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3483 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11887), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11969), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11837));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12089), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[39]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11887), .B(N20355));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3486 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[39]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3487 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12326), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12187), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12242), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12326), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12187));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12309), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[38]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12242), .B(N20382));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[38]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3493 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11912), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11966), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12048), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11912));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11895), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[37]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11966), .B(N20370));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[37]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12268), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12323), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12407), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12268));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3503 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12114), .AN(N21559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3504 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[36]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12323), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12114));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[36]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12061), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12333), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[35]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12061), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12333));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[35]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11930), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11919), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3514 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[34]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11930), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11919));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[34]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12133), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[33]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12133));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3519 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[33]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3520 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12356), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[32]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12356));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[32]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11941), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[31]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11941));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3529 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[31]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12158), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12158));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[30]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12380), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3535 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12380));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[29]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11963), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11963));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3542 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13289), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3543 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3544 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13344), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13289), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13325));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13285), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13344), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13285));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3547 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12181), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[27]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12181));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[27]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12402), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12402));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3554 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13287), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3555 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13305), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13335), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13287));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13297), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3557 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3558 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13330), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13297), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13313));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13277), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13305), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13330));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13321), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13312), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13321), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3562 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13277), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13312));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3563 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11985), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3564 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11985));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[25]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13278), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13314), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13331), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13278), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13314));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13322), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3570 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13340), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3571 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13275), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13322), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13340));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3572 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13317), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13331), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13275));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3573 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13347), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13300), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13347), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13281));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3576 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13290), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3578 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13326), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13290), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13306));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13272), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13300), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13326));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13298), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13317), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13272));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3581 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13315), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13270), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13315), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13333));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13342), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13336), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13296), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13342), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13336));
OA21X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13332), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13270), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13296));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3588 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13298), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13332));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3589 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13413), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13413), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3592 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13410), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3595 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[0]));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3600 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3603 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3604 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3605 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13478), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13430), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3610 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3611 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3612 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3613 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13428), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13478), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3614 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13529), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13428), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0]));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3623 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3624 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3625 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N683), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13529), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N683));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3627 (.Y(x[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N739), .B(N18245), .S0(N22962));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3630 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3635 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13449), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13550), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3638 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13548), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13449), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3642 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13496), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13548), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3643 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3644 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3645 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3646 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3647 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N682), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13496), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N738), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N682));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3652 (.Y(x[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N738), .B(N18245), .S0(N22964));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3653 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3654 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3655 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3656 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13566), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13514), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13566), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13460), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13514), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3663 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3664 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N681), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13460), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N737), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N681));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3666 (.Y(x[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N737), .B(N18245), .S0(N22966));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13534), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13477), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13534), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13429), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13477), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N680), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13429), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N736), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N680));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3679 (.Y(x[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N736), .B(N18245), .S0(N22965));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13448), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13549), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13448), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N679), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13549), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N679));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3687 (.Y(x[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N735), .B(N18245), .S0(N22963));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13565), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13516), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13565), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N678), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13516), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N678));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3695 (.Y(x[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N734), .B(N18245), .S0(N22964));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13533), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13480), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13533), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N677), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13480), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N733), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N677));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3703 (.Y(x[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N733), .B(N18245), .S0(N22963));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13500), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13451), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13500), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N732), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13451));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3708 (.Y(x[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N732), .B(N18245), .S0(N22965));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13568), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3710 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N731), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13568));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3711 (.Y(x[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N731), .B(N18245), .S0(N22965));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13535), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N730), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13535));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3714 (.Y(x[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N730), .B(N18245), .S0(N22964));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13502), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N729), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13502));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3717 (.Y(x[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N729), .B(N18245), .S0(N22962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13466), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3719 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N728), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13466));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3720 (.Y(x[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N728), .B(N18245), .S0(N22962));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3721 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13436), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N727), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13436));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3723 (.Y(x[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N727), .B(N18245), .S0(N22964));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13556), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N726), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13556));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3726 (.Y(x[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N726), .B(N18245), .S0(N22966));
AOI22XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13522), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N725), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13522));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3729 (.Y(x[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N725), .B(N18245), .S0(N22965));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18874));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3732 (.Y(x[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N724), .B(N18245), .S0(N22962));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N723), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3734 (.Y(x[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N723), .B(N18245), .S0(N22963));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N722), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3736 (.Y(x[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N722), .B(N18245), .S0(N22963));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N721), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3738 (.Y(x[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N721), .B(N18245), .S0(N22963));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N720), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3740 (.Y(x[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N720), .B(N18245), .S0(N22965));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N719), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3742 (.Y(x[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N719), .B(N18245), .S0(N22966));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N718), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3744 (.Y(x[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N718), .B(N18245), .S0(N22964));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3745 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N717), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3746 (.Y(x[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N717), .B(N18245), .S0(N22962));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N595), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N585));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N595));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N713), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3751 (.Y(x[27]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N713), .B(N18406), .S0(N18402));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N712), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3753 (.Y(x[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N712), .B(N18406), .S0(N18402));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N711), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3755 (.Y(x[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N711), .B(N18406), .S0(N18402));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N710), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3757 (.Y(x[24]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N710), .B(N18406), .S0(N18402));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N709), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3759 (.Y(x[23]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N709), .B(N18406), .S0(N18402));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13872), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_3_I3761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707));
NOR4BBX1 DFT_compute_cynw_cm_float_cos_E8_M23_3_I3763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[31]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13872), .BN(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N493), .C(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[8]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[7]));
EDFFHQX1 x_reg_28__I3792 (.Q(x[28]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__I3794 (.Q(x[30]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[30]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__I3795 (.Q(x[31]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[31]), .E(bdw_enable), .CK(aclk));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[0] = x[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[1] = x[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[2] = x[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[3] = x[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[4] = x[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[5] = x[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[6] = x[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[7] = x[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[8] = x[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[9] = x[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[10] = x[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[11] = x[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[12] = x[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[13] = x[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[14] = x[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[15] = x[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[16] = x[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[17] = x[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[18] = x[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[19] = x[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[20] = x[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[21] = x[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[22] = x[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[23] = x[23];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[24] = x[24];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[25] = x[25];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[26] = x[26];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[27] = x[27];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[28] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[29] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[30] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[4] = 1'B0;
assign x[29] = x[28];
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urX3TAHWrBlO : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



