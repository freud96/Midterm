/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:30 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_mul_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x;
wire  DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__33;
wire [9:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34;
wire  DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__41,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__42;
wire [47:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43;
wire [7:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54;
wire  DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__60,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__61,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N267,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N268,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N269,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N270,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N272,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N273,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N274,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N276,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1314,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1318,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1338,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1340,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1361,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1369,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1372,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1374,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1378,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1380,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1383,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1389,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1393,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1425,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1429,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1451,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1483,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1485,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1489,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1491,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1494,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1500,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1504,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1551,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1552,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1553,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1554,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1555,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1556,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1557,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1558,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1559,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1561,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1563,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1564,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1566,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1567,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1569,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1570,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1571,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1572,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1574,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1576,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1577,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1578,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1579,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1580,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1581,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1582,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1583,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1584,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1585,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1586,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1587,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1588,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1589,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1590,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1591,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1592,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1593,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1594,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1595,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1596,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1597,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1600,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1601,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1602,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1603,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1604,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1605,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1606,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1607,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1608,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1609,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1610,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1611,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1612,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1613,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1614,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1616,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1617,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1618,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1619,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1620,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1622,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1624,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1625,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1626,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1627,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1628,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1631,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1632,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1633,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1634,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1636,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1637,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1638,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1639,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1640,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1641,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1642,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1643,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1644,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1645,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1646,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1647,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1648,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1650,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1651,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1652,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1654,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1655,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1656,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1657,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1659,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1660,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1661,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1662,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1664,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1665,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1666,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1667,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1668,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1669,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1670,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1671,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1673,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1674,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1675,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1676,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1677,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1678,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1679,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1680,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1681,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1683,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1684,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1685,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1686,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1687,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1690,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1691,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1692,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1693,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1694,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1696,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1698,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1699,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1700,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1701,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1703,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1704,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1705,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1707,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1708,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1709,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1710,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1711,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1712,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1713,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1714,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1715,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1716,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1717,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1718,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1719,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1720,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1721,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1722,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1723,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1725,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1727,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1728,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1729,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1730,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1731,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1733,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1734,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1735,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1736,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1737,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1738,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1739,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1740,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1741,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1742,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1743,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1744,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1745,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1746,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1747,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1748,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1750,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1751,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1752,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1753,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1754,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1755,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1757,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1759,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1760,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1761,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1762,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1763,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1764,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1766,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1767,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1769,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1771,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1773,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1774,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1775,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1776,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1779,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1780,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1781,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1782,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1783,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1784,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1785,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1786,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1787,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1788,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1791,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1792,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1793,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1796,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1799,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1800,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1801,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1802,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1804,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1805,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1806,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1807,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1808,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1809,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1810,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1811,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1812,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1813,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1815,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1816,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1817,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1818,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1819,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1821,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1822,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1824,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1825,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1826,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1827,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1828,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1830,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1832,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1834,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1835,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1837,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1838,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1839,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1840,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1841,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1842,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1843,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1844,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1845,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1847,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1848,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1849,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1852,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1853,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1855,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1856,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1858,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1859,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1860,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1861,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1862,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1863,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1864,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1865,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1866,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1867,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1869,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1870,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1872,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1873,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1874,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1875,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1876,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1877,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1878,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1879,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1880,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1881,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1882,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1883,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1884,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1885,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1886,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1887,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1888,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1889,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1890,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1891,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1892,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1893,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1894,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1896,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1897,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1899,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1900,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1903,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1905,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1906,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1907,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1908,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1909,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1910,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1911,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1912,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1913,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1914,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1915,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1916,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1918,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1919,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1920,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1921,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1922,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1924,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1925,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1926,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1927,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1929,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1930,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1932,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1934,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1935,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1936,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1938,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1939,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1940,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1942,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1944,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1946,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1947,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1949,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1950,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1951,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1952,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1953,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1954,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1956,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1957,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1958,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1959,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1960,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1961,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1962,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1963,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1964,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1965,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1966,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1967,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1968,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1969,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1972,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1973,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1974,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1975,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1976,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1977,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1978,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1979,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1980,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1981,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1982,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1983,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1984,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1985,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1986,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1987,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1988,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1990,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1991,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1993,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1994,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1995,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1996,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1997,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1998,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1999,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2000,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2001,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2003,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2004,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2005,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2007,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2008,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2009,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2010,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2011,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2012,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2013,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2014,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2015,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2016,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2017,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2018,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2019,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2020,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2022,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2023,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2024,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2026,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2027,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2028,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2029,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2030,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2031,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2032,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2034,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2035,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2036,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2037,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2038,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2039,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2040,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2041,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2042,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2043,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2044,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2046,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2047,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2048,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2051,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2052,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2053,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2055,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2056,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2057,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2058,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2060,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2061,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2062,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2064,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2065,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2066,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2067,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2069,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2070,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2071,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2073,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2074,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2075,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2076,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2077,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2079,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2080,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2082,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2083,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2084,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2085,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2086,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2087,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2089,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2090,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2091,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2092,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2093,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2094,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2095,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2096,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2097,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2098,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2101,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2102,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2103,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2104,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2105,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2106,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2108,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2109,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2110,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2111,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2112,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2113,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2114,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2116,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2117,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2118,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2119,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2121,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2123,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2124,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2125,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2126,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2127,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2128,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2129,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2130,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2131,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2132,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2133,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2134,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2136,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2137,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2138,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2140,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2141,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2143,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2144,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2145,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2148,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2149,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2151,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2153,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2154,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2156,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2157,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2158,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2160,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2161,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2162,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2163,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2164,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2165,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2166,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2167,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2168,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2170,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2171,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2172,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2173,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2174,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2175,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2176,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2177,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2179,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2180,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2181,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2183,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2184,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2185,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2186,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2187,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2188,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2190,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2193,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2194,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2195,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2197,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2198,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2199,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2200,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2203,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2204,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2205,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2207,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2208,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2209,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2210,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2211,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2212,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2213,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2214,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2215,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2216,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2217,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2219,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2220,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2221,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2223,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2224,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2225,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2226,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2227,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2228,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2229,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2231,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2233,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2234,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2235,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2236,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2238,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2239,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2240,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2242,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2243,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2244,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2246,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2247,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2248,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2249,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2250,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2251,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2253,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2254,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2255,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2256,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2257,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2258,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2259,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2260,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2262,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2263,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2264,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2265,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2266,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2267,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2269,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2270,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2271,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2272,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2273,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2274,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2276,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2277,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2278,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2279,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2280,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2282,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2283,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2284,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2286,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2287,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2288,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2290,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2291,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2292,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2293,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2295,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2296,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2298,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2299,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2300,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2302,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2303,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2304,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2305,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2306,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2308,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2309,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2310,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2311,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2313,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2314,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2315,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2317,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2318,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2319,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2320,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2321,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2322,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2324,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2325,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2326,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2328,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2329,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2332,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2333,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2334,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2336,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2337,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2338,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2339,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2340,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2341,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2342,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2343,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2344,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2345,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2346,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2347,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2348,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2350,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2352,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2353,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2355,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2356,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2357,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2358,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2360,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2361,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2362,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2363,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2364,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2365,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2366,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2367,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2368,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2369,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2370,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2371,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2373,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2374,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2376,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2377,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2378,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2379,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2380,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2382,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2383,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2384,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2385,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2386,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2387,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2388,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2389,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2390,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2391,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2392,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2393,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2395,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2396,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2397,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2398,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2401,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2402,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2404,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2405,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2406,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2407,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2409,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2410,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2411,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2412,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2413,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2414,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2415,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2416,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2417,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2419,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2420,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2421,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2422,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2424,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2425,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2426,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2427,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2428,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2429,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2430,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2431,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2432,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2434,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2435,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2436,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2437,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2438,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2439,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2441,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2442,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2443,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2444,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2445,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2446,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2448,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2451,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2452,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2454,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2455,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2456,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2457,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2459,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2460,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2461,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2463,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2464,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2465,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2466,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2467,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2468,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2469,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2471,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2473,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2474,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2475,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2476,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2477,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2478,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2479,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2481,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2482,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2483,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2484,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2485,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2486,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2487,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2488,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2490,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2491,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2492,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2493,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2494,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2495,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2497,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2498,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2499,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2500,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2501,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2502,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2503,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2505,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2506,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2507,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2508,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2509,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2511,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2512,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2514,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2515,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2516,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2517,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2518,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2519,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2521,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2522,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2523,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2524,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2525,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2526,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2527,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2529,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2531,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2532,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2533,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2534,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2535,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2536,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2537,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2538,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2540,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2542,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2543,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2545,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2546,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2547,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2548,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2550,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2551,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2553,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2554,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2555,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2557,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2558,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2559,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2560,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2561,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2562,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2563,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2564,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2565,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2566,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2567,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2568,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2569,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2571,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2572,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2574,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2575,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2576,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2577,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2579,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2580,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2581,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2582,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2585,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2586,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2588,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2589,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2590,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2591,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2592,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2593,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2594,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2595,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2596,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2597,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2600,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2601,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2602,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2603,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2604,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2605,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2606,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2608,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2610,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2611,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2612,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2613,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2614,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2615,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2616,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2617,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2618,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2619,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2620,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2624,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2625,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2626,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2627,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2628,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2629,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2631,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2632,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2633,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2634,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2635,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2637,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2638,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2640,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2641,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2642,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2643,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2644,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2645,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2646,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2648,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2650,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2651,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2652,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2653,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2654,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2655,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2657,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2658,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2659,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2661,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2662,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2663,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2664,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2665,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2666,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2667,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2668,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2669,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2672,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2673,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2674,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2675,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2676,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2678,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2679,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2680,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2681,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2683,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2684,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2685,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2686,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2687,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2689,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2690,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2691,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2692,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2693,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2695,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2696,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2698,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2699,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2700,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2701,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2702,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2703,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2704,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2707,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2708,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2709,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2710,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2711,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2713,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2714,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2717,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2719,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2721,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2722,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2723,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2724,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2725,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2727,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2728,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2730,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2731,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2732,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2733,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2734,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2735,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2736,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2737,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2738,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2739,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2740,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2742,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2743,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2744,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2745,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2748,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2749,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2750,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2751,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2752,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2754,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2755,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2756,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2757,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2758,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2760,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2761,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2763,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2764,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2765,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2766,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2767,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2768,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2769,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2770,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2771,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2772,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2773,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2774,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2775,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2776,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2778,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2779,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2780,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2781,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2782,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2783,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2784,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2785,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2786,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2788,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2789,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2790,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2792,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2793,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2794,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2795,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2796,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2797,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2798,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2799,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2800,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2803,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2804,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2805,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2807,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2808,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2809,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2810,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2811,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2813,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2814,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2815,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2816,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2817,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2818,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2819,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2820,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2821,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2823,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2824,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2825,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2827,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2828,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2829,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2830,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2833,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2834,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2836,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2837,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2838,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2839,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2840,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2841,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2842,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2843,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2844,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2845,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2846,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2847,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2849,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2850,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2851,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2852,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2853,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2854,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2855,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2856,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2857,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2859,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2860,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2861,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2862,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2863,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2864,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2865,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2867,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2868,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2869,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2872,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2873,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2874,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2875,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2876,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2878,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2879,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2880,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2882,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2883,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2884,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2885,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2886,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2887,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2888,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2889,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2890,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2892,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2893,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2894,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2895,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2896,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2897,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2898,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2899,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2900,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2901,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2903,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2904,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2906,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2907,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2908,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2909,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2910,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2913,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2914,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2915,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2916,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2917,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2918,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2919,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2920,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2922,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2923,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2924,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2925,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2926,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2927,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2928,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2931,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2932,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2933,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2934,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2935,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2936,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2937,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2939,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2940,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2941,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2942,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2944,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2945,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2946,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2947,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2948,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2949,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2950,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2951,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2952,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2953,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2955,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2956,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2957,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2958,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2959,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2962,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2963,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2964,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2965,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2966,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2968,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2969,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2970,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2971,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2972,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2973,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2974,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2975,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2976,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2979,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2980,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2981,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2982,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2983,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2985,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2986,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2987,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2988,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2989,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2990,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2991,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2993,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2994,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2995,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2996,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2997,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2998,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2999,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3000,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3001,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3003,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3004,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3005,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3007,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3008,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3009,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3010,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3012,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3013,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3014,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3015,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3016,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3017,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3018,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3019,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3020,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3021,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3022,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3023,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3025,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3026,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3027,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3028,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3030,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3031,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3034,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3035,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3036,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3037,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3039,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3040,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3041,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3042,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3043,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3044,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3046,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3047,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3048,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3049,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3051,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3052,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3053,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3054,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3055,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3057,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3058,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3059,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3061,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3063,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3064,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3065,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3067,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3069,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3070,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3071,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3073,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3075,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3076,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3078,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3079,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3080,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3081,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3082,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3083,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3086,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3087,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3088,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3089,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3090,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3092,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3093,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3094,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3096,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3097,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3098,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3100,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3101,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3102,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3103,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3104,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3105,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3107,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3108,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3109,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3110,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3111,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3112,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3113,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3115,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3116,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3117,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3118,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3119,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3120,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3121,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3122,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3124,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3125,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3126,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3127,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3128,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3130,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3131,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3133,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3134,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3135,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3136,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3137,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3138,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3139,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3140,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3141,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3142,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3143,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3144,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3147,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3149,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3150,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3151,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3152,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3153,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3155,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3156,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3158,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3159,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3160,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3161,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3162,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3163,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3164,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3165,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3166,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3167,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3168,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3169,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3170,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3171,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3173,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3174,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3175,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3176,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3177,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3178,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3179,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3181,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3182,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3183,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3185,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3186,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3187,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3188,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3189,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3191,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3192,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3193,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3194,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3195,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3196,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3197,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3198,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3199,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3200,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3201,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3203,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3205,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3206,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3208,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3209,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3210,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3211,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3212,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3213,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3215,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3216,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3217,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3219,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3220,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3221,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3222,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3223,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3224,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3225,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3226,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3227,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3229,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3230,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3231,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3232,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3233,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3234,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3235,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3238,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3239,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3240,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3241,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3242,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3243,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3244,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3245,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3246,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3247,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3248,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3249,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3250,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3252,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3253,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3255,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3256,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3257,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3258,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3259,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3261,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3262,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3264,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3265,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3266,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3267,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3268,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3269,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3270,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3271,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3272,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3273,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3274,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3275,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3276,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3277,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3279,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3280,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3282,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3283,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3284,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3285,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3286,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3288,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3289,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3290,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3292,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3293,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3295,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3296,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3297,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3298,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3300,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3301,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3302,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3304,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3305,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3307,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3308,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3309,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3310,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3313,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3314,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3315,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3316,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3317,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3318,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3319,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3320,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3321,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3323,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3324,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3325,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3327,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3328,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3329,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3330,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3331,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3333,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3334,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3336,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3337,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3338,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3339,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3340,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3341,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3342,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3343,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3344,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3345,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3346,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3348,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3349,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3350,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3351,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3353,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3354,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3355,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3356,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3357,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3358,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3360,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3361,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3364,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3366,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3368,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3369,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3371,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3372,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3373,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3374,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3375,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3376,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3377,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3378,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3379,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3380,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3381,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3384,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3385,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3387,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3389,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3390,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3391,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3392,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3393,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3395,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3396,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3397,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3399,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3400,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3401,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3402,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3403,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3404,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3405,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3406,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3407,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3410,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3411,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3413,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3414,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3415,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3416,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3417,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3418,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3419,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3420,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3421,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3422,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3423,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3424,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3425,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3426,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3427,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3429,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3430,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3431,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3433,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3434,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3435,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3436,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3437,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3438,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3439,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3442,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3443,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3444,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3446,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3447,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3448,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3450,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3451,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3452,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3453,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3454,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3455,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3456,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3457,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3458,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3459,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3461,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3462,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3465,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3466,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3468,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3470,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3471,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3473,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3474,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3475,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3476,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3478,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3479,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3481,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3482,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3483,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3485,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3486,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3487,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3488,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3489,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3491,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3492,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3493,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3495,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3496,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3497,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3498,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3500,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3501,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3502,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3504,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3505,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3506,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3507,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3508,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3510,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3511,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3512,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5430,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5437,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5452,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5456,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5457,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5462,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5468,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5477,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5501,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5505,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5507,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5529,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5530,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5534,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5538,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5564,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5566,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5575,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5580,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5618,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5625,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5627,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5669,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5672,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5677,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5680,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5684,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5687,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5692,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5694,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5697,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5700,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5705,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5707,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5711,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5714,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5719,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5722,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5727,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5729,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5732,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5735,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5741,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5743,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5747,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5750,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5755,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5759,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5762,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5766,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5770,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5776,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5778,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8064,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8072,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8078,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8085,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N16704;
INVX3 DFT_compute_cynw_cm_float_mul_E8_M23_2_I0 (.Y(bdw_enable), .A(astall));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1425), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I2 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1429), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I3 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1425), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1429));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I4 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1449), .A(b_exp[0]), .B(b_exp[1]));
AND4XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I5 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1451), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I6 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8072), .A(b_exp[7]), .B(b_exp[6]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1451));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I7 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1449), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8072));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I8 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1485), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I9 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1489), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1485));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I10 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1472), .A(b_man[10]), .B(b_man[9]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I11 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1491), .A(b_man[6]), .B(b_man[5]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I12 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1480), .A(b_man[8]), .B(b_man[7]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I13 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1500), .A(b_man[4]), .B(b_man[3]));
NAND4XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I14 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1483), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1472), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1491), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1480), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1500));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I15 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1494), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I16 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1504), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I17 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1489), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1483), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1494), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1504));
NOR2BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I18 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I19 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20));
NOR3BXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I20 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N269), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I21 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1314), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I22 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1318), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I23 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1314), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1318));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I24 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1338), .A(a_exp[0]), .B(a_exp[1]));
AND4XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I25 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1340), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I26 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8064), .A(a_exp[7]), .B(a_exp[6]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1340));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I27 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1338), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8064));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I28 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1374), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I29 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1378), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1374));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I30 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1361), .A(a_man[10]), .B(a_man[9]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I31 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1380), .A(a_man[6]), .B(a_man[5]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I32 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1369), .A(a_man[8]), .B(a_man[7]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I33 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1389), .A(a_man[4]), .B(a_man[3]));
NAND4XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I34 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1372), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1361), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1380), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1369), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1389));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I35 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1383), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I36 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1393), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I37 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1378), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1372), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1383), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1393));
NOR2BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I38 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I39 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19));
NOR3BXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I40 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N270), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I41 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N269), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N270));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I42 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N268), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I43 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N267), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I44 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N268), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N267));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I45 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5452), .A(a_exp[7]));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I46 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5456), .A(b_exp[0]), .B(a_exp[0]));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I47 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5449), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]), .A(b_exp[1]), .B(a_exp[1]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5456));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I48 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5468), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]), .A(b_exp[2]), .B(a_exp[2]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5449));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I49 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5480), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]), .A(b_exp[3]), .B(a_exp[3]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5468));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I50 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5462), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]), .A(b_exp[4]), .B(a_exp[4]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I51 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5477), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]), .A(b_exp[5]), .B(a_exp[5]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5462));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I52 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5457), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]), .A(b_exp[6]), .B(a_exp[6]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I53 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5452), .B(b_exp[7]), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5457));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I54 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]), .A(a_exp[7]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472));
NOR3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I55 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5564), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]));
OR3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I56 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5529), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I57 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5538), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I58 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0]), .A(b_exp[0]), .B(a_exp[0]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I59 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5530), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I60 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8]), .A(a_exp[7]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472));
NOR4BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I61 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5534), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5530), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]));
NAND3BXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I62 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N273), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5529), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5538), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5534));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I63 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5566), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5564), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N273));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I64 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5430), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I65 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5437), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I66 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N272), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5437), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24));
OAI2BB1X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I67 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30), .A0N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5430), .A1N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N272));
NAND3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I68 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5507), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]));
AND4XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I69 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5505), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I70 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5501), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5505));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I71 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N276), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5507), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5501));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I72 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8078), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N276));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I73 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__41), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8078), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I74 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__41));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I75 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__60), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5566), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37));
NAND3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I76 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5580), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]));
NAND4XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I77 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5575), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I78 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N274), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5580), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5575));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I79 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8085), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N274));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I80 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__42), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8085), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I81 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__42));
NOR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I82 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__61), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I83 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .A(a_man[22]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I84 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1991), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I85 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905), .A(b_man[22]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I86 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3087), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I87 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3094), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I88 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480), .A(b_man[21]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I89 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2231), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I90 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .A(a_man[21]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I91 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2250), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I92 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2066), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1641), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3094), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2231), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2250));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I93 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1991), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3087), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2066));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I94 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3357), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I95 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049), .A(b_man[20]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I96 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3341), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I97 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2240), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I98 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3426), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2994), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3357), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3341), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2240));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I99 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .A(a_man[20]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I100 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1657), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I101 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623), .A(b_man[19]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I102 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2486), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I103 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2502), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I104 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1962), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3495), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1657), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2486), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2502));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I105 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2512), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I106 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2319), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1887), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1962), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2512), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2994));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I107 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1641), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3426), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2319));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I108 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I109 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3349), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I110 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .A(a_man[19]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I111 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2769), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I112 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1911), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I113 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157), .A(b_man[18]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I114 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1628), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I115 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2761), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I116 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1610), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3141), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1911), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1628), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2761));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I117 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2820), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2390), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3349), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2769), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1610));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I118 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1647), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I119 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .A(a_man[18]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I120 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3026), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I121 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2494), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I122 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2466), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2030), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1647), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3026), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2494));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I123 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1716), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3245), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3495), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2466), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2390));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I124 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1887), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2820), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1716));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I125 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I126 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .A(a_man[17]));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I127 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2436), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I128 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301), .A(b_man[16]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I129 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1878), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I130 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3277), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I131 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2253), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1824), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2436), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1878), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3277));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I132 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1638), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I133 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2163), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I134 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .A(a_man[16]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I135 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1587), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I136 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3010), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I137 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3107), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2683), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2163), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1587), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3010));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I138 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2108), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1684), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2253), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1638), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3107));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I139 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1903), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I140 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3286), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I141 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2751), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I142 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3215), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2788), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1903), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3286), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2751));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I143 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2170), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I144 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729), .A(b_man[17]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I145 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2736), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I146 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3018), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I147 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2362), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1929), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2170), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2736), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3018));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I148 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2743), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I149 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1893), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I150 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2690), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I151 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871), .A(b_man[15]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I152 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2983), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I153 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1574), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I154 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3255), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2829), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2690), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2983), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1574));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I155 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2003), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1576), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2743), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1893), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3255));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I156 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2964), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2540), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2788), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1929), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2003));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I157 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2212), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1781), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2108), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2030), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2964));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I158 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3319), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2890), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3215), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2362), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3141));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I159 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2212), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3319), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3245));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I160 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I161 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2999), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I162 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2154), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I163 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1885), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I164 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3003), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2579), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2999), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2154), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1885));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I165 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2426), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I166 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .A(a_man[15]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I167 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1843), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I168 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3270), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I169 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2149), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1725), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2426), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1843), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3270));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I170 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2859), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2434), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3003), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2149), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1824));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I171 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2681), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I172 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .A(a_man[14]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I173 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2102), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I174 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1564), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I175 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2293), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1866), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2681), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2102), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1564));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I176 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2949), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I177 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412), .A(b_man[14]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I178 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2128), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I179 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1835), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I180 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3404), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2972), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2949), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2128), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1835));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I181 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3262), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I182 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2416), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I183 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2145), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I184 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3150), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2722), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3262), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2416), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2145));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I185 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1896), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3435), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2293), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3404), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3150));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I186 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1750), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3288), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1896), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2683), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1576));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I187 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1858), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3395), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1684), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2859), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1750));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I188 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1858), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2890), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1781));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I189 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I190 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I191 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2756), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2328), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1725), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2829), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2579));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I192 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1556), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I193 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2672), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I194 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2407), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I195 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2444), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2010), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1556), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2672), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2407));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I196 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2898), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2475), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2972), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2444), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1866));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I197 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3209), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I198 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978), .A(b_man[13]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I199 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3235), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I200 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2092), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I201 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2691), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2263), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3209), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3235), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2092));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I202 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2991), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I203 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2941), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I204 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .A(a_man[13]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I205 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2365), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I206 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1826), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I207 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1585), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3117), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2941), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2365), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1826));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I208 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2039), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1619), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2691), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2991), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1585));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I209 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1650), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3181), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2898), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2039), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3435));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I210 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2610), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2179), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2434), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2756), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1650));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I211 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2610), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2540), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3395));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I212 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I213 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2137), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I214 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3253), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I215 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3466), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I216 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556), .A(b_man[12]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I217 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2380), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I218 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2357), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I219 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3083), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2659), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3466), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2380), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2357));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I220 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3296), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2868), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2137), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3253), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3083));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I221 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1816), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I222 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2928), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I223 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2664), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I224 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2839), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2411), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1816), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2928), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2664));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I225 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3199), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I226 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .A(a_man[12]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I227 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2620), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I228 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2083), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I229 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1979), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1553), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3199), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2620), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2083));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I230 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2397), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I231 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3511), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I232 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3244), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I233 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1734), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3264), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2397), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3511), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3244));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I234 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2188), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1760), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2839), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1979), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1734));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I235 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1791), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3327), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3296), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2722), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2188));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I236 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3043), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2618), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3117), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2263), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2010));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I237 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2650), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2221), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1619), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3043), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2475));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I238 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2505), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2075), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2328), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1791), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2650));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I239 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2505), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3288), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2179));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I240 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I241 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I242 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3457), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I243 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .A(a_man[11]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I244 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2880), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I245 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2345), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I246 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3479), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3054), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3457), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2880), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2345));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I247 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1762), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I248 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122), .A(b_man[11]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I249 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3483), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I250 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2613), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I251 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2626), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2197), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3483), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2613));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I252 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2074), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I253 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3192), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I254 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2920), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I255 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2379), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1950), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2074), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3192), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2920));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I256 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2588), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2160), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3479), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2626), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2379));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I257 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2658), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I258 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1809), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I259 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3502), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I260 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3232), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2807), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1809), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3502));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I261 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3443), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3013), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2659), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3232), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1553));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I262 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1939), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3472), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2868), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2588), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3443));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I263 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2018), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I264 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702), .A(b_man[10]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I265 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2629), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I266 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2873), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I267 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3273), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2846), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2018), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2629), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2873));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I268 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2388), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I269 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1755), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I270 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .A(a_man[10]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I271 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3139), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I272 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2604), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I273 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2166), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1739), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1755), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3139), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2604));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I274 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2124), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1704), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3273), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2388), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2166));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I275 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2336), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1905), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3264), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2411), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2124));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I276 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2797), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2370), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2336), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1760), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2618));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I277 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3505), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3075), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3327), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1939), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2797));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I278 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3505), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3181), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2075));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I279 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I280 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1875), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3413), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1950), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3054), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2807));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I281 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2914), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I282 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2065), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I283 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1801), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I284 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1914), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3450), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2914), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2065), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1801));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I285 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2338), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I286 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3449), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I287 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3183), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I288 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3020), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2597), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2338), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3449), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3183));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I289 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2982), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2559), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1914), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3020), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2197));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I290 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3193), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2765), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1875), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2982), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2160));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I291 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2595), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I292 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1747), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I293 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3442), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I294 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2814), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2387), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2595), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1747), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3442));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I295 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2012), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I296 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .A(a_man[9]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I297 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3401), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I298 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2861), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I299 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1958), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3487), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2012), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3401), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2861));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I300 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3174), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I301 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2326), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I302 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2057), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I303 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1712), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3241), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3174), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2326), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2057));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I304 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1667), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3200), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2814), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1958), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1712));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I305 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3492), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I306 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2648), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I307 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2283), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I308 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228), .A(b_man[9]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I309 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1769), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I310 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3128), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I311 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3063), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2635), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2283), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1769), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3128));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I312 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2772), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2343), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3492), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2648), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3063));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I313 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1787), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I314 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2904), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I315 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2638), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I316 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2566), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2131), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1787), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2904), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2638));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I317 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2525), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2094), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2846), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2566), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1739));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I318 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2731), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2304), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1667), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2772), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2525));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I319 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2084), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1660), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2731), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3013), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1905));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I320 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1694), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3223), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3472), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3193), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2084));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I321 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1694), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2221), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3075));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I322 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I323 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I324 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2274), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I325 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .A(a_man[8]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I326 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1701), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I327 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3119), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I328 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2854), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2428), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2274), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1701), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3119));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I329 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2547), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I330 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806), .A(b_man[8]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I331 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2879), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I332 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3391), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I333 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1998), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1569), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2547), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2879), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3391));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I334 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2853), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I335 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2005), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I336 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1741), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I337 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1745), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3282), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2853), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2005), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1741));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I338 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3420), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2990), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2854), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1998), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1745));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I339 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3377), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2947), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3450), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2597), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3420));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I340 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1627), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3161), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3377), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1704), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2559));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I341 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2048), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I342 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3167), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I343 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2896), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I344 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3459), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3028), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2048), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3167), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2896));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I345 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3434), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I346 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2590), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I347 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2318), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I348 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2605), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2174), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3434), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2590), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2318));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I349 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2314), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1880), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3459), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2605), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2635));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I350 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3168), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2738), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2387), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3487), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3241));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I351 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2270), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1844), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2314), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2343), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3168));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I352 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2483), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2051), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2270), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3413), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2304));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I353 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2939), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2517), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2765), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1627), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2483));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I354 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2939), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2370), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3223));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I355 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I356 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2803), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I357 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375), .A(b_man[7]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I358 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2020), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I359 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1692), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I360 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2034), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1611), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2803), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2020), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1692));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I361 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1779), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I362 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2537), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I363 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .A(a_man[7]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I364 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1954), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I365 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3379), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I366 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2894), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2469), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2537), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1954), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3379));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I367 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2355), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1924), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2034), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1779), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2894));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I368 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1733), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I369 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2844), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I370 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2581), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I371 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2642), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2215), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1733), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2844), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2581));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I372 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3111), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I373 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2265), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I374 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1997), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I375 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1785), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3323), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3111), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2265), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1997));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I376 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2309), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I377 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3425), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I378 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3159), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I379 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3500), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3069), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2309), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3425), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3159));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I380 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3211), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2782), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2642), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1785), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3500));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I381 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2060), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1636), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2355), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2131), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3211));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I382 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3126), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2699), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2094), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3200), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2060));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I383 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2103), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1676), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2428), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1569), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3282));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I384 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2888), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I385 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2038), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I386 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3059), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I387 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948), .A(b_man[6]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I388 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3127), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I389 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1947), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I390 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3185), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2760), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3059), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3127), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1947));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I391 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2395), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1965), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2888), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2038), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3185));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I392 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2957), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2535), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3028), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2174), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2395));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I393 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2916), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2490), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2990), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2103), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2957));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I394 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2016), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1593), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2916), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2947), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1844));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I395 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3336), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2909), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3161), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3126), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2016));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I396 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3336), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1660), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2517));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I397 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I398 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I399 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I400 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3147), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I401 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2300), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I402 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2029), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I403 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1580), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3109), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3147), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2300), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2029));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I404 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2572), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I405 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1723), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I406 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3419), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I407 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2686), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2257), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2572), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1723), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3419));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I408 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2143), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1719), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1580), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2686), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1611));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I409 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3372), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I410 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2527), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I411 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2255), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I412 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2934), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2507), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3372), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2527), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2255));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I413 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2794), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I414 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .A(a_man[6]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I415 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2211), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I416 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1681), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I417 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2079), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1654), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2794), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2211), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1681));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I418 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1987), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I419 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3101), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I420 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2838), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I421 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1828), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3366), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1987), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3101), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2838));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I422 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3248), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2823), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2934), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2079), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1828));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I423 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2997), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2574), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3323), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2469), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2215));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I424 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1853), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3389), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2143), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3248), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2997));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I425 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1810), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3346), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2738), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1880), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1853));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I426 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3049), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I427 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .A(a_man[5]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I428 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2474), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I429 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1936), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I430 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2373), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1944), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3049), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2474), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1936));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I431 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3318), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I432 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477), .A(b_man[5]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I433 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2273), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I434 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2205), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I435 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3474), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3046), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3318), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2273), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2205));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I436 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1671), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I437 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2784), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I438 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2519), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I439 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3226), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2800), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1671), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2784), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2519));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I440 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2438), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2007), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2373), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3474), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3226));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I441 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2828), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I442 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1981), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I443 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1715), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I444 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2975), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2553), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2828), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1981), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1715));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I445 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2246), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I446 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3364), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I447 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3092), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I448 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2118), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1698), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2246), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3364), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3092));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I449 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3411), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I450 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2565), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I451 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2291), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I452 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1869), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3407), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3411), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2565), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2291));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I453 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3292), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2863), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2975), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2118), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1869));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I454 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1889), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3429), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2438), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3069), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3292));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I455 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2708), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2279), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2782), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1924), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1889));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I456 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2667), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2238), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2708), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1636), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2490));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I457 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2876), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2451), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2699), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1810), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2667));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I458 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2876), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2051), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2909));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I459 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I460 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2183), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1753), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1654), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2760), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2507));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I461 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2750), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2322), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2183), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1965), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2823));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I462 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1603), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3137), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2535), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1676), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2750));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I463 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3036), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2615), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2257), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3366), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3109));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I464 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1644), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3175), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1719), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3036), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2574));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I465 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2461), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2026), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1644), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3389), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2279));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I466 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1559), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3090), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3346), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1603), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2461));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I467 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1559), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1593), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2451));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I468 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I469 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I470 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3330), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2903), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1698), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2800), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2553));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I471 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2792), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2363), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2007), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3330), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2863));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I472 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2509), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I473 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1662), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I474 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3354), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I475 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1555), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3086), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2509), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1662), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3354));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I476 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1926), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I477 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3041), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I478 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2774), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I479 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2661), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2233), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1926), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3041), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2774));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I480 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3082), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I481 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2236), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I482 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1973), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I483 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2414), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1983), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3082), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2236), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1973));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I484 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1622), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3155), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1555), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2661), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2414));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I485 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1618), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I486 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050), .A(b_man[4]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I487 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3381), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I488 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2465), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I489 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2913), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2485), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1618), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3381), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2465));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I490 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3138), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I491 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3310), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I492 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .A(a_man[4]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I493 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2730), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I494 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2193), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I495 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1807), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3340), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3310), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2730), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2193));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I496 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2725), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2298), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2913), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3138), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1807));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I497 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1708), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I498 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2819), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I499 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2555), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I500 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3267), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2840), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1708), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2819), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2555));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I501 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2478), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2042), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3046), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3267), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1944));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I502 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1934), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3468), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1622), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2725), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2478));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I503 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2498), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2069), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2792), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1934), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3429));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I504 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2282), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I505 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3403), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I506 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1874), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I507 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623), .A(b_man[3]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I508 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2526), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I509 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2721), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I510 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3453), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3022), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1874), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2526), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2721));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I511 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2162), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1736), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2282), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3403), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3453));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I512 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2185), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I513 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3302), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I514 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3031), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I515 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3203), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2775), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2185), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3302), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3031));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I516 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1609), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I517 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .A(a_man[3]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I518 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2989), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I519 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2457), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I520 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2348), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1918), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1609), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2989), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2457));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I521 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2767), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I522 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1916), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I523 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1652), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I524 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2097), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1669), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2767), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1916), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1652));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I525 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3016), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2591), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3203), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2348), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2097));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I526 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2224), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1796), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2162), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3407), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3016));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I527 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1686), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3219), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1753), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2224), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2615));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I528 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3356), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2924), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1686), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2322), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3175));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I529 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3315), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2885), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3137), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2498), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3356));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I530 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3315), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2238), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3090));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I531 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I532 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1664), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3195), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1983), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3086), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2840));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I533 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1974), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3510), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1664), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2042));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I534 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2768), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2340), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3340), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2485), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2233));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I535 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1964), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I536 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3073), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I537 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2813), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I538 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1847), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3380), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1964), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3073), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2813));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I539 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3345), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I540 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2500), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I541 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2229), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I542 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2952), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2529), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3345), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2500), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2229));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I543 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2546), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I544 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1700), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I545 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3393), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I546 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2702), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2272), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2546), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1700), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3393));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I547 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1908), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3446), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1847), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2952), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I548 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3078), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2653), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2768), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1908), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2298));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I549 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2545), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2111), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1974), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3078), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2363));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I550 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1643), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I551 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2758), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I552 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2492), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I553 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2637), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2208), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1643), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2758), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2492));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I554 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3023), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I555 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2176), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I556 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1909), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I557 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1780), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3317), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3023), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2176), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1909));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I558 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2220), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I559 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3338), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I560 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3065), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I561 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3491), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3064), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2220), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3338), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3065));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I562 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2454), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2019), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2637), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1780), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3491));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I563 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1865), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I564 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .A(a_man[2]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I565 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3247), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I566 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2711), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I567 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2028), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1606), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1865), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3247), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2711));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I568 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2134), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I569 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196), .A(b_man[2]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I570 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1670), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I571 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2981), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I572 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3140), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2710), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2134), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1670), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2981));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I573 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2449), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I574 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1602), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I575 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3293), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I576 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2887), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2463), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2449), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1602), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3293));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I577 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1597), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3130), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2028), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3140), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2887));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I578 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2518), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2087), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2454), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1597), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1736));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I579 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2833), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2404), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2518), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2903), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1796));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I580 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3399), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2965), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3468), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3219));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I581 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2247), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1818), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2069), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2545), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3399));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I582 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2247), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2026), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2885));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I583 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I584 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I585 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I586 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765), .A(b_man[1]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I587 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2776), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I588 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2393), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I589 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1969), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3501), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2776), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2393));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I590 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2536), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I591 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3239), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I592 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .A(a_man[1]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I593 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3508), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I594 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2123), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I595 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2824), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2398), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3239), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3508), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2123));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I596 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3243), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2816), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1969), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2536), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2824));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I597 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3057), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2628), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2272), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3380), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3243));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I598 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2200), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1771), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1669), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2775), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2529));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I599 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2267), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1838), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3057), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2200), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2340));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I600 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2805), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I601 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1957), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I602 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1691), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I603 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2389), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1960), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2805), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1957), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1691));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I604 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3309), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2878), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3022), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2389), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1918));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I605 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3374), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2944), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2591), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3309), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3446));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I606 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1728), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3257), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2267), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3374), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2653));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I607 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2210), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I608 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3329), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I609 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3058), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I610 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3178), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2752), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2210), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3329), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3058));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I611 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1634), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I612 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2748), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I613 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2482), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I614 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2325), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1892), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1634), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2748), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2482));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I615 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2796), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I616 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1946), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I617 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1680), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I618 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2071), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1646), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2796), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1946), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1680));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I619 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2993), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2569), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3178), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2325), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2071));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I620 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2442), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I621 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1591), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I622 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3283), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I623 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2576), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2144), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2442), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1591), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3283));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I624 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1856), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I625 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2971), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I626 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2704), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I627 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1722), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3252), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1856), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2971), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2704));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I628 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3015), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I629 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2168), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I630 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1900), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I631 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3430), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3000), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3015), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2168), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1900));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I632 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2136), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1714), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2576), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1722), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3430));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I633 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1884), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3422), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1606), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2710), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2463));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I634 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1953), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3482), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2993), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2136), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1884));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I635 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2742), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2317), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2208), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3317), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3064));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I636 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2811), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2382), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3130), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2742), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2019));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I637 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3118), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2695), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1953), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3195), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2811));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I638 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2582), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2153), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3510), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3118), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2404));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I639 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2286), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1862), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2111), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1728), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2582));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I640 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2286), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2924), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1818));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I641 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I642 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303), .A(b_man[0]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I643 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1915), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I644 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2652), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I645 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2763), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2334), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1915), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2652));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I646 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3498), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I647 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .A(a_man[0]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I648 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1806), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I649 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2386), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I650 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1656), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3188), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3498), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1806), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2386));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I651 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2927), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2501), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3501), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2763), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1656));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I652 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2696), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I653 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1849), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I654 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1582), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I655 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3368), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2937), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2696), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1849), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1582));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I656 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2114), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I657 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3231), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I658 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2963), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I659 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2511), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2082), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3231), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2963));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I660 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3275), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I661 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2431), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I662 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2161), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I663 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2260), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1830), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3275), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2431), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2161));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I664 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1821), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3358), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3368), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2511), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2260));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I665 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1639), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3171), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2927), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1960), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1821));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I666 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1707), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3234), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2878), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1639), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1771));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I667 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2014), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1590), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2944), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2087), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1707));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I668 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2473), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I669 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1626), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I670 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3321), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I671 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2008), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1583), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2473), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1626), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3321));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I672 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1891), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I673 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3005), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I674 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2740), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I675 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3113), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2689), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1891), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3005), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2740));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I676 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3048), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I677 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2204), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I678 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1935), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I679 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2865), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2441), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3048), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2204), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1935));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I680 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2679), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2249), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2008), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3113), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2865));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I681 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1572), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3103), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3252), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2398), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2144));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I682 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2493), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2061), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2816), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2679), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1572));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I683 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2430), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1999), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1892), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3000), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2752));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I684 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3348), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2919), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1714), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2430), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2569));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I685 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2563), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2127), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2493), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2628), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3348));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I686 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2872), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2445), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1838), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2563), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2695));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I687 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3438), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3007), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3257), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2014), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2872));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I688 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3438), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2965), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1862));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I689 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I690 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I691 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I692 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I693 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1592), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I694 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2786), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I695 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1757), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3295), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1592), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2786), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2334));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I696 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2106), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I697 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3222), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I698 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2953), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I699 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2194), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1764), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2106), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3222), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2953));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I700 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3486), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I701 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2641), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I702 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2378), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I703 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3304), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2874), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3486), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2641), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2378));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I704 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2687), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I705 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1841), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I706 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1571), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I707 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3047), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2624), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2687), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1841), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1571));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I708 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2616), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2186), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2194), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3304), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3047));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I709 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3284), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2856), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1757), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1646), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2616));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I710 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2242), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1813), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3422), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3284), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2317));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I711 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3416), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2985), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2382), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3482), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2242));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I712 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1882), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I713 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2996), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I714 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2733), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I715 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2804), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2374), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1882), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2996), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2733));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I716 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3268), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I717 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2421), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I718 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2151), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I719 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1949), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3476), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3268), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2421), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2151));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I720 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2464), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I721 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1617), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I722 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3314), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I723 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1699), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3229), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2464), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1617), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3314));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I724 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3470), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3039), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2804), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1949), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1699));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I725 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3040), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I726 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2195), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I727 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1925), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I728 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2557), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2121), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3040), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2195), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1925));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I729 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2367), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1938), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3188), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2557), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2082));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I730 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2177), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1748), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2501), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3470), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2367));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I731 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3220), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2795), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1830), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2937), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2689));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I732 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3030), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2606), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3358), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3220), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2249));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I733 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3093), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2668), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3171), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2177), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3030));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I734 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2308), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1877), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3234), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3093), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2127));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I735 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1761), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3300), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1590), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3416), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2308));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I736 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1761), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2153), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3007));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I737 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I738 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3121), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I739 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2053), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I740 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2901), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I741 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2129), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1709), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2053), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2901));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I742 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2634), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I743 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1784), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I744 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3478), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I745 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2986), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2564), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2634), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1784), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3478));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I746 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3410), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2976), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3121), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2129), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2986));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I747 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2113), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1690), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2441), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1583), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3410));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I748 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1927), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3461), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3103), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2113), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1999));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I749 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1990), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1563), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2919), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2061), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1927));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I750 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1832), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I751 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2945), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I752 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2678), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I753 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2737), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2310), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1832), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2945), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2678));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I754 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3213), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I755 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2369), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I756 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2098), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I757 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1879), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3418), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3213), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2369), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2098));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I758 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2413), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I759 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1561), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I760 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3259), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I761 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1633), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3166), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2413), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1561), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3259));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I762 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2299), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1872), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2737), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1879), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1633));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I763 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1608), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I764 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2724), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I765 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2456), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I766 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3342), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2915), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1608), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2724), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2456));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I767 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2988), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I768 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2141), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I769 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1873), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I770 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2488), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2056), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2988), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2141), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1873));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I771 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2187), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I772 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3301), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I773 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3164), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I774 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2041), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I775 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1566), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3098), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3164), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2041));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I776 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2235), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1808), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2187), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3301), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1566));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I777 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3158), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2728), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3342), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2488), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2235));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I778 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2968), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2548), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3295), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2299), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3158));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I779 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2047), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1624), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1764), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2874), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2624));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I780 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1863), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3402), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2186), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2047), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3039));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I781 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2785), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2358), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2856), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2968), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1863));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I782 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2849), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2422), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1813), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2785), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2668));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I783 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3165), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2735), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2985), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1990), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2849));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I784 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3165), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2445), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3300));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I785 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I786 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I787 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I788 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2906), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2481), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2374), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3476), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3229));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I789 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2719), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2290), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2906), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2795));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I790 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1679), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3212), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2606), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1748), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2719));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I791 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1776), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I792 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2893), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I793 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2625), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I794 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2425), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1993), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1776), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2893), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2625));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I795 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2361), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I796 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3471), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I797 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3206), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I798 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3276), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2852), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2361), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3471), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3206));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I799 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3089), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2663), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2425), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1709), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3276));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I800 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1554), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I801 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2669), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I802 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2402), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I803 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3025), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2600), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1554), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2669), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2402));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I804 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2936), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I805 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2089), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I806 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1822), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I807 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2172), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1744), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2936), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2089), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1822));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I808 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2133), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I809 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3250), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I810 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2980), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I811 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1919), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3456), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2133), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3250), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2980));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I812 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1984), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1557), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3025), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2172), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1919));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I813 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1800), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3333), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3089), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2121), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1984));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I814 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2714), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I815 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1864), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I816 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1601), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I817 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2779), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2353), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2714), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1864), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1601));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I818 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2843), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2415), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2564), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2779), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3418));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I819 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2657), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2227), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2843), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2976), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1872));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I820 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1614), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3149), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1690), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1800), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2657));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I821 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2306), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I822 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3153), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I823 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1859), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3396), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2306), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3153));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I824 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2448), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I825 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1674), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3205), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1859), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2448), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3098));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I826 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2592), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2164), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1674), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2915), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1808));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I827 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1738), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3269), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3166), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2310), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2056));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I828 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3512), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3081), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2592), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1738), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2728));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I829 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2472), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2037), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3512), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2548), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3402));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I830 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2538), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2105), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3461), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1614), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2472));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I831 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1742), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3274), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1563), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1679), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2538));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I832 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1742), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1877), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2735));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I833 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I834 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3238), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I835 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2392), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I836 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2126), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I837 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2209), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1782), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3238), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2392), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2126));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I838 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2662), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I839 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1812), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I840 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3507), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I841 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3320), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2889), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2662), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1812), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3507));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I842 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1855), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I843 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2970), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I844 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2703), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I845 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3067), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2640), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1855), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2970), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2703));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I846 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3385), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2956), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2209), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3320), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3067));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I847 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3462), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I848 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2617), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I849 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2350), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I850 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1607), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3142), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3462), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2617), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2350));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I851 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2884), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I852 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2032), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I853 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1767), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I854 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2713), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2284), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2884), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2032), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1767));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I855 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2080), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I856 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3197), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I857 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2926), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I858 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2467), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2031), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2080), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3197), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2926));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I859 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2531), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2101), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1607), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2713), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2467));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I860 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2277), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1848), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2852), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1993), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1744));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I861 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3448), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3017), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3385), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2531), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2277));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I862 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2406), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1977), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2481), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1624), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3448));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I863 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3325), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2895), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2290), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2406), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3149));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I864 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3392), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2959), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3212), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2358), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3325));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I865 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3392), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2422), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3274));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I866 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I867 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I868 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3131), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2707), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3456), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2600), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2353));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I869 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2342), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1910), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2663), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3131), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1557));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I870 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3261), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2836), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3333), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2342), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2227));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I871 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3189), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I872 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2341), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I873 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2070), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I874 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1651), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3182), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3189), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2341), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2070));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I875 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2608), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I876 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1759), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I877 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3454), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I878 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2754), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2329), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2608), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1759), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3454));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I879 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1805), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I880 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2918), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I881 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2655), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I882 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2506), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2073), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1805), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2918), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2655));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I883 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2818), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2391), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1651), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2754), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2506));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I884 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3415), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I885 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2296), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I886 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3004), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2580), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3415), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2296));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I887 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2024), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I888 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3144), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I889 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2875), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I890 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1897), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3433), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2024), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3144), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2875));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I891 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1963), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3493), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3396), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3004), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1897));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I892 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2023), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1600), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2818), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1963), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3205));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I893 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3196), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2770), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3269), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2415), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2023));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I894 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2156), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1731), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3196), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1977));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I895 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2216), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1788), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2037), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3261), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2156));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I896 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2216), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2105), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2959));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I897 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I898 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2962), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I899 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2117), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I900 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2562), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I901 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3406), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I902 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3042), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2619), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2562), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3406));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I903 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2254), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1825), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2962), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2117), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3042));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I904 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2385), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I905 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3497), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I906 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3230), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I907 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3360), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2931), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2385), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3497), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3230));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I908 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1717), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3246), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2254), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3360), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2284));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I909 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2883), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2455), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2101), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1717), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2956));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I910 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2091), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1665), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2883), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2164), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3017));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I911 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3135), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I912 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2288), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I913 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2015), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I914 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1940), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3473), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3135), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2288), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2015));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I915 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1752), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I916 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2867), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I917 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2601), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I918 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2798), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2368), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1752), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2867), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2601));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I919 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3108), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2680), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1940), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2580), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2798));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I920 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3424), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2995), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2640), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1782), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3108));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I921 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2571), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2138), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2031), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3142), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2889));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I922 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1773), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3313), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3424), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2571), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1848));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I923 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2910), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I924 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2062), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I925 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1793), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I926 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2550), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2116), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2910), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2062), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1793));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I927 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2333), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I928 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3447), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I929 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3179), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I930 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1693), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3224), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2333), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3447), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3179));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I931 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3489), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I932 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2644), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I933 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2377), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I934 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3405), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2969), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3489), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2644), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2377));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I935 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2000), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1577), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2550), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1693), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3405));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I936 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2860), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2435), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2329), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3433), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3182));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I937 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2320), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1888), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3493), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2000), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2860));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I938 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2632), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2203), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2320), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2707), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1600));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I939 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2946), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2521), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1910), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1773), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2632));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I940 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3009), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2585), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2836), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2091), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2946));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I941 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3009), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2895), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1788));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I942 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I943 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I944 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I945 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2749), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I946 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1705), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I947 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2551), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I948 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1980), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1551), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1705), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2551));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I949 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3221), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I950 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2292), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1867), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1980), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3221), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2619));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I951 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1751), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3285), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2931), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2073), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2292));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I952 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3173), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2744), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1751), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2391), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3246));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I953 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2857), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I954 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2009), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I955 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1743), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I956 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1735), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3265), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2857), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2009), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1743));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I957 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2278), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I958 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3397), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I959 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3124), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I960 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2837), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2412), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2278), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3397), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3124));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I961 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3439), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I962 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2593), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I963 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2324), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I964 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2589), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2157), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3439), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2593), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2324));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I965 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3151), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2723), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1735), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2837), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2589));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I966 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2633), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I967 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1783), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I968 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3481), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I969 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2337), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1906), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2633), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1783), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3481));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I970 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2055), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I971 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3170), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I972 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2900), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I973 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3444), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3014), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2055), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3170), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2900));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I974 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2040), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1616), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2337), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3444), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3473));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I975 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2611), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2180), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3151), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1825), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2040));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I976 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2064), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1642), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2611), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2138), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2995));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I977 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3485), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3061), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2455), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3173), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2064));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I978 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1840), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3375), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3485), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2770), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1665));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I979 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1840), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1731), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2585));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I980 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I981 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2897), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2476), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3224), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2368), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2116));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I982 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3465), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3034), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2680), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2897), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1577));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I983 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2810), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I984 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1696), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I985 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1766), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3307), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2810), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1696));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I986 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3387), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I987 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2543), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I988 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2269), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I989 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2627), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2198), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3387), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2543), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2269));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I990 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3191), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2766), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1551), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1766), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2627));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I991 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2586), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I992 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1737), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I993 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3431), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I994 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2376), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1951), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2586), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1737), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3431));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I995 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2001), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I996 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3116), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I997 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2850), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I998 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3480), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3052), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2001), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3116), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2850));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I999 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3163), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1000 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2315), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1001 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2044), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1002 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3233), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2808), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3163), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2315), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2044));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1003 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2085), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1661), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2376), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3480), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3233));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1004 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1792), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3328), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3191), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2969), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2085));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1005 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2360), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1930), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2435), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1792), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3285));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1006 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2922), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2497), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1888), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3465), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2360));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1007 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2383), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1956), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2922), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3313), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2203));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1008 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2383), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2521), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3375));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1009 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1010 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1011 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1775), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1012 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2892), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1013 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1952), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1014 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2799), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1015 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2419), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1986), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1952), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2799));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1016 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2125), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1703), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1775), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2892), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2419));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1017 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2940), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2515), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2412), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2125), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3265));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1018 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2651), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2219), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2940), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1867), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2723));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1019 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1834), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3371), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3014), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2157), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1906));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1020 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3504), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3076), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1616), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1834), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2476));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1021 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3216), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2789), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2180), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2651), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3504));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1022 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1815), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3350), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1642), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2744), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3216));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1023 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1815), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3061), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1956));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1024 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1025 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2305), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1026 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3423), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1027 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3152), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1028 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1912), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3451), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2305), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3423), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3152));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1029 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1730), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1030 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2841), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1031 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2577), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1032 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3021), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2594), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1730), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2841), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2577));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1033 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1876), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3414), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1912), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3021), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2198));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1034 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2534), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1035 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1685), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1036 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3376), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1037 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3271), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2847), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2534), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1685), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3376));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1038 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3105), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1039 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2262), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1040 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1994), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1041 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2167), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1740), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3105), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2262), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1994));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1042 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2979), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2560), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3271), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3307), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2167));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1043 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2732), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2302), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1951), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3052), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2808));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1044 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2692), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2264), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1876), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2979), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2732));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1045 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3055), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1046 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1942), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1047 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1959), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3488), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3055), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1942));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1048 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2036), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1049 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2773), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2344), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1959), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2036), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1986));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1050 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2251), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1051 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3369), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1052 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3096), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1053 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1710), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3242), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2251), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3369), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3096));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1054 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1675), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1055 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2790), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1056 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2523), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1057 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2815), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2384), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1675), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2790), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2523));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1058 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2834), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1059 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1985), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1060 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1721), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1061 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2567), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2132), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2834), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1985), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1721));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1062 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1668), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3198), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1710), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2815), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2567));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1063 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1625), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3162), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1703), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2773), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1668));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1064 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1586), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3115), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1661), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2766), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1625));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1065 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2401), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1972), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3328), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2692), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1586));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1066 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2109), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1683), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1930), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3034), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2401));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1067 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2109), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2497), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3350));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1068 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1589), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1069 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1589));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1070 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2645), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1071 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3417), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1072 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2568), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1073 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2295), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1074 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3421), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2987), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3417), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2568), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2295));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1075 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2522), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2095), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2847), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3421), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1740));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1076 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2199), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1077 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3044), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1078 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2356), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1921), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2199), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3044));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1079 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2780), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1080 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1932), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1081 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1666), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1082 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3208), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2783), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2780), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1932), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1666));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1083 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2311), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1881), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3488), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2356), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3208));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1084 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3378), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2948), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3451), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2594), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2311));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1085 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2484), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2052), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2560), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2522), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3378));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1086 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2443), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2011), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3371), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2515), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2484));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1087 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3256), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2827), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3076), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2219), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2443));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1088 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3256), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2789), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1683));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1089 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1090 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1978), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1091 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3088), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1092 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2825), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1093 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2958), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2533), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1978), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3088), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2825));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1094 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3361), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1095 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2516), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1096 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2243), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1097 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2104), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1677), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3361), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2516), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2243));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1098 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2561), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1099 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1713), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1100 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3308), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1101 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2190), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1102 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1645), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3176), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3308), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2190));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1103 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1852), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3390), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2561), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1713), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1645));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1104 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3169), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2739), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2958), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2104), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1852));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1105 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2058), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1637), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3242), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2384), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2132));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1106 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2271), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1842), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3169), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2344), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2058));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1107 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3337), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2907), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2302), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3414), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2271));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1108 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3297), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2869), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3337), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2264), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3115));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1109 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3297), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1972), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2827));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1110 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1839), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1111 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1579), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1839));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1112 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3122), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2700), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2095), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3198), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2948));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1113 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2228), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1804), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2052), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3162), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3122));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1114 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2228), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2011), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2869));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1115 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N16704), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1116 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2452), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1117 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3298), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1118 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1786), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3324), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2452), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3298));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1119 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2817), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1120 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3100), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2674), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1786), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2817), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3176));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1121 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2460), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2027), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3100), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2533), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3390));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1122 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3080), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1123 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2234), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1124 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1968), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1125 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2248), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1819), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3080), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2234), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1968));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1126 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1604), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3134), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2783), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2248), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1677));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1127 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1811), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3344), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2460), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1604), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2739));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1128 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1922), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1129 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3035), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1130 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2771), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1131 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2499), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2067), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1922), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3035), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2771));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1132 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2503), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1133 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1659), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1134 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3351), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1135 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3353), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2925), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2503), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1659), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3351));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1136 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2709), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2280), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2499), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1921), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3353));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1137 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2917), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2491), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2709), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2987), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1881));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1138 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2017), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1594), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1811), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2917), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1842));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1139 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2017), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2907), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1804));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1140 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1141 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2855), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2429), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2925), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2067), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1819));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1142 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1648), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1143 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2764), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1144 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2495), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1145 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3496), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3070), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1648), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2764), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2495));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1146 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3027), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1147 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2181), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1148 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1913), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1149 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2643), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2213), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3027), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2181), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1913));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1150 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2225), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1151 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3343), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1152 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3071), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1153 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2396), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1966), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2225), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3343), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3071));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1154 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1996), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1570), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3496), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2643), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2396));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1155 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3316), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2886), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2855), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1996), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2280));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1156 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2665), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2239), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3316), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1637), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2491));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1157 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2665), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2700), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1594));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1158 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2459), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1159 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3280), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1160 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2437), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1161 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2165), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1162 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1581), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3110), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3280), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2437), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2165));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1163 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1596), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1164 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2446), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1165 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2793), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2364), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1596), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2446));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1166 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1894), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1167 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3012), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1168 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2745), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1169 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2439), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2004), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1894), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3012), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2745));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1170 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2287), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1860), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1581), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2364), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2439));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1171 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2998), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2575), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1966), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3070), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2287));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1172 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2603), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2175), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2998), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1570), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2429));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1173 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2173), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1174 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3290), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1175 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3019), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1176 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1687), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3217), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2173), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3290), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3019));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1177 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3249), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2821), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3324), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2793), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1687));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1178 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3334), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1179 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2487), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1180 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2701), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1181 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1588), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1182 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2684), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2258), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1588));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1183 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3400), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2966), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3334), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2487), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2684));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1184 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2755), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1185 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1907), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1186 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1640), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1187 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2542), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2112), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2755), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1907), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1640));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1188 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2140), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1720), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3400), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2542), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2213));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1189 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1746), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3279), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2674), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3249), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2140));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1190 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2207), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1774), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1746), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3134), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2027));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1191 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2886), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2603), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1774));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1192 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2207), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3344), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2239));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1193 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450));
OAI2BB1X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1194 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2646), .A0N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062), .A1N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1195 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1845), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1196 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2693), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1197 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3436), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3008), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1845), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2693));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1198 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1631), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1199 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3289), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2864), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3436), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1631), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2258));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1200 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3143), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2717), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2112), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3217), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3289));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1201 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1890), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3427), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3143), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2821), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1720));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1202 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1890), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3279), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2175));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1203 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1204 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3001), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1205 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2158), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1206 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1886), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1207 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3186), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2757), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3001), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2158), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1886));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1208 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2427), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1209 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1578), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1210 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3272), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1211 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2332), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1899), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2427), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1578), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3272));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1212 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2184), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1754), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3186), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2332), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3110));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1213 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2035), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1612), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2184), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2966), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1860));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1214 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2035), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2575), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3427));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1215 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2955), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1216 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2148), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1217 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3266), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1218 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2096), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1219 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2942), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1220 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1620), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3156), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2096), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2942));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1221 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2830), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2405), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2148), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3266), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1620));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1222 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2935), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2508), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1899), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2830), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2757));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1223 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2951), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1224 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1837), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1225 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3079), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2654), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2951), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1837));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1226 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1567), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1227 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2685), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1228 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2417), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1229 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1975), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3506), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1567), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2685), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2417));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1230 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2076), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1655), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3008), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3079), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1975));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1231 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3037), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2612), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2076), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2004), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2864));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1232 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1754), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2935), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2612));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1233 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3037), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2717), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1612));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1234 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323));
OAI2BB1X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1235 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2226), .A0N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931), .A1N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1236 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2675), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1237 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1827), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1238 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1558), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1239 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2479), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2043), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2675), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1827), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1558));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1240 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1729), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3258), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2479), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2654), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3506));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1241 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1655), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1729), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2508));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1242 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2352), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1243 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3201), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1244 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2086), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1245 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2973), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2554), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3201), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2086));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1246 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2409), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1247 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3331), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2899), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2973), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2409), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3156));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1248 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2405), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3331), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3258));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1249 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3455), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1250 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1817), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1251 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2932), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1252 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2666), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1253 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1870), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1817), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2932), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2666));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1254 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2043), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1870), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2899));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1255 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2602), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1256 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2347), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1257 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3194), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1258 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3227), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2347), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3194));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1259 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2077), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1260 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2923), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1261 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3452), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1262 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2339), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
ADDHX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1263 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2371), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3452), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2339));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1264 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2119), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2077), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2923), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2371));
ADDFX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1265 (.CO(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726), .S(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2554), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3227), .CI(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2119));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1266 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1584), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1267 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2851), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294));
AND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1268 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1995), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1269 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1270 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3097), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945));
OR4X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1271 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2244), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1272 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2673), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1273 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2631), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3097), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2244), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2673));
OAI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1274 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2130), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1995), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2631), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1275 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2424), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1276 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1632), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2851), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2130), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2424));
OAI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1277 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2842), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1584), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1632), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1278 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2171), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1279 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2090), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2602), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2842), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2171));
OAI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1280 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3051), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3455), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2090), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1281 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1920), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1282 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2046), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2352), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3051), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1920));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1283 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2778), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1284 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1673), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1285 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1799), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2778), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1673));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1286 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2514), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2226), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2046), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1799));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1287 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2532), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1288 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3384), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1289 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2259), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2532), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3384));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1290 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3104), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2259));
AOI31X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1291 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2471), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2955), .A2(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2514), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3104));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1292 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2276), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1293 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3133), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1294 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2217), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2276), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3133));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1295 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2432), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2646), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2471), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2217));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1296 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2022), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1297 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2882), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758));
AO21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1298 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1961), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2022), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2882));
AOI31X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1299 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1883), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2459), .A2(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2432), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1961));
AO22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1300 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2256), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N16704), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1883), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1301 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3373), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1302 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2266), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1303 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3112), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3373), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2266));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1304 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1579), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2256), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3112));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1305 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3120), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1306 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2013), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1307 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3120), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2013));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1308 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1309 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1763), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1310 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2862), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1763));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1311 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2214), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2862));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1312 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2645), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2214));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1313 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1314 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3475), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1315 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3475));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1316 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1317 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3225), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1318 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2614), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3225));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1319 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2614));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1320 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1321 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2974), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1322 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2974));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1323 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1324 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2727), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1325 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2366), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2727));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1326 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1967), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2366));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1327 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2321), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1967));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1328 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2749), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2321));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1329 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1330 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2477), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1331 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2477));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1332 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1333 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2223), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1334 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2110), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2223));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1335 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2110));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1336 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1337 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1976), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1338 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1976));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1339 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1340 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1727), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1341 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1861), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1727));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1342 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1718), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1861));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1343 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3177), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1718));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1344 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3355), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3177));
AOI31X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1345 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251), .A2(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3355));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1346 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1347 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3437), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1348 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3437));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1349 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1350 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3187), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1351 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1613), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3187));
OA21X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1352 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3458), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1613));
OAI31X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1353 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145), .A2(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3458));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1354 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1355 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2933), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1356 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2468), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2933));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1357 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2313), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2468));
AOI31X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1358 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510), .A2(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2313));
OR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1359 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741));
MXI2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1360 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__60), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__61), .S0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47]));
NAND2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1361 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1362 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[46]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159));
NOR2BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1363 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56));
NOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1364 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1365 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1552), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1366 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1367 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1982), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1368 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2410), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1552), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1982));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1369 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[45]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2410), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1370 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5705), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[46]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[45]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1371 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[22]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5705));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1372 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[44]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1373 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5766), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[45]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[44]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1374 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[21]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5766));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1375 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2908), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1376 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3240), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1377 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1378 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1711), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1379 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3240), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1711));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1380 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3339), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1381 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1802), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2908), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3339));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1382 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[43]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1802), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1383 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5719), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[44]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[43]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1384 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[20]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5719));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1385 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[42]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1386 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5669), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[43]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[42]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1387 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[19]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5669));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1388 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2303), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1389 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1390 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2734), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1391 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3160), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2303), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2734));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1392 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[41]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3160), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1393 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5732), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[42]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[41]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1394 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[18]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5732));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1395 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[40]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1396 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5684), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[41]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[40]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1397 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[17]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5684));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1398 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1399 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1400 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2558), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1401 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[39]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2558), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1402 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5747), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[40]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[39]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1403 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[16]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5747));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1404 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[38]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1405 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5697), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[39]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[38]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1406 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[15]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5697));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1407 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1408 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2809), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1409 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[37]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2809), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1410 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5759), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[38]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[37]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1411 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[14]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5759));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1412 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[36]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1413 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5711), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[37]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[36]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1414 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[13]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5711));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1415 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1416 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1417 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3053), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1418 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[35]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3053), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1419 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5776), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[36]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[35]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1420 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[12]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5776));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1421 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[34]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1422 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5727), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[35]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[34]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1423 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[11]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5727));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1424 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1425 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3305), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1426 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[33]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3305), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1427 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5677), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[34]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[33]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1428 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[10]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5677));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1429 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[32]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1430 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5741), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[33]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[32]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1431 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[9]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5741));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1432 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2698), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1433 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3136), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1434 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2676), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1435 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3102), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1436 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2676), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3102));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1437 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1605), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1438 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3136), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1605));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1439 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3125), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1440 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1595), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2698), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3125));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1441 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[31]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1595), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1442 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5692), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[32]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[31]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1443 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[8]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5692));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1444 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[30]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1445 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5755), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[31]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[30]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1446 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[7]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5755));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1447 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2093), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1448 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1449 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2524), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1450 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2950), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2093), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2524));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1451 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[29]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2950), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1452 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5707), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[30]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[29]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1453 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[6]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5707));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1454 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[28]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1455 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5770), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[29]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[28]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1456 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[5]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5770));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1457 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1458 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2346), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1459 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[27]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2346), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1460 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5722), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[28]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[27]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1461 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[4]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5722));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1462 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[26]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1463 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5672), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[27]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[26]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1464 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[3]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5672));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1465 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1466 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2596), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1467 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[25]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2596), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1468 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5735), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[26]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[25]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1469 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[2]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5735));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1470 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[24]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1471 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5687), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[25]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[24]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1472 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[1]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5687));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1473 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1988), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1474 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2781), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1475 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3210), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006));
AOI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1476 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1678), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2781), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3210));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1477 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2420), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871));
OAI21XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1478 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2845), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1988), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1678), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2420));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1479 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[23]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2845), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1480 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5750), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[24]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[23]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1481 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[0]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5750));
OR3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1482 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[7]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1483 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1484 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]));
INVXL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1485 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0]));
NOR2BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1486 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1487 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641));
NOR3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1488 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631));
NAND3XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1489 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5625), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620), .C(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1490 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[7]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5625), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1491 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5700), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[7]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]));
OAI2BB1X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1492 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[30]), .A0N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56), .A1N(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[7]), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5700));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1493 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[7]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1494 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5627), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1495 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[6]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5627), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1496 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5762), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[6]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1497 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[29]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5762));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1498 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[5]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1499 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5714), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[5]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1500 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[28]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5714));
NOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1501 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5618), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1502 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[4]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5618));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1503 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5778), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[4]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1504 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[27]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5778));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1505 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[3]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1506 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5729), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[3]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1507 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[26]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5729));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1508 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[2]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1509 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5680), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[2]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1510 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[25]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5680));
XNOR2X1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1511 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[1]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0]), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1512 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5743), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[1]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1513 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[24]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5743));
AOI22XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1514 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5694), .A0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0]), .A1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682), .B0(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767), .B1(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0]));
NAND2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1515 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[23]), .A(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5694));
XOR2XL DFT_compute_cynw_cm_float_mul_E8_M23_2_I1516 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__33), .A(a_sign), .B(b_sign));
NOR2BX1 DFT_compute_cynw_cm_float_mul_E8_M23_2_I1517 (.Y(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[31]), .AN(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__33), .B(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29));
EDFFHQX1 x_reg_0__I1518 (.Q(x[0]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_1__I1519 (.Q(x[1]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_2__I1520 (.Q(x[2]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_3__I1521 (.Q(x[3]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_4__I1522 (.Q(x[4]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_5__I1523 (.Q(x[5]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_6__I1524 (.Q(x[6]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__I1525 (.Q(x[7]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_8__I1526 (.Q(x[8]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_9__I1527 (.Q(x[9]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_10__I1528 (.Q(x[10]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_11__I1529 (.Q(x[11]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_12__I1530 (.Q(x[12]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_13__I1531 (.Q(x[13]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_14__I1532 (.Q(x[14]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_15__I1533 (.Q(x[15]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_16__I1534 (.Q(x[16]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_17__I1535 (.Q(x[17]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_18__I1536 (.Q(x[18]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_19__I1537 (.Q(x[19]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__I1538 (.Q(x[20]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__I1539 (.Q(x[21]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__I1540 (.Q(x[22]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__I1541 (.Q(x[23]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[23]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__I1542 (.Q(x[24]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_25__I1543 (.Q(x[25]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_26__I1544 (.Q(x[26]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[26]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_27__I1545 (.Q(x[27]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[27]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_28__I1546 (.Q(x[28]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[28]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_29__I1547 (.Q(x[29]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__I1548 (.Q(x[30]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[30]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__I1549 (.Q(x[31]), .D(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[31]), .E(bdw_enable), .CK(aclk));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[0] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[1] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[2] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[3] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[4] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[5] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[6] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[7] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[8] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[9] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[10] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[11] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[12] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[13] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[14] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[15] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[16] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[17] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[18] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[19] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[20] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[21] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[22] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[0] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[1] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[2] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[3] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[4] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[5] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[6] = 1'B0;
endmodule

/* CADENCE  vbH1Swjbrhk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



