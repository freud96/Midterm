/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:13 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_div_ieee_E8_M23_0 (
	clk,
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	accept,
	x
	); /* architecture "gate_level" */ 
input  clk;
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input  accept;
output [31:0] x;
wire [31:0] inst_cellmath__8,
	inst_cellmath__9;
wire  inst_cellmath__11;
wire [3:0] inst_cellmath__12,
	inst_cellmath__13;
wire [25:0] inst_cellmath__14,
	inst_cellmath__16,
	inst_cellmath__17;
wire [4:0] inst_cellmath__22,
	inst_cellmath__23;
wire [6:0] inst_lookup0_cellmath__27;
wire [2:0] inst_lookup0_cellmath__29;
wire [25:0] inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__34,
	inst_cellmath__35,
	inst_cellmath__38__W0,
	inst_cellmath__38__W1,
	inst_cellmath__39__W0,
	inst_cellmath__39__W1;
wire [28:0] inst_cellmath__40,
	inst_cellmath__41,
	inst_cellmath__42,
	inst_cellmath__43,
	inst_cellmath__44,
	inst_cellmath__45,
	inst_cellmath__46,
	inst_cellmath__47;
wire [6:0] inst_it2_lookup1_cellmath__53;
wire [2:0] inst_it2_lookup1_cellmath__55;
wire [25:0] inst_it2_cellmath__56,
	inst_it2_cellmath__57,
	inst_it2_cellmath__60,
	inst_it2_cellmath__61,
	inst_it2_cellmath__62__W0,
	inst_it2_cellmath__62__W1,
	inst_it2_cellmath__63__W1;
wire [9:0] inst_cellmath__67,
	inst_cellmath__68;
wire  inst_cellmath__69,
	inst_cellmath__70,
	inst_cellmath__71,
	inst_cellmath__72,
	inst_cellmath__73,
	inst_cellmath__74,
	inst_cellmath__75,
	inst_cellmath__76,
	inst_cellmath__77,
	inst_cellmath__78,
	inst_cellmath__79,
	inst_cellmath__80,
	inst_cellmath__83,
	inst_cellmath__84,
	inst_cellmath__85,
	inst_cellmath__86,
	inst_cellmath__87,
	inst_cellmath__88,
	inst_cellmath__89,
	inst_cellmath__91,
	inst_cellmath__96,
	inst_cellmath__100,
	inst_cellmath__101,
	inst_cellmath__102,
	inst_cellmath__103,
	inst_cellmath__104,
	inst_cellmath__105,
	inst_cellmath__106,
	inst_cellmath__109;
wire [7:0] inst_cellmath__110,
	inst_cellmath__111;
wire [21:0] inst_cellmath__112;
wire [31:0] inst_cellmath__113;
wire [25:0] inst_cellmath__120;
wire  inst_cellmath__122;
wire [28:0] inst_cellmath__124;
wire [22:0] inst_cellmath__125;
wire  inst_cellmath__126,
	inst_cellmath__127;
wire [22:0] inst_cellmath__129;
wire  inst_cellmath__135,
	inst_cellmath__136,
	inst_cellmath__137;
wire N1322,N1324,N1325,N1326,N1327,N1386,N1387 
	,N1388,N1417,N1555,N1675,N1677,N1678,N1679,N1680 
	,N1681,N1682,N1750,N1751,N1752,N1753,N1754,N1755 
	,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763 
	,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771 
	,N1772,N1922,N2045,N2046,N2047,N2048,N2049,N2050 
	,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058 
	,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066 
	,N2067,N2068,N2150,N2151,N2152,N2153,N2154,N2155 
	,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163 
	,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171 
	,N2172,N2173,N2201,N2202,N2203,N2204,N2205,N2206 
	,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214 
	,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222 
	,N2223,N2224,N2254,N2255,N2256,N2257,N2258,N2259 
	,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267 
	,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275 
	,N2276,N2277,N4587,N4594,N12283,N12286,N12290,N12294 
	,N12297,N12310,N12313,N12314,N12315,N12318,N12322,N12323 
	,N12326,N12362,N12363,N12364,N12365,N12366,N12368,N12369 
	,N12371,N12373,N12375,N12376,N12377,N12378,N12379,N12380 
	,N12381,N12383,N12384,N12385,N12386,N12387,N12389,N12392 
	,N12394,N12395,N12396,N12397,N12399,N12400,N12401,N12403 
	,N12404,N12405,N12407,N12408,N12409,N12410,N12411,N12414 
	,N12417,N12418,N12419,N12421,N12573,N12658,N12720,N12723 
	,N12729,N12732,N12736,N12738,N12740,N12744,N12751,N12754 
	,N12761,N12764,N12771,N12774,N12782,N12785,N12791,N12794 
	,N12797,N12803,N12806,N12811,N12813,N12870,N12983,N13206 
	,N13373,N13376,N13380,N13384,N13387,N13401,N13402,N13403 
	,N13404,N13405,N13408,N13410,N13412,N13414,N13415,N13417 
	,N13419,N13420,N13422,N13423,N13424,N13425,N13426,N13428 
	,N13431,N13433,N13434,N13435,N13436,N13438,N13439,N13440 
	,N13442,N13444,N13447,N13448,N13449,N13450,N13453,N13456 
	,N13457,N13458,N13460,N13614,N13658,N13661,N13665,N13667 
	,N13673,N13677,N13680,N13685,N13689,N13692,N13697,N13704 
	,N13705,N13712,N13716,N13719,N13722,N13725,N13730,N13737 
	,N13738,N13745,N13750,N13753,N13758,N13935,N13952,N14010 
	,N14012,N14016,N14018,N14020,N14025,N14027,N14030,N14033 
	,N14035,N14038,N14043,N14045,N14047,N14053,N14055,N14058 
	,N14061,N14063,N14070,N14072,N14077,N14146,N14149,N14153 
	,N14158,N14160,N14165,N14169,N14173,N14177,N14179,N14181 
	,N14182,N14185,N14213,N14214,N14594,N14648,N14981,N15334 
	,N15398,N15400,N15401,N15403,N15404,N15406,N15409,N15411 
	,N15412,N15413,N15415,N15417,N15418,N15421,N15423,N15424 
	,N15426,N15429,N15430,N15431,N15432,N15434,N15435,N15436 
	,N15440,N15443,N15444,N15486,N15491,N15495,N15497,N15503 
	,N15504,N15506,N15511,N15518,N15523,N15552,N15554,N15560 
	,N15579,N15582,N15583,N15585,N15589,N15605,N15608,N15618 
	,N15631,N15636,N15640,N15656,N15660,N15663,N15666,N15679 
	,N15681,N15699,N15702,N15710,N15711,N15720,N15722,N15724 
	,N15726,N15728,N15730,N15732,N15733,N15736,N15758,N15759 
	,N15762,N15770,N15779,N15780,N15782,N15784,N15786,N15788 
	,N15790,N15792,N15795,N15830,N15834,N15837,N15840,N15848 
	,N15852,N15855,N15858,N15898,N15943,N15964,N16014,N16016 
	,N16019,N16030,N16033,N16051,N16052,N16055,N16059,N16064 
	,N16067,N16070,N16076,N16080,N16083,N16086,N16122,N16178 
	,N18408,N18417,N28016,N28021,N28027;
reg inst_cellmath__0_0_0__I0_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_0__I0_QOUT <= inst_cellmath__113[0];
	end
assign x[0] = inst_cellmath__0_0_0__I0_QOUT;
reg inst_cellmath__0_0_1__I1_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_1__I1_QOUT <= inst_cellmath__113[1];
	end
assign x[1] = inst_cellmath__0_0_1__I1_QOUT;
reg inst_cellmath__0_0_2__I2_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_2__I2_QOUT <= inst_cellmath__113[2];
	end
assign x[2] = inst_cellmath__0_0_2__I2_QOUT;
reg inst_cellmath__0_0_3__I3_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_3__I3_QOUT <= inst_cellmath__113[3];
	end
assign x[3] = inst_cellmath__0_0_3__I3_QOUT;
reg inst_cellmath__0_0_4__I4_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_4__I4_QOUT <= inst_cellmath__113[4];
	end
assign x[4] = inst_cellmath__0_0_4__I4_QOUT;
reg inst_cellmath__0_0_5__I5_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_5__I5_QOUT <= inst_cellmath__113[5];
	end
assign x[5] = inst_cellmath__0_0_5__I5_QOUT;
reg inst_cellmath__0_0_6__I6_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_6__I6_QOUT <= inst_cellmath__113[6];
	end
assign x[6] = inst_cellmath__0_0_6__I6_QOUT;
reg inst_cellmath__0_0_7__I7_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_7__I7_QOUT <= inst_cellmath__113[7];
	end
assign x[7] = inst_cellmath__0_0_7__I7_QOUT;
reg inst_cellmath__0_0_8__I8_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_8__I8_QOUT <= inst_cellmath__113[8];
	end
assign x[8] = inst_cellmath__0_0_8__I8_QOUT;
reg inst_cellmath__0_0_9__I9_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_9__I9_QOUT <= inst_cellmath__113[9];
	end
assign x[9] = inst_cellmath__0_0_9__I9_QOUT;
reg inst_cellmath__0_0_10__I10_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_10__I10_QOUT <= inst_cellmath__113[10];
	end
assign x[10] = inst_cellmath__0_0_10__I10_QOUT;
reg inst_cellmath__0_0_11__I11_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_11__I11_QOUT <= inst_cellmath__113[11];
	end
assign x[11] = inst_cellmath__0_0_11__I11_QOUT;
reg inst_cellmath__0_0_12__I12_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_12__I12_QOUT <= inst_cellmath__113[12];
	end
assign x[12] = inst_cellmath__0_0_12__I12_QOUT;
reg inst_cellmath__0_0_13__I13_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_13__I13_QOUT <= inst_cellmath__113[13];
	end
assign x[13] = inst_cellmath__0_0_13__I13_QOUT;
reg inst_cellmath__0_0_14__I14_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_14__I14_QOUT <= inst_cellmath__113[14];
	end
assign x[14] = inst_cellmath__0_0_14__I14_QOUT;
reg inst_cellmath__0_0_15__I15_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_15__I15_QOUT <= inst_cellmath__113[15];
	end
assign x[15] = inst_cellmath__0_0_15__I15_QOUT;
reg inst_cellmath__0_0_16__I16_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_16__I16_QOUT <= inst_cellmath__113[16];
	end
assign x[16] = inst_cellmath__0_0_16__I16_QOUT;
reg inst_cellmath__0_0_17__I17_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_17__I17_QOUT <= inst_cellmath__113[17];
	end
assign x[17] = inst_cellmath__0_0_17__I17_QOUT;
reg inst_cellmath__0_0_18__I18_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_18__I18_QOUT <= inst_cellmath__113[18];
	end
assign x[18] = inst_cellmath__0_0_18__I18_QOUT;
reg inst_cellmath__0_0_19__I19_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_19__I19_QOUT <= inst_cellmath__113[19];
	end
assign x[19] = inst_cellmath__0_0_19__I19_QOUT;
reg inst_cellmath__0_0_20__I20_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_20__I20_QOUT <= inst_cellmath__113[20];
	end
assign x[20] = inst_cellmath__0_0_20__I20_QOUT;
reg inst_cellmath__0_0_21__I21_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_21__I21_QOUT <= inst_cellmath__113[21];
	end
assign x[21] = inst_cellmath__0_0_21__I21_QOUT;
reg inst_cellmath__0_0_22__I22_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_22__I22_QOUT <= inst_cellmath__113[22];
	end
assign x[22] = inst_cellmath__0_0_22__I22_QOUT;
reg inst_cellmath__0_0_23__I23_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_23__I23_QOUT <= inst_cellmath__113[23];
	end
assign x[23] = inst_cellmath__0_0_23__I23_QOUT;
reg inst_cellmath__0_0_24__I24_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_24__I24_QOUT <= inst_cellmath__113[24];
	end
assign x[24] = inst_cellmath__0_0_24__I24_QOUT;
reg inst_cellmath__0_0_25__I25_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_25__I25_QOUT <= inst_cellmath__113[25];
	end
assign x[25] = inst_cellmath__0_0_25__I25_QOUT;
reg inst_cellmath__0_0_26__I26_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_26__I26_QOUT <= inst_cellmath__113[26];
	end
assign x[26] = inst_cellmath__0_0_26__I26_QOUT;
reg inst_cellmath__0_0_27__I27_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_27__I27_QOUT <= inst_cellmath__113[27];
	end
assign x[27] = inst_cellmath__0_0_27__I27_QOUT;
reg inst_cellmath__0_0_28__I28_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_28__I28_QOUT <= inst_cellmath__113[28];
	end
assign x[28] = inst_cellmath__0_0_28__I28_QOUT;
reg inst_cellmath__0_0_29__I29_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_29__I29_QOUT <= inst_cellmath__113[29];
	end
assign x[29] = inst_cellmath__0_0_29__I29_QOUT;
reg inst_cellmath__0_0_30__I30_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_30__I30_QOUT <= inst_cellmath__113[30];
	end
assign x[30] = inst_cellmath__0_0_30__I30_QOUT;
reg inst_cellmath__0_0_31__I31_QOUT;
always @ (posedge clk)
	if (N4594==1'b1) begin inst_cellmath__0_0_31__I31_QOUT <= inst_cellmath__113[31];
	end
assign x[31] = inst_cellmath__0_0_31__I31_QOUT;
reg inst_cellmath__9_0_0__I32_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_0__I32_QOUT <= b_man[0];
	end
assign inst_cellmath__9[0] = inst_cellmath__9_0_0__I32_QOUT;
reg inst_cellmath__9_0_1__I33_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_1__I33_QOUT <= b_man[1];
	end
assign inst_cellmath__9[1] = inst_cellmath__9_0_1__I33_QOUT;
reg inst_cellmath__9_0_2__I34_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_2__I34_QOUT <= b_man[2];
	end
assign inst_cellmath__9[2] = inst_cellmath__9_0_2__I34_QOUT;
reg inst_cellmath__9_0_3__I35_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_3__I35_QOUT <= b_man[3];
	end
assign inst_cellmath__9[3] = inst_cellmath__9_0_3__I35_QOUT;
reg inst_cellmath__9_0_4__I36_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_4__I36_QOUT <= b_man[4];
	end
assign inst_cellmath__9[4] = inst_cellmath__9_0_4__I36_QOUT;
reg inst_cellmath__9_0_5__I37_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_5__I37_QOUT <= b_man[5];
	end
assign inst_cellmath__9[5] = inst_cellmath__9_0_5__I37_QOUT;
reg inst_cellmath__9_0_6__I38_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_6__I38_QOUT <= b_man[6];
	end
assign inst_cellmath__9[6] = inst_cellmath__9_0_6__I38_QOUT;
reg inst_cellmath__9_0_7__I39_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_7__I39_QOUT <= b_man[7];
	end
assign inst_cellmath__9[7] = inst_cellmath__9_0_7__I39_QOUT;
reg inst_cellmath__9_0_8__I40_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_8__I40_QOUT <= b_man[8];
	end
assign inst_cellmath__9[8] = inst_cellmath__9_0_8__I40_QOUT;
reg inst_cellmath__9_0_9__I41_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_9__I41_QOUT <= b_man[9];
	end
assign inst_cellmath__9[9] = inst_cellmath__9_0_9__I41_QOUT;
reg inst_cellmath__9_0_10__I42_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_10__I42_QOUT <= b_man[10];
	end
assign inst_cellmath__9[10] = inst_cellmath__9_0_10__I42_QOUT;
reg inst_cellmath__9_0_11__I43_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_11__I43_QOUT <= b_man[11];
	end
assign inst_cellmath__9[11] = inst_cellmath__9_0_11__I43_QOUT;
reg inst_cellmath__9_0_12__I44_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_12__I44_QOUT <= b_man[12];
	end
assign inst_cellmath__9[12] = inst_cellmath__9_0_12__I44_QOUT;
reg inst_cellmath__9_0_13__I45_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_13__I45_QOUT <= b_man[13];
	end
assign inst_cellmath__9[13] = inst_cellmath__9_0_13__I45_QOUT;
reg inst_cellmath__9_0_14__I46_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_14__I46_QOUT <= b_man[14];
	end
assign inst_cellmath__9[14] = inst_cellmath__9_0_14__I46_QOUT;
reg inst_cellmath__9_0_15__I47_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_15__I47_QOUT <= b_man[15];
	end
assign inst_cellmath__9[15] = inst_cellmath__9_0_15__I47_QOUT;
reg inst_cellmath__9_0_16__I48_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_16__I48_QOUT <= b_man[16];
	end
assign inst_cellmath__9[16] = inst_cellmath__9_0_16__I48_QOUT;
reg inst_cellmath__9_0_17__I49_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_17__I49_QOUT <= b_man[17];
	end
assign inst_cellmath__9[17] = inst_cellmath__9_0_17__I49_QOUT;
reg inst_cellmath__9_0_18__I50_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_18__I50_QOUT <= b_man[18];
	end
assign inst_cellmath__9[18] = inst_cellmath__9_0_18__I50_QOUT;
reg inst_cellmath__9_0_19__I51_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_19__I51_QOUT <= b_man[19];
	end
assign inst_cellmath__9[19] = inst_cellmath__9_0_19__I51_QOUT;
reg inst_cellmath__9_0_20__I52_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_20__I52_QOUT <= b_man[20];
	end
assign inst_cellmath__9[20] = inst_cellmath__9_0_20__I52_QOUT;
reg inst_cellmath__9_0_21__I53_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_21__I53_QOUT <= b_man[21];
	end
assign inst_it2_lookup1_cellmath__53[0] = inst_cellmath__9_0_21__I53_QOUT;
reg inst_cellmath__9_0_22__I54_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_22__I54_QOUT <= b_man[22];
	end
assign inst_it2_lookup1_cellmath__53[1] = inst_cellmath__9_0_22__I54_QOUT;
reg inst_cellmath__9_0_23__I55_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_23__I55_QOUT <= b_exp[0];
	end
assign inst_cellmath__9[23] = inst_cellmath__9_0_23__I55_QOUT;
reg inst_cellmath__9_0_24__I56_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_24__I56_QOUT <= b_exp[1];
	end
assign inst_cellmath__9[24] = inst_cellmath__9_0_24__I56_QOUT;
reg inst_cellmath__9_0_25__I57_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_25__I57_QOUT <= b_exp[2];
	end
assign inst_cellmath__9[25] = inst_cellmath__9_0_25__I57_QOUT;
reg inst_cellmath__9_0_26__I58_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_26__I58_QOUT <= b_exp[3];
	end
assign inst_cellmath__9[26] = inst_cellmath__9_0_26__I58_QOUT;
reg inst_cellmath__9_0_27__I59_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_27__I59_QOUT <= b_exp[4];
	end
assign inst_cellmath__9[27] = inst_cellmath__9_0_27__I59_QOUT;
reg inst_cellmath__9_0_28__I60_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_28__I60_QOUT <= b_exp[5];
	end
assign inst_cellmath__9[28] = inst_cellmath__9_0_28__I60_QOUT;
reg inst_cellmath__9_0_29__I61_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_29__I61_QOUT <= b_exp[6];
	end
assign inst_cellmath__9[29] = inst_cellmath__9_0_29__I61_QOUT;
reg inst_cellmath__9_0_30__I62_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_30__I62_QOUT <= b_exp[7];
	end
assign inst_cellmath__9[30] = inst_cellmath__9_0_30__I62_QOUT;
reg inst_cellmath__9_0_31__I63_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__9_0_31__I63_QOUT <= b_sign;
	end
assign inst_cellmath__9[31] = inst_cellmath__9_0_31__I63_QOUT;
reg inst_cellmath__11_0_I64_QOUT;
always @ (posedge clk)
	inst_cellmath__11_0_I64_QOUT <= accept;
assign inst_cellmath__11 = inst_cellmath__11_0_I64_QOUT;
reg inst_cellmath__16_0_1__I65_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_1__I65_QOUT <= inst_cellmath__14[1];
assign inst_cellmath__16[1] = inst_cellmath__16_0_1__I65_QOUT;
reg inst_cellmath__16_0_2__I66_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_2__I66_QOUT <= inst_cellmath__14[2];
assign inst_cellmath__16[2] = inst_cellmath__16_0_2__I66_QOUT;
reg inst_cellmath__16_0_3__I67_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_3__I67_QOUT <= inst_cellmath__14[3];
assign inst_cellmath__16[3] = inst_cellmath__16_0_3__I67_QOUT;
reg inst_cellmath__16_0_4__I68_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_4__I68_QOUT <= inst_cellmath__14[4];
assign inst_cellmath__16[4] = inst_cellmath__16_0_4__I68_QOUT;
reg inst_cellmath__16_0_5__I69_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_5__I69_QOUT <= inst_cellmath__14[5];
assign inst_cellmath__16[5] = inst_cellmath__16_0_5__I69_QOUT;
reg inst_cellmath__16_0_6__I70_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_6__I70_QOUT <= inst_cellmath__14[6];
assign inst_cellmath__16[6] = inst_cellmath__16_0_6__I70_QOUT;
reg inst_cellmath__16_0_7__I71_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_7__I71_QOUT <= inst_cellmath__14[7];
assign inst_cellmath__16[7] = inst_cellmath__16_0_7__I71_QOUT;
reg inst_cellmath__16_0_8__I72_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_8__I72_QOUT <= inst_cellmath__14[8];
assign inst_cellmath__16[8] = inst_cellmath__16_0_8__I72_QOUT;
reg inst_cellmath__16_0_9__I73_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_9__I73_QOUT <= inst_cellmath__14[9];
assign inst_cellmath__16[9] = inst_cellmath__16_0_9__I73_QOUT;
reg inst_cellmath__16_0_10__I74_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_10__I74_QOUT <= inst_cellmath__14[10];
assign inst_cellmath__16[10] = inst_cellmath__16_0_10__I74_QOUT;
reg inst_cellmath__16_0_11__I75_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_11__I75_QOUT <= inst_cellmath__14[11];
assign inst_cellmath__16[11] = inst_cellmath__16_0_11__I75_QOUT;
reg inst_cellmath__16_0_12__I76_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_12__I76_QOUT <= inst_cellmath__14[12];
assign inst_cellmath__16[12] = inst_cellmath__16_0_12__I76_QOUT;
reg inst_cellmath__16_0_13__I77_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_13__I77_QOUT <= inst_cellmath__14[13];
assign inst_cellmath__16[13] = inst_cellmath__16_0_13__I77_QOUT;
reg inst_cellmath__16_0_14__I78_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_14__I78_QOUT <= inst_cellmath__14[14];
assign inst_cellmath__16[14] = inst_cellmath__16_0_14__I78_QOUT;
reg inst_cellmath__16_0_15__I79_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_15__I79_QOUT <= inst_cellmath__14[15];
assign inst_cellmath__16[15] = inst_cellmath__16_0_15__I79_QOUT;
reg inst_cellmath__16_0_16__I80_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_16__I80_QOUT <= inst_cellmath__14[16];
assign inst_cellmath__16[16] = inst_cellmath__16_0_16__I80_QOUT;
reg inst_cellmath__16_0_17__I81_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_17__I81_QOUT <= inst_cellmath__14[17];
assign inst_cellmath__16[17] = inst_cellmath__16_0_17__I81_QOUT;
reg inst_cellmath__16_0_18__I82_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_18__I82_QOUT <= inst_cellmath__14[18];
assign inst_cellmath__16[18] = inst_cellmath__16_0_18__I82_QOUT;
reg inst_cellmath__16_0_19__I83_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_19__I83_QOUT <= inst_cellmath__14[19];
assign inst_cellmath__16[19] = inst_cellmath__16_0_19__I83_QOUT;
reg inst_cellmath__16_0_20__I84_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_20__I84_QOUT <= inst_cellmath__14[20];
assign inst_cellmath__16[20] = inst_cellmath__16_0_20__I84_QOUT;
reg inst_cellmath__16_0_21__I85_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_21__I85_QOUT <= inst_cellmath__14[21];
assign inst_cellmath__16[21] = inst_cellmath__16_0_21__I85_QOUT;
reg inst_cellmath__16_0_22__I86_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_22__I86_QOUT <= inst_cellmath__14[22];
assign inst_cellmath__16[22] = inst_cellmath__16_0_22__I86_QOUT;
reg inst_cellmath__16_0_23__I87_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_23__I87_QOUT <= inst_cellmath__14[23];
assign inst_cellmath__16[23] = inst_cellmath__16_0_23__I87_QOUT;
reg inst_cellmath__16_0_24__I88_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_24__I88_QOUT <= inst_cellmath__14[24];
assign inst_cellmath__16[24] = inst_cellmath__16_0_24__I88_QOUT;
reg inst_cellmath__16_0_25__I89_QOUT;
always @ (posedge clk)
	inst_cellmath__16_0_25__I89_QOUT <= inst_cellmath__14[25];
assign inst_cellmath__16[25] = inst_cellmath__16_0_25__I89_QOUT;
reg inst_cellmath__17_0_1__I91_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_1__I91_QOUT <= inst_it2_cellmath__63__W1[1];
assign inst_cellmath__17[1] = inst_cellmath__17_0_1__I91_QOUT;
reg inst_cellmath__17_0_2__I92_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_2__I92_QOUT <= inst_it2_cellmath__63__W1[2];
assign inst_cellmath__17[2] = inst_cellmath__17_0_2__I92_QOUT;
reg inst_cellmath__17_0_3__I93_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_3__I93_QOUT <= inst_it2_cellmath__63__W1[3];
assign inst_cellmath__17[3] = inst_cellmath__17_0_3__I93_QOUT;
reg inst_cellmath__17_0_4__I94_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_4__I94_QOUT <= inst_it2_cellmath__63__W1[4];
assign inst_cellmath__17[4] = inst_cellmath__17_0_4__I94_QOUT;
reg inst_cellmath__17_0_5__I95_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_5__I95_QOUT <= inst_it2_cellmath__63__W1[5];
assign inst_cellmath__17[5] = inst_cellmath__17_0_5__I95_QOUT;
reg inst_cellmath__17_0_6__I96_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_6__I96_QOUT <= inst_it2_cellmath__63__W1[6];
assign inst_cellmath__17[6] = inst_cellmath__17_0_6__I96_QOUT;
reg inst_cellmath__17_0_7__I97_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_7__I97_QOUT <= inst_it2_cellmath__63__W1[7];
assign inst_cellmath__17[7] = inst_cellmath__17_0_7__I97_QOUT;
reg inst_cellmath__17_0_8__I98_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_8__I98_QOUT <= inst_it2_cellmath__63__W1[8];
assign inst_cellmath__17[8] = inst_cellmath__17_0_8__I98_QOUT;
reg inst_cellmath__17_0_9__I99_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_9__I99_QOUT <= inst_it2_cellmath__63__W1[9];
assign inst_cellmath__17[9] = inst_cellmath__17_0_9__I99_QOUT;
reg inst_cellmath__17_0_10__I100_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_10__I100_QOUT <= inst_it2_cellmath__63__W1[10];
assign inst_cellmath__17[10] = inst_cellmath__17_0_10__I100_QOUT;
reg inst_cellmath__17_0_11__I101_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_11__I101_QOUT <= inst_it2_cellmath__63__W1[11];
assign inst_cellmath__17[11] = inst_cellmath__17_0_11__I101_QOUT;
reg inst_cellmath__17_0_12__I102_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_12__I102_QOUT <= inst_it2_cellmath__63__W1[12];
assign inst_cellmath__17[12] = inst_cellmath__17_0_12__I102_QOUT;
reg inst_cellmath__17_0_13__I103_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_13__I103_QOUT <= inst_it2_cellmath__63__W1[13];
assign inst_cellmath__17[13] = inst_cellmath__17_0_13__I103_QOUT;
reg inst_cellmath__17_0_14__I104_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_14__I104_QOUT <= inst_it2_cellmath__63__W1[14];
assign inst_cellmath__17[14] = inst_cellmath__17_0_14__I104_QOUT;
reg inst_cellmath__17_0_15__I105_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_15__I105_QOUT <= inst_it2_cellmath__63__W1[15];
assign inst_cellmath__17[15] = inst_cellmath__17_0_15__I105_QOUT;
reg inst_cellmath__17_0_16__I106_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_16__I106_QOUT <= inst_it2_cellmath__63__W1[16];
assign inst_cellmath__17[16] = inst_cellmath__17_0_16__I106_QOUT;
reg inst_cellmath__17_0_17__I107_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_17__I107_QOUT <= inst_it2_cellmath__63__W1[17];
assign inst_cellmath__17[17] = inst_cellmath__17_0_17__I107_QOUT;
reg inst_cellmath__17_0_18__I108_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_18__I108_QOUT <= inst_it2_cellmath__63__W1[18];
assign inst_cellmath__17[18] = inst_cellmath__17_0_18__I108_QOUT;
reg inst_cellmath__17_0_19__I109_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_19__I109_QOUT <= inst_it2_cellmath__63__W1[19];
assign inst_cellmath__17[19] = inst_cellmath__17_0_19__I109_QOUT;
reg inst_cellmath__17_0_20__I110_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_20__I110_QOUT <= inst_it2_cellmath__63__W1[20];
assign inst_cellmath__17[20] = inst_cellmath__17_0_20__I110_QOUT;
reg inst_cellmath__17_0_21__I111_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_21__I111_QOUT <= inst_it2_cellmath__63__W1[21];
assign inst_cellmath__17[21] = inst_cellmath__17_0_21__I111_QOUT;
reg inst_cellmath__17_0_22__I112_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_22__I112_QOUT <= inst_it2_cellmath__63__W1[22];
assign inst_cellmath__17[22] = inst_cellmath__17_0_22__I112_QOUT;
reg inst_cellmath__17_0_23__I113_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_23__I113_QOUT <= inst_it2_cellmath__63__W1[23];
assign inst_cellmath__17[23] = inst_cellmath__17_0_23__I113_QOUT;
reg inst_cellmath__17_0_24__I114_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_24__I114_QOUT <= inst_it2_cellmath__63__W1[24];
assign inst_cellmath__17[24] = inst_cellmath__17_0_24__I114_QOUT;
reg inst_cellmath__17_0_25__I115_QOUT;
always @ (posedge clk)
	inst_cellmath__17_0_25__I115_QOUT <= inst_it2_cellmath__63__W1[25];
assign inst_cellmath__17[25] = inst_cellmath__17_0_25__I115_QOUT;
assign {N12290, inst_cellmath__23[0]} = {1'B0, inst_cellmath__17[21]} + {1'B0, inst_cellmath__16[21]};
assign {N12286, inst_cellmath__23[1]} = {1'B0, inst_cellmath__17[22]} + {1'B0, inst_cellmath__16[22]} + {1'B0, N12290};
assign {N12297, inst_cellmath__23[2]} = {1'B0, inst_cellmath__17[23]} + {1'B0, inst_cellmath__16[23]} + {1'B0, N12286};
assign {N12283, inst_cellmath__23[3]} = {1'B0, inst_cellmath__17[24]} + {1'B0, inst_cellmath__16[24]} + {1'B0, N12297};
assign {N12294, inst_cellmath__23[4]} = {1'B0, inst_cellmath__17[25]} + {1'B0, inst_cellmath__16[25]} + {1'B0, N12283};
reg inst_cellmath__8_0_0__I117_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_0__I117_QOUT <= a_man[0];
	end
assign inst_cellmath__8[0] = inst_cellmath__8_0_0__I117_QOUT;
reg inst_cellmath__8_0_1__I118_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_1__I118_QOUT <= a_man[1];
	end
assign inst_cellmath__8[1] = inst_cellmath__8_0_1__I118_QOUT;
reg inst_cellmath__8_0_2__I119_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_2__I119_QOUT <= a_man[2];
	end
assign inst_cellmath__8[2] = inst_cellmath__8_0_2__I119_QOUT;
reg inst_cellmath__8_0_3__I120_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_3__I120_QOUT <= a_man[3];
	end
assign inst_cellmath__8[3] = inst_cellmath__8_0_3__I120_QOUT;
reg inst_cellmath__8_0_4__I121_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_4__I121_QOUT <= a_man[4];
	end
assign inst_cellmath__8[4] = inst_cellmath__8_0_4__I121_QOUT;
reg inst_cellmath__8_0_5__I122_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_5__I122_QOUT <= a_man[5];
	end
assign inst_cellmath__8[5] = inst_cellmath__8_0_5__I122_QOUT;
reg inst_cellmath__8_0_6__I123_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_6__I123_QOUT <= a_man[6];
	end
assign inst_cellmath__8[6] = inst_cellmath__8_0_6__I123_QOUT;
reg inst_cellmath__8_0_7__I124_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_7__I124_QOUT <= a_man[7];
	end
assign inst_cellmath__8[7] = inst_cellmath__8_0_7__I124_QOUT;
reg inst_cellmath__8_0_8__I125_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_8__I125_QOUT <= a_man[8];
	end
assign inst_cellmath__8[8] = inst_cellmath__8_0_8__I125_QOUT;
reg inst_cellmath__8_0_9__I126_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_9__I126_QOUT <= a_man[9];
	end
assign inst_cellmath__8[9] = inst_cellmath__8_0_9__I126_QOUT;
reg inst_cellmath__8_0_10__I127_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_10__I127_QOUT <= a_man[10];
	end
assign inst_cellmath__8[10] = inst_cellmath__8_0_10__I127_QOUT;
reg inst_cellmath__8_0_11__I128_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_11__I128_QOUT <= a_man[11];
	end
assign inst_cellmath__8[11] = inst_cellmath__8_0_11__I128_QOUT;
reg inst_cellmath__8_0_12__I129_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_12__I129_QOUT <= a_man[12];
	end
assign inst_cellmath__8[12] = inst_cellmath__8_0_12__I129_QOUT;
reg inst_cellmath__8_0_13__I130_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_13__I130_QOUT <= a_man[13];
	end
assign inst_cellmath__8[13] = inst_cellmath__8_0_13__I130_QOUT;
reg inst_cellmath__8_0_14__I131_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_14__I131_QOUT <= a_man[14];
	end
assign inst_cellmath__8[14] = inst_cellmath__8_0_14__I131_QOUT;
reg inst_cellmath__8_0_15__I132_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_15__I132_QOUT <= a_man[15];
	end
assign inst_cellmath__8[15] = inst_cellmath__8_0_15__I132_QOUT;
reg inst_cellmath__8_0_16__I133_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_16__I133_QOUT <= a_man[16];
	end
assign inst_cellmath__8[16] = inst_cellmath__8_0_16__I133_QOUT;
reg inst_cellmath__8_0_17__I134_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_17__I134_QOUT <= a_man[17];
	end
assign inst_cellmath__8[17] = inst_cellmath__8_0_17__I134_QOUT;
reg inst_cellmath__8_0_18__I135_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_18__I135_QOUT <= a_man[18];
	end
assign inst_cellmath__8[18] = inst_cellmath__8_0_18__I135_QOUT;
reg inst_cellmath__8_0_19__I136_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_19__I136_QOUT <= a_man[19];
	end
assign inst_cellmath__8[19] = inst_cellmath__8_0_19__I136_QOUT;
reg inst_cellmath__8_0_20__I137_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_20__I137_QOUT <= a_man[20];
	end
assign inst_cellmath__8[20] = inst_cellmath__8_0_20__I137_QOUT;
reg inst_cellmath__8_0_21__I138_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_21__I138_QOUT <= a_man[21];
	end
assign inst_cellmath__8[21] = inst_cellmath__8_0_21__I138_QOUT;
reg inst_cellmath__8_0_22__I139_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_22__I139_QOUT <= a_man[22];
	end
assign inst_cellmath__8[22] = inst_cellmath__8_0_22__I139_QOUT;
reg inst_cellmath__8_0_23__I140_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_23__I140_QOUT <= a_exp[0];
	end
assign inst_cellmath__8[23] = inst_cellmath__8_0_23__I140_QOUT;
reg inst_cellmath__8_0_24__I141_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_24__I141_QOUT <= a_exp[1];
	end
assign inst_cellmath__8[24] = inst_cellmath__8_0_24__I141_QOUT;
reg inst_cellmath__8_0_25__I142_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_25__I142_QOUT <= a_exp[2];
	end
assign inst_cellmath__8[25] = inst_cellmath__8_0_25__I142_QOUT;
reg inst_cellmath__8_0_26__I143_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_26__I143_QOUT <= a_exp[3];
	end
assign inst_cellmath__8[26] = inst_cellmath__8_0_26__I143_QOUT;
reg inst_cellmath__8_0_27__I144_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_27__I144_QOUT <= a_exp[4];
	end
assign inst_cellmath__8[27] = inst_cellmath__8_0_27__I144_QOUT;
reg inst_cellmath__8_0_28__I145_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_28__I145_QOUT <= a_exp[5];
	end
assign inst_cellmath__8[28] = inst_cellmath__8_0_28__I145_QOUT;
reg inst_cellmath__8_0_29__I146_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_29__I146_QOUT <= a_exp[6];
	end
assign inst_cellmath__8[29] = inst_cellmath__8_0_29__I146_QOUT;
reg inst_cellmath__8_0_30__I147_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_30__I147_QOUT <= a_exp[7];
	end
assign inst_cellmath__8[30] = inst_cellmath__8_0_30__I147_QOUT;
reg inst_cellmath__8_0_31__I148_QOUT;
always @ (posedge clk)
	if (accept==1'b1) begin inst_cellmath__8_0_31__I148_QOUT <= a_sign;
	end
assign inst_cellmath__8[31] = inst_cellmath__8_0_31__I148_QOUT;
assign N1386 = !inst_cellmath__9[20];
assign N1387 = !inst_it2_lookup1_cellmath__53[0];
assign N1388 = !inst_it2_lookup1_cellmath__53[1];
assign N12322 = !(inst_cellmath__8[20] & N1386);
assign N12326 = !(inst_cellmath__8[21] | N1387);
assign N12313 = !(inst_cellmath__8[21] & N1387);
assign N12315 = !(inst_cellmath__8[22] | N1388);
assign N12318 = !(inst_cellmath__8[22] & N1388);
assign N12314 = (N12322 & N12313) | N12326;
assign inst_cellmath__22[4] = (N12314 & N12318) | N12315;
assign N12310 = !(N12313 & (!N12326));
assign N12323 = !(N12318 & (!N12315));
assign inst_cellmath__22[0] = inst_cellmath__8[20] ^ N1386;
assign inst_cellmath__22[1] = N12322 ^ N12310;
assign inst_cellmath__22[2] = N12314 ^ N12323;
assign inst_lookup0_cellmath__27[2] = (inst_cellmath__11 & inst_cellmath__22[0]) | ((!inst_cellmath__11) & inst_cellmath__23[0]);
assign inst_lookup0_cellmath__27[3] = (inst_cellmath__11 & inst_cellmath__22[1]) | ((!inst_cellmath__11) & inst_cellmath__23[1]);
assign inst_lookup0_cellmath__27[4] = (inst_cellmath__11 & inst_cellmath__22[2]) | ((!inst_cellmath__11) & inst_cellmath__23[2]);
assign inst_lookup0_cellmath__27[5] = (inst_cellmath__11 & inst_cellmath__22[4]) | ((!inst_cellmath__11) & inst_cellmath__23[3]);
assign inst_lookup0_cellmath__27[6] = (inst_cellmath__11 & inst_cellmath__22[4]) | ((!inst_cellmath__11) & inst_cellmath__23[4]);
assign N12397 = !inst_lookup0_cellmath__27[2];
assign N12386 = !inst_lookup0_cellmath__27[3];
assign N12381 = !(N12386 | N12397);
assign N12418 = !(N12397 | N1388);
assign N12379 = !(N1387 & N1388);
assign N12366 = !((inst_it2_lookup1_cellmath__53[1] & N12397) | (N12379 & inst_lookup0_cellmath__27[2]));
assign N12421 = !((N12366 & N12386) | (N12418 & inst_lookup0_cellmath__27[3]));
assign N12365 = !(inst_it2_lookup1_cellmath__53[1] & inst_lookup0_cellmath__27[2]);
assign N12373 = !(N12386 | N12365);
assign N12363 = !inst_lookup0_cellmath__27[4];
assign N12394 = !((N12421 & N12363) | (N12381 & inst_lookup0_cellmath__27[4]));
assign N12385 = !(N12381 & inst_lookup0_cellmath__27[4]);
assign N12404 = !(N1387 | N1388);
assign N12407 = !(inst_it2_lookup1_cellmath__53[0] | inst_it2_lookup1_cellmath__53[1]);
assign N12401 = !(N12397 & N12407);
assign N12411 = !(inst_lookup0_cellmath__27[3] | N12401);
assign N12408 = !((N1388 & N12397) | (N12407 & inst_lookup0_cellmath__27[2]));
assign N12368 = !(inst_it2_lookup1_cellmath__53[1] & inst_it2_lookup1_cellmath__53[0]);
assign N12376 = !((N12368 & N12397) | (N1388 & inst_lookup0_cellmath__27[2]));
assign N12396 = !((N12376 & N12386) | (N12408 & inst_lookup0_cellmath__27[3]));
assign N12419 = !((((!N12386) & inst_lookup0_cellmath__27[2]) & inst_lookup0_cellmath__27[4]) & N12404);
assign N12403 = !((N12396 & N12363) | (N12411 & inst_lookup0_cellmath__27[4]));
assign N12409 = !inst_lookup0_cellmath__27[5];
assign N12362 = !((N12419 & N12409) | (N12394 & inst_lookup0_cellmath__27[5]));
assign N12369 = !(inst_lookup0_cellmath__27[4] | N12373);
assign N12380 = !(N12369 | N12409);
assign N12417 = !((N12403 & N12409) | (N12385 & inst_lookup0_cellmath__27[5]));
assign N12364 = !((((!inst_lookup0_cellmath__27[3]) & N12404) & N12363) & N12397);
assign N12377 = !((N1388 & N1387) | (inst_it2_lookup1_cellmath__53[1] & inst_it2_lookup1_cellmath__53[0]));
assign N12395 = !((N1388 & N12397) | (N12377 & inst_lookup0_cellmath__27[2]));
assign N12410 = !((inst_it2_lookup1_cellmath__53[1] & N12397) | (N12404 & inst_lookup0_cellmath__27[2]));
assign N12400 = !((N12395 & N12386) | (N1388 & inst_lookup0_cellmath__27[3]));
assign N12414 = !(inst_lookup0_cellmath__27[3] | N12410);
assign N12375 = !(N12407 & inst_lookup0_cellmath__27[2]);
assign N12405 = !(N12397 | N12379);
assign N12387 = !(N12397 | inst_it2_lookup1_cellmath__53[1]);
assign N12371 = !((N12387 & N12386) | (N12375 & inst_lookup0_cellmath__27[3]));
assign N12384 = !(N12405 & inst_lookup0_cellmath__27[3]);
assign N12378 = !((N12371 & N12363) | (N12400 & inst_lookup0_cellmath__27[4]));
assign N12392 = !((N12384 & N12363) | (N12414 & inst_lookup0_cellmath__27[4]));
assign N12383 = !((N12378 & N12409) | (N12364 & inst_lookup0_cellmath__27[5]));
assign N12399 = !(inst_lookup0_cellmath__27[5] | N12392);
assign N12389 = !inst_lookup0_cellmath__27[6];
assign inst_cellmath__42[0] = !((N12362 & inst_lookup0_cellmath__27[6]) | (N12389 & N12383));
assign inst_lookup0_cellmath__29[1] = !((N12399 & N12389) | (N12380 & inst_lookup0_cellmath__27[6]));
assign inst_lookup0_cellmath__29[2] = !(N12389 | N12417);
assign inst_cellmath__43[0] = !inst_cellmath__42[0];
assign N2068 = !inst_cellmath__43[0];
assign N2045 = N2068 & inst_cellmath__9[0];
assign N2046 = N2068 & inst_cellmath__9[1];
assign N2047 = N2068 & inst_cellmath__9[2];
assign N2048 = N2068 & inst_cellmath__9[3];
assign N2049 = N2068 & inst_cellmath__9[4];
assign N2050 = N2068 & inst_cellmath__9[5];
assign N2051 = N2068 & inst_cellmath__9[6];
assign N2052 = N2068 & inst_cellmath__9[7];
assign N2053 = N2068 & inst_cellmath__9[8];
assign N2054 = N2068 & inst_cellmath__9[9];
assign N2055 = N2068 & inst_cellmath__9[10];
assign N2056 = N2068 & inst_cellmath__9[11];
assign N2057 = N2068 & inst_cellmath__9[12];
assign N2058 = N2068 & inst_cellmath__9[13];
assign N2059 = N2068 & inst_cellmath__9[14];
assign N2060 = N2068 & inst_cellmath__9[15];
assign N2061 = N2068 & inst_cellmath__9[16];
assign N2062 = N2068 & inst_cellmath__9[17];
assign N2063 = N2068 & inst_cellmath__9[18];
assign N2064 = N2068 & inst_cellmath__9[19];
assign N2065 = N2068 & inst_cellmath__9[20];
assign N2066 = N2068 & inst_it2_lookup1_cellmath__53[0];
assign N2067 = N2068 & inst_it2_lookup1_cellmath__53[1];
assign N12573 = !inst_lookup0_cellmath__29[1];
assign N2173 = !N12573;
assign N2150 = !(N2173 & inst_cellmath__9[0]);
assign N2151 = !(N2173 & inst_cellmath__9[1]);
assign N2152 = !(N2173 & inst_cellmath__9[2]);
assign N2153 = !(N2173 & inst_cellmath__9[3]);
assign N2154 = !(N2173 & inst_cellmath__9[4]);
assign N2155 = !(N2173 & inst_cellmath__9[5]);
assign N2156 = !(N2173 & inst_cellmath__9[6]);
assign N2157 = !(N2173 & inst_cellmath__9[7]);
assign N2158 = !(N2173 & inst_cellmath__9[8]);
assign N2159 = !(N2173 & inst_cellmath__9[9]);
assign N2160 = !(N2173 & inst_cellmath__9[10]);
assign N2161 = !(N2173 & inst_cellmath__9[11]);
assign N2162 = !(N2173 & inst_cellmath__9[12]);
assign N2163 = !(N2173 & inst_cellmath__9[13]);
assign N2164 = !(N2173 & inst_cellmath__9[14]);
assign N2165 = !(N2173 & inst_cellmath__9[15]);
assign N2166 = !(N2173 & inst_cellmath__9[16]);
assign N2167 = !(N2173 & inst_cellmath__9[17]);
assign N2168 = !(N2173 & inst_cellmath__9[18]);
assign N2169 = !(N2173 & inst_cellmath__9[19]);
assign N2170 = !(N2173 & inst_cellmath__9[20]);
assign N2171 = !(N2173 & inst_it2_lookup1_cellmath__53[0]);
assign N2172 = !(N2173 & inst_it2_lookup1_cellmath__53[1]);
assign N12658 = !inst_cellmath__11;
assign inst_cellmath__38__W0[2] = !N12658;
assign inst_cellmath__34[3] = (inst_cellmath__38__W0[2] & inst_cellmath__8[0]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[1]);
assign inst_cellmath__34[4] = (inst_cellmath__38__W0[2] & inst_cellmath__8[1]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[2]);
assign inst_cellmath__34[5] = (inst_cellmath__38__W0[2] & inst_cellmath__8[2]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[3]);
assign inst_cellmath__34[6] = (inst_cellmath__38__W0[2] & inst_cellmath__8[3]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[4]);
assign inst_cellmath__34[7] = (inst_cellmath__38__W0[2] & inst_cellmath__8[4]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[5]);
assign inst_cellmath__34[8] = (inst_cellmath__38__W0[2] & inst_cellmath__8[5]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[6]);
assign inst_cellmath__34[9] = (inst_cellmath__38__W0[2] & inst_cellmath__8[6]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[7]);
assign inst_cellmath__34[10] = (inst_cellmath__38__W0[2] & inst_cellmath__8[7]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[8]);
assign inst_cellmath__34[11] = (inst_cellmath__38__W0[2] & inst_cellmath__8[8]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[9]);
assign inst_cellmath__34[12] = (inst_cellmath__38__W0[2] & inst_cellmath__8[9]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[10]);
assign inst_cellmath__34[13] = (inst_cellmath__38__W0[2] & inst_cellmath__8[10]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[11]);
assign inst_cellmath__34[14] = (inst_cellmath__38__W0[2] & inst_cellmath__8[11]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[12]);
assign inst_cellmath__34[15] = (inst_cellmath__38__W0[2] & inst_cellmath__8[12]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[13]);
assign inst_cellmath__34[16] = (inst_cellmath__38__W0[2] & inst_cellmath__8[13]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[14]);
assign inst_cellmath__34[17] = (inst_cellmath__38__W0[2] & inst_cellmath__8[14]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[15]);
assign inst_cellmath__34[18] = (inst_cellmath__38__W0[2] & inst_cellmath__8[15]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[16]);
assign inst_cellmath__34[19] = (inst_cellmath__38__W0[2] & inst_cellmath__8[16]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[17]);
assign inst_cellmath__34[20] = (inst_cellmath__38__W0[2] & inst_cellmath__8[17]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[18]);
assign inst_cellmath__34[21] = (inst_cellmath__38__W0[2] & inst_cellmath__8[18]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[19]);
assign inst_cellmath__34[22] = (inst_cellmath__38__W0[2] & inst_cellmath__8[19]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[20]);
assign inst_cellmath__34[23] = (inst_cellmath__38__W0[2] & inst_cellmath__8[20]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[21]);
assign inst_cellmath__34[24] = (inst_cellmath__38__W0[2] & inst_cellmath__8[21]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[22]);
assign inst_cellmath__34[25] = (inst_cellmath__38__W0[2] & inst_cellmath__8[22]) | ((!inst_cellmath__38__W0[2]) & inst_cellmath__16[23]);
assign inst_it2_cellmath__60[4] = !inst_lookup0_cellmath__29[2];
assign N12797 = !inst_cellmath__17[1];
assign N12723 = !inst_cellmath__17[2];
assign N12744 = !inst_cellmath__17[3];
assign N12764 = !inst_cellmath__17[4];
assign N12785 = !inst_cellmath__17[5];
assign N12806 = !inst_cellmath__17[6];
assign N12732 = !inst_cellmath__17[7];
assign N12754 = !inst_cellmath__17[8];
assign N12774 = !inst_cellmath__17[9];
assign N12794 = !inst_cellmath__17[10];
assign N12720 = !inst_cellmath__17[11];
assign N12740 = !inst_cellmath__17[12];
assign N12761 = !inst_cellmath__17[13];
assign N12782 = !inst_cellmath__17[14];
assign N12803 = !inst_cellmath__17[15];
assign N12729 = !inst_cellmath__17[16];
assign N12751 = !inst_cellmath__17[17];
assign N12771 = !inst_cellmath__17[18];
assign N12791 = !inst_cellmath__17[19];
assign N12813 = !inst_cellmath__17[20];
assign N12738 = !inst_cellmath__17[21];
assign inst_cellmath__35[3] = !((N12797 & N12658) | (inst_cellmath__9[0] & inst_cellmath__11));
assign inst_cellmath__35[4] = !((N12723 & N12658) | (inst_cellmath__9[1] & inst_cellmath__11));
assign inst_cellmath__35[5] = !((N12744 & N12658) | (inst_cellmath__9[2] & inst_cellmath__11));
assign inst_cellmath__35[6] = !((N12764 & N12658) | (inst_cellmath__9[3] & inst_cellmath__11));
assign inst_cellmath__35[7] = !((N12785 & N12658) | (inst_cellmath__9[4] & inst_cellmath__11));
assign inst_cellmath__35[8] = !((N12806 & N12658) | (inst_cellmath__9[5] & inst_cellmath__11));
assign inst_cellmath__35[9] = !((N12732 & N12658) | (inst_cellmath__9[6] & inst_cellmath__11));
assign inst_cellmath__35[10] = !((N12754 & N12658) | (inst_cellmath__9[7] & inst_cellmath__11));
assign inst_cellmath__35[11] = !((N12774 & N12658) | (inst_cellmath__9[8] & inst_cellmath__11));
assign inst_cellmath__35[12] = !((N12794 & N12658) | (inst_cellmath__9[9] & inst_cellmath__11));
assign inst_cellmath__35[13] = !((N12720 & N12658) | (inst_cellmath__9[10] & inst_cellmath__11));
assign inst_cellmath__35[14] = !((N12740 & N12658) | (inst_cellmath__9[11] & inst_cellmath__11));
assign inst_cellmath__35[15] = !((N12761 & N12658) | (inst_cellmath__9[12] & inst_cellmath__11));
assign inst_cellmath__35[16] = !((N12782 & N12658) | (inst_cellmath__9[13] & inst_cellmath__11));
assign inst_cellmath__35[17] = !((N12803 & N12658) | (inst_cellmath__9[14] & inst_cellmath__11));
assign inst_cellmath__35[18] = !((N12729 & N12658) | (inst_cellmath__9[15] & inst_cellmath__11));
assign inst_cellmath__35[19] = !((N12751 & N12658) | (inst_cellmath__9[16] & inst_cellmath__11));
assign inst_cellmath__35[20] = !((N12771 & N12658) | (inst_cellmath__9[17] & inst_cellmath__11));
assign inst_cellmath__35[21] = !((N12791 & N12658) | (inst_cellmath__9[18] & inst_cellmath__11));
assign inst_cellmath__35[22] = !((N12813 & N12658) | (inst_cellmath__9[19] & inst_cellmath__11));
assign inst_cellmath__35[23] = !((N12738 & N12658) | (inst_cellmath__9[20] & inst_cellmath__11));
assign N12811 = !inst_cellmath__17[22];
assign inst_cellmath__35[24] = !((N12811 & N12658) | (inst_it2_lookup1_cellmath__53[0] & inst_cellmath__11));
assign N12736 = !inst_cellmath__17[23];
assign inst_cellmath__35[25] = !((N12736 & N12658) | (inst_it2_lookup1_cellmath__53[1] & inst_cellmath__11));
assign N12870 = !inst_it2_cellmath__60[4];
assign inst_it2_cellmath__61[3] = (!N2045) ^ N12870;
assign inst_cellmath__38__W1[2] = (!N2046) ^ N12870;
assign inst_cellmath__30[3] = (!N2047) ^ N12870;
assign inst_cellmath__30[4] = (!N2048) ^ N12870;
assign inst_cellmath__30[5] = (!N2049) ^ N12870;
assign inst_cellmath__30[6] = (!N2050) ^ N12870;
assign inst_cellmath__30[7] = (!N2051) ^ N12870;
assign inst_cellmath__30[8] = (!N2052) ^ N12870;
assign inst_cellmath__30[9] = (!N2053) ^ N12870;
assign inst_cellmath__30[10] = (!N2054) ^ N12870;
assign inst_cellmath__30[11] = (!N2055) ^ N12870;
assign inst_cellmath__30[12] = (!N2056) ^ N12870;
assign inst_cellmath__30[13] = (!N2057) ^ N12870;
assign inst_cellmath__30[14] = (!N2058) ^ N12870;
assign inst_cellmath__30[15] = (!N2059) ^ N12870;
assign inst_cellmath__30[16] = (!N2060) ^ N12870;
assign inst_cellmath__30[17] = (!N2061) ^ N12870;
assign inst_cellmath__30[18] = (!N2062) ^ N12870;
assign inst_cellmath__30[19] = (!N2063) ^ N12870;
assign inst_cellmath__30[20] = (!N2064) ^ N12870;
assign inst_cellmath__30[21] = (!N2065) ^ N12870;
assign inst_cellmath__30[22] = (!N2066) ^ N12870;
assign inst_cellmath__30[23] = (!N2067) ^ N12870;
assign inst_cellmath__30[24] = (!N2068) ^ N12870;
assign {inst_cellmath__38__W0[3], inst_cellmath__38__W1[3]} = {1'B0, inst_cellmath__34[3]} + {1'B0, inst_cellmath__35[3]} + {1'B0, inst_cellmath__30[3]};
assign {inst_cellmath__38__W0[4], inst_cellmath__38__W1[4]} = {1'B0, inst_cellmath__34[4]} + {1'B0, inst_cellmath__35[4]} + {1'B0, inst_cellmath__30[4]};
assign {inst_cellmath__38__W0[5], inst_cellmath__38__W1[5]} = {1'B0, inst_cellmath__34[5]} + {1'B0, inst_cellmath__35[5]} + {1'B0, inst_cellmath__30[5]};
assign {inst_cellmath__38__W0[6], inst_cellmath__38__W1[6]} = {1'B0, inst_cellmath__34[6]} + {1'B0, inst_cellmath__35[6]} + {1'B0, inst_cellmath__30[6]};
assign {inst_cellmath__38__W0[7], inst_cellmath__38__W1[7]} = {1'B0, inst_cellmath__34[7]} + {1'B0, inst_cellmath__35[7]} + {1'B0, inst_cellmath__30[7]};
assign {inst_cellmath__38__W0[8], inst_cellmath__38__W1[8]} = {1'B0, inst_cellmath__34[8]} + {1'B0, inst_cellmath__35[8]} + {1'B0, inst_cellmath__30[8]};
assign {inst_cellmath__38__W0[9], inst_cellmath__38__W1[9]} = {1'B0, inst_cellmath__34[9]} + {1'B0, inst_cellmath__35[9]} + {1'B0, inst_cellmath__30[9]};
assign {inst_cellmath__38__W0[10], inst_cellmath__38__W1[10]} = {1'B0, inst_cellmath__34[10]} + {1'B0, inst_cellmath__35[10]} + {1'B0, inst_cellmath__30[10]};
assign {inst_cellmath__38__W0[11], inst_cellmath__38__W1[11]} = {1'B0, inst_cellmath__34[11]} + {1'B0, inst_cellmath__35[11]} + {1'B0, inst_cellmath__30[11]};
assign {inst_cellmath__38__W0[12], inst_cellmath__38__W1[12]} = {1'B0, inst_cellmath__34[12]} + {1'B0, inst_cellmath__35[12]} + {1'B0, inst_cellmath__30[12]};
assign {inst_cellmath__38__W0[13], inst_cellmath__38__W1[13]} = {1'B0, inst_cellmath__34[13]} + {1'B0, inst_cellmath__35[13]} + {1'B0, inst_cellmath__30[13]};
assign {inst_cellmath__38__W0[14], inst_cellmath__38__W1[14]} = {1'B0, inst_cellmath__34[14]} + {1'B0, inst_cellmath__35[14]} + {1'B0, inst_cellmath__30[14]};
assign {inst_cellmath__38__W0[15], inst_cellmath__38__W1[15]} = {1'B0, inst_cellmath__34[15]} + {1'B0, inst_cellmath__35[15]} + {1'B0, inst_cellmath__30[15]};
assign {inst_cellmath__38__W0[16], inst_cellmath__38__W1[16]} = {1'B0, inst_cellmath__34[16]} + {1'B0, inst_cellmath__35[16]} + {1'B0, inst_cellmath__30[16]};
assign {inst_cellmath__38__W0[17], inst_cellmath__38__W1[17]} = {1'B0, inst_cellmath__34[17]} + {1'B0, inst_cellmath__35[17]} + {1'B0, inst_cellmath__30[17]};
assign {inst_cellmath__38__W0[18], inst_cellmath__38__W1[18]} = {1'B0, inst_cellmath__34[18]} + {1'B0, inst_cellmath__35[18]} + {1'B0, inst_cellmath__30[18]};
assign {inst_cellmath__38__W0[19], inst_cellmath__38__W1[19]} = {1'B0, inst_cellmath__34[19]} + {1'B0, inst_cellmath__35[19]} + {1'B0, inst_cellmath__30[19]};
assign {inst_cellmath__38__W0[20], inst_cellmath__38__W1[20]} = {1'B0, inst_cellmath__34[20]} + {1'B0, inst_cellmath__35[20]} + {1'B0, inst_cellmath__30[20]};
assign {inst_cellmath__38__W0[21], inst_cellmath__38__W1[21]} = {1'B0, inst_cellmath__34[21]} + {1'B0, inst_cellmath__35[21]} + {1'B0, inst_cellmath__30[21]};
assign {inst_cellmath__38__W0[22], inst_cellmath__38__W1[22]} = {1'B0, inst_cellmath__34[22]} + {1'B0, inst_cellmath__35[22]} + {1'B0, inst_cellmath__30[22]};
assign {inst_cellmath__38__W0[23], inst_cellmath__38__W1[23]} = {1'B0, inst_cellmath__34[23]} + {1'B0, inst_cellmath__35[23]} + {1'B0, inst_cellmath__30[23]};
assign {inst_cellmath__38__W0[24], inst_cellmath__38__W1[24]} = {1'B0, inst_cellmath__34[24]} + {1'B0, inst_cellmath__35[24]} + {1'B0, inst_cellmath__30[24]};
assign {N12983, inst_cellmath__38__W1[25]} = {1'B0, inst_cellmath__34[25]} + {1'B0, inst_cellmath__35[25]} + {1'B0, inst_it2_cellmath__60[4]};
assign inst_cellmath__31[1] = !N12870;
assign inst_cellmath__31[2] = !((N2150 & N12870) | ((!N2150) & inst_cellmath__31[1]));
assign inst_cellmath__31[3] = !((N2151 & N12870) | ((!N2151) & inst_cellmath__31[1]));
assign inst_cellmath__31[4] = !((N2152 & N12870) | ((!N2152) & inst_cellmath__31[1]));
assign inst_cellmath__31[5] = !((N2153 & N12870) | ((!N2153) & inst_cellmath__31[1]));
assign inst_cellmath__31[6] = !((N2154 & N12870) | ((!N2154) & inst_cellmath__31[1]));
assign inst_cellmath__31[7] = !((N2155 & N12870) | ((!N2155) & inst_cellmath__31[1]));
assign inst_cellmath__31[8] = !((N2156 & N12870) | ((!N2156) & inst_cellmath__31[1]));
assign inst_cellmath__31[9] = !((N2157 & N12870) | ((!N2157) & inst_cellmath__31[1]));
assign inst_cellmath__31[10] = !((N2158 & N12870) | ((!N2158) & inst_cellmath__31[1]));
assign inst_cellmath__31[11] = !((N2159 & N12870) | ((!N2159) & inst_cellmath__31[1]));
assign inst_cellmath__31[12] = !((N2160 & N12870) | ((!N2160) & inst_cellmath__31[1]));
assign inst_cellmath__31[13] = !((N2161 & N12870) | ((!N2161) & inst_cellmath__31[1]));
assign inst_cellmath__31[14] = !((N2162 & N12870) | ((!N2162) & inst_cellmath__31[1]));
assign inst_cellmath__31[15] = !((N2163 & N12870) | ((!N2163) & inst_cellmath__31[1]));
assign inst_cellmath__31[16] = !((N2164 & N12870) | ((!N2164) & inst_cellmath__31[1]));
assign inst_cellmath__31[17] = !((N2165 & N12870) | ((!N2165) & inst_cellmath__31[1]));
assign inst_cellmath__31[18] = !((N2166 & N12870) | ((!N2166) & inst_cellmath__31[1]));
assign inst_cellmath__31[19] = !((N2167 & N12870) | ((!N2167) & inst_cellmath__31[1]));
assign inst_cellmath__31[20] = !((N2168 & N12870) | ((!N2168) & inst_cellmath__31[1]));
assign inst_cellmath__31[21] = !((N2169 & N12870) | ((!N2169) & inst_cellmath__31[1]));
assign inst_cellmath__31[22] = !((N2170 & N12870) | ((!N2170) & inst_cellmath__31[1]));
assign inst_cellmath__31[23] = !((N2171 & N12870) | ((!N2171) & inst_cellmath__31[1]));
assign inst_cellmath__31[24] = !((N2172 & N12870) | ((!N2172) & inst_cellmath__31[1]));
assign inst_cellmath__31[25] = !((N2173 & inst_cellmath__31[1]) | ((!N2173) & N12870));
assign N28016 = !inst_it2_cellmath__60[4];
assign inst_it2_cellmath__60[3] = !N28016;
assign {inst_it2_cellmath__60[5], inst_it2_cellmath__61[4]} = {1'B0, inst_cellmath__38__W1[2]} + {1'B0, inst_cellmath__31[2]};
assign {inst_it2_cellmath__60[6], inst_it2_cellmath__61[5]} = {1'B0, inst_cellmath__38__W1[3]} + {1'B0, inst_cellmath__38__W0[2]} + {1'B0, inst_cellmath__31[3]};
assign {inst_it2_cellmath__60[7], inst_it2_cellmath__61[6]} = {1'B0, inst_cellmath__38__W1[4]} + {1'B0, inst_cellmath__38__W0[3]} + {1'B0, inst_cellmath__31[4]};
assign {inst_it2_cellmath__60[8], inst_it2_cellmath__61[7]} = {1'B0, inst_cellmath__38__W1[5]} + {1'B0, inst_cellmath__38__W0[4]} + {1'B0, inst_cellmath__31[5]};
assign {inst_it2_cellmath__60[9], inst_it2_cellmath__61[8]} = {1'B0, inst_cellmath__38__W1[6]} + {1'B0, inst_cellmath__38__W0[5]} + {1'B0, inst_cellmath__31[6]};
assign {inst_it2_cellmath__60[10], inst_it2_cellmath__61[9]} = {1'B0, inst_cellmath__38__W1[7]} + {1'B0, inst_cellmath__38__W0[6]} + {1'B0, inst_cellmath__31[7]};
assign {inst_it2_cellmath__60[11], inst_it2_cellmath__61[10]} = {1'B0, inst_cellmath__38__W1[8]} + {1'B0, inst_cellmath__38__W0[7]} + {1'B0, inst_cellmath__31[8]};
assign {inst_it2_cellmath__60[12], inst_it2_cellmath__61[11]} = {1'B0, inst_cellmath__38__W1[9]} + {1'B0, inst_cellmath__38__W0[8]} + {1'B0, inst_cellmath__31[9]};
assign {inst_it2_cellmath__60[13], inst_it2_cellmath__61[12]} = {1'B0, inst_cellmath__38__W1[10]} + {1'B0, inst_cellmath__38__W0[9]} + {1'B0, inst_cellmath__31[10]};
assign {inst_it2_cellmath__60[14], inst_it2_cellmath__61[13]} = {1'B0, inst_cellmath__38__W1[11]} + {1'B0, inst_cellmath__38__W0[10]} + {1'B0, inst_cellmath__31[11]};
assign {inst_it2_cellmath__60[15], inst_it2_cellmath__61[14]} = {1'B0, inst_cellmath__38__W1[12]} + {1'B0, inst_cellmath__38__W0[11]} + {1'B0, inst_cellmath__31[12]};
assign {inst_it2_cellmath__60[16], inst_it2_cellmath__61[15]} = {1'B0, inst_cellmath__38__W1[13]} + {1'B0, inst_cellmath__38__W0[12]} + {1'B0, inst_cellmath__31[13]};
assign {inst_it2_cellmath__60[17], inst_it2_cellmath__61[16]} = {1'B0, inst_cellmath__38__W1[14]} + {1'B0, inst_cellmath__38__W0[13]} + {1'B0, inst_cellmath__31[14]};
assign {inst_it2_cellmath__60[18], inst_it2_cellmath__61[17]} = {1'B0, inst_cellmath__38__W1[15]} + {1'B0, inst_cellmath__38__W0[14]} + {1'B0, inst_cellmath__31[15]};
assign {inst_it2_cellmath__60[19], inst_it2_cellmath__61[18]} = {1'B0, inst_cellmath__38__W1[16]} + {1'B0, inst_cellmath__38__W0[15]} + {1'B0, inst_cellmath__31[16]};
assign {inst_it2_cellmath__60[20], inst_it2_cellmath__61[19]} = {1'B0, inst_cellmath__38__W1[17]} + {1'B0, inst_cellmath__38__W0[16]} + {1'B0, inst_cellmath__31[17]};
assign {inst_it2_cellmath__60[21], inst_it2_cellmath__61[20]} = {1'B0, inst_cellmath__38__W1[18]} + {1'B0, inst_cellmath__38__W0[17]} + {1'B0, inst_cellmath__31[18]};
assign {inst_it2_cellmath__60[22], inst_it2_cellmath__61[21]} = {1'B0, inst_cellmath__38__W1[19]} + {1'B0, inst_cellmath__38__W0[18]} + {1'B0, inst_cellmath__31[19]};
assign {inst_it2_cellmath__60[23], inst_it2_cellmath__61[22]} = {1'B0, inst_cellmath__38__W1[20]} + {1'B0, inst_cellmath__38__W0[19]} + {1'B0, inst_cellmath__31[20]};
assign {inst_it2_cellmath__60[24], inst_it2_cellmath__61[23]} = {1'B0, inst_cellmath__38__W1[21]} + {1'B0, inst_cellmath__38__W0[20]} + {1'B0, inst_cellmath__31[21]};
assign {inst_it2_cellmath__60[25], inst_it2_cellmath__61[24]} = {1'B0, inst_cellmath__38__W1[22]} + {1'B0, inst_cellmath__38__W0[21]} + {1'B0, inst_cellmath__31[22]};
assign {inst_cellmath__39__W0[23], inst_it2_cellmath__61[25]} = {1'B0, inst_cellmath__38__W1[23]} + {1'B0, inst_cellmath__38__W0[22]} + {1'B0, inst_cellmath__31[23]};
assign {inst_cellmath__39__W0[24], inst_cellmath__39__W1[24]} = {1'B0, inst_cellmath__38__W1[24]} + {1'B0, inst_cellmath__38__W0[23]} + {1'B0, inst_cellmath__31[24]};
assign {N13206, inst_cellmath__39__W1[25]} = {1'B0, inst_cellmath__38__W1[25]} + {1'B0, inst_cellmath__38__W0[24]} + {1'B0, inst_cellmath__31[25]};
assign {N13380, inst_it2_lookup1_cellmath__53[2]} = {1'B0, inst_it2_cellmath__60[23]} + {1'B0, inst_it2_cellmath__61[23]};
assign {N13376, inst_it2_lookup1_cellmath__53[3]} = {1'B0, inst_it2_cellmath__60[24]} + {1'B0, inst_it2_cellmath__61[24]} + {1'B0, N13380};
assign {N13387, inst_it2_lookup1_cellmath__53[4]} = {1'B0, inst_it2_cellmath__60[25]} + {1'B0, inst_it2_cellmath__61[25]} + {1'B0, N13376};
assign {N13373, inst_it2_lookup1_cellmath__53[5]} = {1'B0, inst_cellmath__39__W0[23]} + {1'B0, inst_cellmath__39__W1[24]} + {1'B0, N13387};
assign {N13384, inst_it2_lookup1_cellmath__53[6]} = {1'B0, inst_cellmath__39__W1[25]} + {1'B0, inst_cellmath__39__W0[24]} + {1'B0, N13373};
assign N13436 = !inst_it2_lookup1_cellmath__53[2];
assign N13425 = !inst_it2_lookup1_cellmath__53[3];
assign N13420 = !(N13425 | N13436);
assign N13457 = !(N13436 | N1388);
assign N13405 = !((inst_it2_lookup1_cellmath__53[1] & N13436) | (N12379 & inst_it2_lookup1_cellmath__53[2]));
assign N13460 = !((N13405 & N13425) | (N13457 & inst_it2_lookup1_cellmath__53[3]));
assign N13404 = !(inst_it2_lookup1_cellmath__53[1] & inst_it2_lookup1_cellmath__53[2]);
assign N13412 = !(N13425 | N13404);
assign N13402 = !inst_it2_lookup1_cellmath__53[4];
assign N13433 = !((N13460 & N13402) | (N13420 & inst_it2_lookup1_cellmath__53[4]));
assign N13424 = !(N13420 & inst_it2_lookup1_cellmath__53[4]);
assign N13440 = !(N13436 & N12407);
assign N13450 = !(inst_it2_lookup1_cellmath__53[3] | N13440);
assign N13447 = !((N1388 & N13436) | (N12407 & inst_it2_lookup1_cellmath__53[2]));
assign N13415 = !((N12368 & N13436) | (N1388 & inst_it2_lookup1_cellmath__53[2]));
assign N13435 = !((N13415 & N13425) | (N13447 & inst_it2_lookup1_cellmath__53[3]));
assign N13458 = !((((!N13425) & N12404) & inst_it2_lookup1_cellmath__53[4]) & inst_it2_lookup1_cellmath__53[2]);
assign N13442 = !((N13435 & N13402) | (N13450 & inst_it2_lookup1_cellmath__53[4]));
assign N13448 = !inst_it2_lookup1_cellmath__53[5];
assign N13401 = !((N13458 & N13448) | (N13433 & inst_it2_lookup1_cellmath__53[5]));
assign N13408 = !(inst_it2_lookup1_cellmath__53[4] | N13412);
assign N13419 = !(N13408 | N13448);
assign N13456 = !((N13442 & N13448) | (N13424 & inst_it2_lookup1_cellmath__53[5]));
assign N13403 = !((((!inst_it2_lookup1_cellmath__53[3]) & N12404) & N13402) & N13436);
assign N13434 = !((N1388 & N13436) | (N12377 & inst_it2_lookup1_cellmath__53[2]));
assign N13449 = !((inst_it2_lookup1_cellmath__53[1] & N13436) | (N12404 & inst_it2_lookup1_cellmath__53[2]));
assign N13439 = !((N13434 & N13425) | (N1388 & inst_it2_lookup1_cellmath__53[3]));
assign N13453 = !(inst_it2_lookup1_cellmath__53[3] | N13449);
assign N13414 = !(N12407 & inst_it2_lookup1_cellmath__53[2]);
assign N13444 = !(N13436 | N12379);
assign N13426 = !(N13436 | inst_it2_lookup1_cellmath__53[1]);
assign N13410 = !((N13426 & N13425) | (N13414 & inst_it2_lookup1_cellmath__53[3]));
assign N13423 = !(N13444 & inst_it2_lookup1_cellmath__53[3]);
assign N13417 = !((N13410 & N13402) | (N13439 & inst_it2_lookup1_cellmath__53[4]));
assign N13431 = !((N13423 & N13402) | (N13453 & inst_it2_lookup1_cellmath__53[4]));
assign N13422 = !((N13417 & N13448) | (N13403 & inst_it2_lookup1_cellmath__53[5]));
assign N13438 = !(inst_it2_lookup1_cellmath__53[5] | N13431);
assign N13428 = !inst_it2_lookup1_cellmath__53[6];
assign inst_cellmath__40[0] = !((N13401 & inst_it2_lookup1_cellmath__53[6]) | (N13428 & N13422));
assign inst_it2_lookup1_cellmath__55[1] = !((N13438 & N13428) | (N13419 & inst_it2_lookup1_cellmath__53[6]));
assign inst_it2_lookup1_cellmath__55[2] = !(N13428 | N13456);
assign inst_cellmath__41[0] = !inst_cellmath__40[0];
assign N2224 = !inst_cellmath__41[0];
assign N2201 = N2224 & inst_cellmath__9[0];
assign N2202 = N2224 & inst_cellmath__9[1];
assign N2203 = N2224 & inst_cellmath__9[2];
assign N2204 = N2224 & inst_cellmath__9[3];
assign N2205 = N2224 & inst_cellmath__9[4];
assign N2206 = N2224 & inst_cellmath__9[5];
assign N2207 = N2224 & inst_cellmath__9[6];
assign N2208 = N2224 & inst_cellmath__9[7];
assign N2209 = N2224 & inst_cellmath__9[8];
assign N2210 = N2224 & inst_cellmath__9[9];
assign N2211 = N2224 & inst_cellmath__9[10];
assign N2212 = N2224 & inst_cellmath__9[11];
assign N2213 = N2224 & inst_cellmath__9[12];
assign N2214 = N2224 & inst_cellmath__9[13];
assign N2215 = N2224 & inst_cellmath__9[14];
assign N2216 = N2224 & inst_cellmath__9[15];
assign N2217 = N2224 & inst_cellmath__9[16];
assign N2218 = N2224 & inst_cellmath__9[17];
assign N2219 = N2224 & inst_cellmath__9[18];
assign N2220 = N2224 & inst_cellmath__9[19];
assign N2221 = N2224 & inst_cellmath__9[20];
assign N2222 = N2224 & inst_it2_lookup1_cellmath__53[0];
assign N2223 = N2224 & inst_it2_lookup1_cellmath__53[1];
assign N13614 = !inst_it2_lookup1_cellmath__55[1];
assign N2277 = !N13614;
assign N2254 = !(N2277 & inst_cellmath__9[0]);
assign N2255 = !(N2277 & inst_cellmath__9[1]);
assign N2256 = !(N2277 & inst_cellmath__9[2]);
assign N2257 = !(N2277 & inst_cellmath__9[3]);
assign N2258 = !(N2277 & inst_cellmath__9[4]);
assign N2259 = !(N2277 & inst_cellmath__9[5]);
assign N2260 = !(N2277 & inst_cellmath__9[6]);
assign N2261 = !(N2277 & inst_cellmath__9[7]);
assign N2262 = !(N2277 & inst_cellmath__9[8]);
assign N2263 = !(N2277 & inst_cellmath__9[9]);
assign N2264 = !(N2277 & inst_cellmath__9[10]);
assign N2265 = !(N2277 & inst_cellmath__9[11]);
assign N2266 = !(N2277 & inst_cellmath__9[12]);
assign N2267 = !(N2277 & inst_cellmath__9[13]);
assign N2268 = !(N2277 & inst_cellmath__9[14]);
assign N2269 = !(N2277 & inst_cellmath__9[15]);
assign N2270 = !(N2277 & inst_cellmath__9[16]);
assign N2271 = !(N2277 & inst_cellmath__9[17]);
assign N2272 = !(N2277 & inst_cellmath__9[18]);
assign N2273 = !(N2277 & inst_cellmath__9[19]);
assign N2274 = !(N2277 & inst_cellmath__9[20]);
assign N2275 = !(N2277 & inst_it2_lookup1_cellmath__53[0]);
assign N2276 = !(N2277 & inst_it2_lookup1_cellmath__53[1]);
reg inst_cellmath__112_0_0__I168_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_0__I168_QOUT <= N1751;
assign inst_cellmath__112[0] = inst_cellmath__112_0_0__I168_QOUT;
reg inst_cellmath__112_0_1__I169_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_1__I169_QOUT <= N1752;
assign inst_cellmath__112[1] = inst_cellmath__112_0_1__I169_QOUT;
reg inst_cellmath__112_0_2__I170_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_2__I170_QOUT <= N1753;
assign inst_cellmath__112[2] = inst_cellmath__112_0_2__I170_QOUT;
reg inst_cellmath__112_0_3__I171_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_3__I171_QOUT <= N1754;
assign inst_cellmath__112[3] = inst_cellmath__112_0_3__I171_QOUT;
reg inst_cellmath__112_0_4__I172_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_4__I172_QOUT <= N1755;
assign inst_cellmath__112[4] = inst_cellmath__112_0_4__I172_QOUT;
reg inst_cellmath__112_0_5__I173_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_5__I173_QOUT <= N1756;
assign inst_cellmath__112[5] = inst_cellmath__112_0_5__I173_QOUT;
reg inst_cellmath__112_0_6__I174_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_6__I174_QOUT <= N1757;
assign inst_cellmath__112[6] = inst_cellmath__112_0_6__I174_QOUT;
reg inst_cellmath__112_0_7__I175_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_7__I175_QOUT <= N1758;
assign inst_cellmath__112[7] = inst_cellmath__112_0_7__I175_QOUT;
reg inst_cellmath__112_0_8__I176_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_8__I176_QOUT <= N1759;
assign inst_cellmath__112[8] = inst_cellmath__112_0_8__I176_QOUT;
reg inst_cellmath__112_0_9__I177_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_9__I177_QOUT <= N1760;
assign inst_cellmath__112[9] = inst_cellmath__112_0_9__I177_QOUT;
reg inst_cellmath__112_0_10__I178_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_10__I178_QOUT <= N1761;
assign inst_cellmath__112[10] = inst_cellmath__112_0_10__I178_QOUT;
reg inst_cellmath__112_0_11__I179_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_11__I179_QOUT <= N1762;
assign inst_cellmath__112[11] = inst_cellmath__112_0_11__I179_QOUT;
reg inst_cellmath__112_0_12__I180_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_12__I180_QOUT <= N1763;
assign inst_cellmath__112[12] = inst_cellmath__112_0_12__I180_QOUT;
reg inst_cellmath__112_0_13__I181_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_13__I181_QOUT <= N1764;
assign inst_cellmath__112[13] = inst_cellmath__112_0_13__I181_QOUT;
reg inst_cellmath__112_0_14__I182_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_14__I182_QOUT <= N1765;
assign inst_cellmath__112[14] = inst_cellmath__112_0_14__I182_QOUT;
reg inst_cellmath__112_0_15__I183_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_15__I183_QOUT <= N1766;
assign inst_cellmath__112[15] = inst_cellmath__112_0_15__I183_QOUT;
reg inst_cellmath__112_0_16__I184_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_16__I184_QOUT <= N1767;
assign inst_cellmath__112[16] = inst_cellmath__112_0_16__I184_QOUT;
reg inst_cellmath__112_0_17__I185_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_17__I185_QOUT <= N1768;
assign inst_cellmath__112[17] = inst_cellmath__112_0_17__I185_QOUT;
reg inst_cellmath__112_0_18__I186_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_18__I186_QOUT <= N1769;
assign inst_cellmath__112[18] = inst_cellmath__112_0_18__I186_QOUT;
reg inst_cellmath__112_0_19__I187_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_19__I187_QOUT <= N1770;
assign inst_cellmath__112[19] = inst_cellmath__112_0_19__I187_QOUT;
reg inst_cellmath__112_0_20__I188_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_20__I188_QOUT <= N1771;
assign inst_cellmath__112[20] = inst_cellmath__112_0_20__I188_QOUT;
reg inst_cellmath__112_0_21__I189_QOUT;
always @ (posedge clk)
	inst_cellmath__112_0_21__I189_QOUT <= N1772;
assign inst_cellmath__112[21] = inst_cellmath__112_0_21__I189_QOUT;
assign {N13719, inst_cellmath__120[1]} = {1'B0, inst_cellmath__16[1]} + {1'B0, inst_cellmath__17[1]};
assign {N13661, inst_cellmath__120[2]} = {1'B0, inst_cellmath__16[2]} + {1'B0, inst_cellmath__17[2]} + {1'B0, N13719};
assign {N13705, inst_cellmath__120[3]} = {1'B0, inst_cellmath__16[3]} + {1'B0, inst_cellmath__17[3]} + {1'B0, N13661};
assign {N13753, inst_cellmath__120[4]} = {1'B0, inst_cellmath__16[4]} + {1'B0, inst_cellmath__17[4]} + {1'B0, N13705};
assign {N13692, inst_cellmath__120[5]} = {1'B0, inst_cellmath__16[5]} + {1'B0, inst_cellmath__17[5]} + {1'B0, N13753};
assign {N13738, inst_cellmath__120[6]} = {1'B0, inst_cellmath__16[6]} + {1'B0, inst_cellmath__17[6]} + {1'B0, N13692};
assign {N13680, inst_cellmath__120[7]} = {1'B0, inst_cellmath__16[7]} + {1'B0, inst_cellmath__17[7]} + {1'B0, N13738};
assign {N13725, inst_cellmath__120[8]} = {1'B0, inst_cellmath__16[8]} + {1'B0, inst_cellmath__17[8]} + {1'B0, N13680};
assign {N13667, inst_cellmath__120[9]} = {1'B0, inst_cellmath__16[9]} + {1'B0, inst_cellmath__17[9]} + {1'B0, N13725};
assign {N13712, inst_cellmath__120[10]} = {1'B0, inst_cellmath__16[10]} + {1'B0, inst_cellmath__17[10]} + {1'B0, N13667};
assign {N13758, inst_cellmath__120[11]} = {1'B0, inst_cellmath__16[11]} + {1'B0, inst_cellmath__17[11]} + {1'B0, N13712};
assign {N13697, inst_cellmath__120[12]} = {1'B0, inst_cellmath__16[12]} + {1'B0, inst_cellmath__17[12]} + {1'B0, N13758};
assign {N13745, inst_cellmath__120[13]} = {1'B0, inst_cellmath__16[13]} + {1'B0, inst_cellmath__17[13]} + {1'B0, N13697};
assign {N13685, inst_cellmath__120[14]} = {1'B0, inst_cellmath__16[14]} + {1'B0, inst_cellmath__17[14]} + {1'B0, N13745};
assign {N13730, inst_cellmath__120[15]} = {1'B0, inst_cellmath__16[15]} + {1'B0, inst_cellmath__17[15]} + {1'B0, N13685};
assign {N13673, inst_cellmath__120[16]} = {1'B0, inst_cellmath__16[16]} + {1'B0, inst_cellmath__17[16]} + {1'B0, N13730};
assign {N13716, inst_cellmath__120[17]} = {1'B0, inst_cellmath__16[17]} + {1'B0, inst_cellmath__17[17]} + {1'B0, N13673};
assign {N13658, inst_cellmath__120[18]} = {1'B0, inst_cellmath__16[18]} + {1'B0, inst_cellmath__17[18]} + {1'B0, N13716};
assign {N13704, inst_cellmath__120[19]} = {1'B0, inst_cellmath__16[19]} + {1'B0, inst_cellmath__17[19]} + {1'B0, N13658};
assign {N13750, inst_cellmath__120[20]} = {1'B0, inst_cellmath__16[20]} + {1'B0, inst_cellmath__17[20]} + {1'B0, N13704};
assign {N13689, inst_cellmath__120[21]} = {1'B0, inst_cellmath__17[21]} + {1'B0, inst_cellmath__16[21]} + {1'B0, N13750};
assign {N13737, inst_cellmath__120[22]} = {1'B0, inst_cellmath__17[22]} + {1'B0, inst_cellmath__16[22]} + {1'B0, N13689};
assign {N13677, inst_cellmath__120[23]} = {1'B0, inst_cellmath__17[23]} + {1'B0, inst_cellmath__16[23]} + {1'B0, N13737};
assign {N13722, inst_cellmath__120[24]} = {1'B0, inst_cellmath__17[24]} + {1'B0, inst_cellmath__16[24]} + {1'B0, N13677};
assign {N13665, inst_cellmath__120[25]} = {1'B0, inst_cellmath__17[25]} + {1'B0, inst_cellmath__16[25]} + {1'B0, N13722};
reg inst_cellmath__44_0_0__I191_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_0__I191_QOUT <= inst_cellmath__40[0];
assign inst_cellmath__44[0] = inst_cellmath__44_0_0__I191_QOUT;
reg inst_cellmath__44_0_1__I192_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_1__I192_QOUT <= inst_cellmath__40[1];
assign inst_cellmath__44[1] = inst_cellmath__44_0_1__I192_QOUT;
reg inst_cellmath__44_0_2__I193_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_2__I193_QOUT <= inst_cellmath__40[2];
assign inst_cellmath__44[2] = inst_cellmath__44_0_2__I193_QOUT;
reg inst_cellmath__44_0_3__I194_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_3__I194_QOUT <= inst_cellmath__40[3];
assign inst_cellmath__44[3] = inst_cellmath__44_0_3__I194_QOUT;
reg inst_cellmath__44_0_4__I195_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_4__I195_QOUT <= inst_cellmath__40[4];
assign inst_cellmath__44[4] = inst_cellmath__44_0_4__I195_QOUT;
reg inst_cellmath__44_0_5__I196_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_5__I196_QOUT <= inst_cellmath__40[5];
assign inst_cellmath__44[5] = inst_cellmath__44_0_5__I196_QOUT;
reg inst_cellmath__44_0_6__I197_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_6__I197_QOUT <= inst_cellmath__40[6];
assign inst_cellmath__44[6] = inst_cellmath__44_0_6__I197_QOUT;
reg inst_cellmath__44_0_7__I198_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_7__I198_QOUT <= inst_cellmath__40[7];
assign inst_cellmath__44[7] = inst_cellmath__44_0_7__I198_QOUT;
reg inst_cellmath__44_0_8__I199_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_8__I199_QOUT <= inst_cellmath__40[8];
assign inst_cellmath__44[8] = inst_cellmath__44_0_8__I199_QOUT;
reg inst_cellmath__44_0_9__I200_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_9__I200_QOUT <= inst_cellmath__40[9];
assign inst_cellmath__44[9] = inst_cellmath__44_0_9__I200_QOUT;
reg inst_cellmath__44_0_10__I201_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_10__I201_QOUT <= inst_cellmath__40[10];
assign inst_cellmath__44[10] = inst_cellmath__44_0_10__I201_QOUT;
reg inst_cellmath__44_0_11__I202_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_11__I202_QOUT <= inst_cellmath__40[11];
assign inst_cellmath__44[11] = inst_cellmath__44_0_11__I202_QOUT;
reg inst_cellmath__44_0_12__I203_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_12__I203_QOUT <= inst_cellmath__40[12];
assign inst_cellmath__44[12] = inst_cellmath__44_0_12__I203_QOUT;
reg inst_cellmath__44_0_13__I204_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_13__I204_QOUT <= inst_cellmath__40[13];
assign inst_cellmath__44[13] = inst_cellmath__44_0_13__I204_QOUT;
reg inst_cellmath__44_0_14__I205_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_14__I205_QOUT <= inst_cellmath__40[14];
assign inst_cellmath__44[14] = inst_cellmath__44_0_14__I205_QOUT;
reg inst_cellmath__44_0_15__I206_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_15__I206_QOUT <= inst_cellmath__40[15];
assign inst_cellmath__44[15] = inst_cellmath__44_0_15__I206_QOUT;
reg inst_cellmath__44_0_16__I207_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_16__I207_QOUT <= inst_cellmath__40[16];
assign inst_cellmath__44[16] = inst_cellmath__44_0_16__I207_QOUT;
reg inst_cellmath__44_0_17__I208_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_17__I208_QOUT <= inst_cellmath__40[17];
assign inst_cellmath__44[17] = inst_cellmath__44_0_17__I208_QOUT;
reg inst_cellmath__44_0_18__I209_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_18__I209_QOUT <= inst_cellmath__40[18];
assign inst_cellmath__44[18] = inst_cellmath__44_0_18__I209_QOUT;
reg inst_cellmath__44_0_19__I210_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_19__I210_QOUT <= inst_cellmath__40[19];
assign inst_cellmath__44[19] = inst_cellmath__44_0_19__I210_QOUT;
reg inst_cellmath__44_0_20__I211_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_20__I211_QOUT <= inst_cellmath__40[20];
assign inst_cellmath__44[20] = inst_cellmath__44_0_20__I211_QOUT;
reg inst_cellmath__44_0_21__I212_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_21__I212_QOUT <= inst_cellmath__40[21];
assign inst_cellmath__44[21] = inst_cellmath__44_0_21__I212_QOUT;
reg inst_cellmath__44_0_22__I213_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_22__I213_QOUT <= inst_cellmath__40[22];
assign inst_cellmath__44[22] = inst_cellmath__44_0_22__I213_QOUT;
reg inst_cellmath__44_0_23__I214_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_23__I214_QOUT <= inst_cellmath__40[23];
assign inst_cellmath__44[23] = inst_cellmath__44_0_23__I214_QOUT;
reg inst_cellmath__44_0_24__I215_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_24__I215_QOUT <= inst_cellmath__40[24];
assign inst_cellmath__44[24] = inst_cellmath__44_0_24__I215_QOUT;
reg inst_cellmath__44_0_25__I216_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_25__I216_QOUT <= inst_cellmath__40[25];
assign inst_cellmath__44[25] = inst_cellmath__44_0_25__I216_QOUT;
reg inst_cellmath__44_0_26__I217_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_26__I217_QOUT <= inst_cellmath__40[26];
assign inst_cellmath__44[26] = inst_cellmath__44_0_26__I217_QOUT;
reg inst_cellmath__44_0_27__I218_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_27__I218_QOUT <= inst_cellmath__40[27];
assign inst_cellmath__44[27] = inst_cellmath__44_0_27__I218_QOUT;
reg inst_cellmath__44_0_28__I219_QOUT;
always @ (posedge clk)
	inst_cellmath__44_0_28__I219_QOUT <= inst_cellmath__40[28];
assign inst_cellmath__44[28] = inst_cellmath__44_0_28__I219_QOUT;
reg inst_cellmath__45_0_0__I220_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_0__I220_QOUT <= inst_cellmath__41[0];
assign inst_cellmath__45[0] = inst_cellmath__45_0_0__I220_QOUT;
reg inst_cellmath__45_0_1__I221_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_1__I221_QOUT <= inst_cellmath__41[1];
assign inst_cellmath__45[1] = inst_cellmath__45_0_1__I221_QOUT;
reg inst_cellmath__45_0_2__I222_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_2__I222_QOUT <= inst_cellmath__41[2];
assign inst_cellmath__45[2] = inst_cellmath__45_0_2__I222_QOUT;
reg inst_cellmath__45_0_3__I223_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_3__I223_QOUT <= inst_cellmath__41[3];
assign inst_cellmath__45[3] = inst_cellmath__45_0_3__I223_QOUT;
reg inst_cellmath__45_0_4__I224_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_4__I224_QOUT <= inst_cellmath__41[4];
assign inst_cellmath__45[4] = inst_cellmath__45_0_4__I224_QOUT;
reg inst_cellmath__45_0_5__I225_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_5__I225_QOUT <= inst_cellmath__41[5];
assign inst_cellmath__45[5] = inst_cellmath__45_0_5__I225_QOUT;
reg inst_cellmath__45_0_6__I226_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_6__I226_QOUT <= inst_cellmath__41[6];
assign inst_cellmath__45[6] = inst_cellmath__45_0_6__I226_QOUT;
reg inst_cellmath__45_0_7__I227_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_7__I227_QOUT <= inst_cellmath__41[7];
assign inst_cellmath__45[7] = inst_cellmath__45_0_7__I227_QOUT;
reg inst_cellmath__45_0_8__I228_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_8__I228_QOUT <= inst_cellmath__41[8];
assign inst_cellmath__45[8] = inst_cellmath__45_0_8__I228_QOUT;
reg inst_cellmath__45_0_9__I229_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_9__I229_QOUT <= inst_cellmath__41[9];
assign inst_cellmath__45[9] = inst_cellmath__45_0_9__I229_QOUT;
reg inst_cellmath__45_0_10__I230_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_10__I230_QOUT <= inst_cellmath__41[10];
assign inst_cellmath__45[10] = inst_cellmath__45_0_10__I230_QOUT;
reg inst_cellmath__45_0_11__I231_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_11__I231_QOUT <= inst_cellmath__41[11];
assign inst_cellmath__45[11] = inst_cellmath__45_0_11__I231_QOUT;
reg inst_cellmath__45_0_12__I232_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_12__I232_QOUT <= inst_cellmath__41[12];
assign inst_cellmath__45[12] = inst_cellmath__45_0_12__I232_QOUT;
reg inst_cellmath__45_0_13__I233_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_13__I233_QOUT <= inst_cellmath__41[13];
assign inst_cellmath__45[13] = inst_cellmath__45_0_13__I233_QOUT;
reg inst_cellmath__45_0_14__I234_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_14__I234_QOUT <= inst_cellmath__41[14];
assign inst_cellmath__45[14] = inst_cellmath__45_0_14__I234_QOUT;
reg inst_cellmath__45_0_15__I235_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_15__I235_QOUT <= inst_cellmath__41[15];
assign inst_cellmath__45[15] = inst_cellmath__45_0_15__I235_QOUT;
reg inst_cellmath__45_0_16__I236_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_16__I236_QOUT <= inst_cellmath__41[16];
assign inst_cellmath__45[16] = inst_cellmath__45_0_16__I236_QOUT;
reg inst_cellmath__45_0_17__I237_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_17__I237_QOUT <= inst_cellmath__41[17];
assign inst_cellmath__45[17] = inst_cellmath__45_0_17__I237_QOUT;
reg inst_cellmath__45_0_18__I238_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_18__I238_QOUT <= inst_cellmath__41[18];
assign inst_cellmath__45[18] = inst_cellmath__45_0_18__I238_QOUT;
reg inst_cellmath__45_0_19__I239_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_19__I239_QOUT <= inst_cellmath__41[19];
assign inst_cellmath__45[19] = inst_cellmath__45_0_19__I239_QOUT;
reg inst_cellmath__45_0_20__I240_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_20__I240_QOUT <= inst_cellmath__41[20];
assign inst_cellmath__45[20] = inst_cellmath__45_0_20__I240_QOUT;
reg inst_cellmath__45_0_21__I241_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_21__I241_QOUT <= inst_cellmath__41[21];
assign inst_cellmath__45[21] = inst_cellmath__45_0_21__I241_QOUT;
reg inst_cellmath__45_0_22__I242_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_22__I242_QOUT <= inst_cellmath__41[22];
assign inst_cellmath__45[22] = inst_cellmath__45_0_22__I242_QOUT;
reg inst_cellmath__45_0_23__I243_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_23__I243_QOUT <= inst_cellmath__41[23];
assign inst_cellmath__45[23] = inst_cellmath__45_0_23__I243_QOUT;
reg inst_cellmath__45_0_24__I244_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_24__I244_QOUT <= inst_cellmath__41[24];
assign inst_cellmath__45[24] = inst_cellmath__45_0_24__I244_QOUT;
reg inst_cellmath__45_0_25__I245_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_25__I245_QOUT <= inst_cellmath__41[25];
assign inst_cellmath__45[25] = inst_cellmath__45_0_25__I245_QOUT;
reg inst_cellmath__45_0_26__I246_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_26__I246_QOUT <= inst_cellmath__41[26];
assign inst_cellmath__45[26] = inst_cellmath__45_0_26__I246_QOUT;
reg inst_cellmath__45_0_27__I247_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_27__I247_QOUT <= inst_cellmath__41[27];
assign inst_cellmath__45[27] = inst_cellmath__45_0_27__I247_QOUT;
reg inst_cellmath__45_0_28__I248_QOUT;
always @ (posedge clk)
	inst_cellmath__45_0_28__I248_QOUT <= inst_cellmath__41[28];
assign inst_cellmath__45[28] = inst_cellmath__45_0_28__I248_QOUT;
assign inst_cellmath__124[0] = (inst_cellmath__120[25] & inst_cellmath__45[0]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[0]);
assign inst_cellmath__124[1] = (inst_cellmath__120[25] & inst_cellmath__45[1]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[1]);
assign inst_cellmath__124[2] = (inst_cellmath__120[25] & inst_cellmath__45[2]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[2]);
assign inst_cellmath__124[3] = (inst_cellmath__120[25] & inst_cellmath__45[3]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[3]);
assign inst_cellmath__124[4] = (inst_cellmath__120[25] & inst_cellmath__45[4]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[4]);
assign inst_cellmath__124[5] = (inst_cellmath__120[25] & inst_cellmath__45[5]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[5]);
assign inst_cellmath__124[6] = (inst_cellmath__120[25] & inst_cellmath__45[6]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[6]);
assign inst_cellmath__124[7] = (inst_cellmath__120[25] & inst_cellmath__45[7]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[7]);
assign inst_cellmath__124[8] = (inst_cellmath__120[25] & inst_cellmath__45[8]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[8]);
assign inst_cellmath__124[9] = (inst_cellmath__120[25] & inst_cellmath__45[9]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[9]);
assign inst_cellmath__124[10] = (inst_cellmath__120[25] & inst_cellmath__45[10]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[10]);
assign inst_cellmath__124[11] = (inst_cellmath__120[25] & inst_cellmath__45[11]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[11]);
assign inst_cellmath__124[12] = (inst_cellmath__120[25] & inst_cellmath__45[12]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[12]);
assign inst_cellmath__124[13] = (inst_cellmath__120[25] & inst_cellmath__45[13]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[13]);
assign inst_cellmath__124[14] = (inst_cellmath__120[25] & inst_cellmath__45[14]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[14]);
assign inst_cellmath__124[15] = (inst_cellmath__120[25] & inst_cellmath__45[15]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[15]);
assign inst_cellmath__124[16] = (inst_cellmath__120[25] & inst_cellmath__45[16]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[16]);
assign inst_cellmath__124[17] = (inst_cellmath__120[25] & inst_cellmath__45[17]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[17]);
assign inst_cellmath__124[18] = (inst_cellmath__120[25] & inst_cellmath__45[18]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[18]);
assign inst_cellmath__124[19] = (inst_cellmath__120[25] & inst_cellmath__45[19]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[19]);
assign inst_cellmath__124[20] = (inst_cellmath__120[25] & inst_cellmath__45[20]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[20]);
assign inst_cellmath__124[21] = (inst_cellmath__120[25] & inst_cellmath__45[21]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[21]);
assign inst_cellmath__124[22] = (inst_cellmath__120[25] & inst_cellmath__45[22]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[22]);
assign inst_cellmath__124[23] = (inst_cellmath__120[25] & inst_cellmath__45[23]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[23]);
assign inst_cellmath__124[24] = (inst_cellmath__120[25] & inst_cellmath__45[24]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[24]);
assign inst_cellmath__124[25] = (inst_cellmath__120[25] & inst_cellmath__45[25]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[25]);
assign inst_cellmath__124[26] = (inst_cellmath__120[25] & inst_cellmath__45[26]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[26]);
assign inst_cellmath__124[27] = (inst_cellmath__120[25] & inst_cellmath__45[27]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[27]);
assign inst_cellmath__122 = !((inst_cellmath__120[25] & inst_cellmath__45[28]) | ((!inst_cellmath__120[25]) & inst_cellmath__44[28]));
assign N13935 = !inst_cellmath__122;
assign N13952 = !N13935;
assign inst_cellmath__125[0] = (N13952 & inst_cellmath__124[4]) | ((!N13952) & inst_cellmath__124[5]);
assign inst_cellmath__125[1] = (N13952 & inst_cellmath__124[5]) | ((!N13952) & inst_cellmath__124[6]);
assign inst_cellmath__125[2] = (N13952 & inst_cellmath__124[6]) | ((!N13952) & inst_cellmath__124[7]);
assign inst_cellmath__125[3] = (N13952 & inst_cellmath__124[7]) | ((!N13952) & inst_cellmath__124[8]);
assign inst_cellmath__125[4] = (N13952 & inst_cellmath__124[8]) | ((!N13952) & inst_cellmath__124[9]);
assign inst_cellmath__125[5] = (N13952 & inst_cellmath__124[9]) | ((!N13952) & inst_cellmath__124[10]);
assign inst_cellmath__125[6] = (N13952 & inst_cellmath__124[10]) | ((!N13952) & inst_cellmath__124[11]);
assign inst_cellmath__125[7] = (N13952 & inst_cellmath__124[11]) | ((!N13952) & inst_cellmath__124[12]);
assign inst_cellmath__125[8] = (N13952 & inst_cellmath__124[12]) | ((!N13952) & inst_cellmath__124[13]);
assign inst_cellmath__125[9] = (N13952 & inst_cellmath__124[13]) | ((!N13952) & inst_cellmath__124[14]);
assign inst_cellmath__125[10] = (N13952 & inst_cellmath__124[14]) | ((!N13952) & inst_cellmath__124[15]);
assign inst_cellmath__125[11] = (N13952 & inst_cellmath__124[15]) | ((!N13952) & inst_cellmath__124[16]);
assign inst_cellmath__125[12] = (N13952 & inst_cellmath__124[16]) | ((!N13952) & inst_cellmath__124[17]);
assign inst_cellmath__125[13] = (N13952 & inst_cellmath__124[17]) | ((!N13952) & inst_cellmath__124[18]);
assign inst_cellmath__125[14] = (N13952 & inst_cellmath__124[18]) | ((!N13952) & inst_cellmath__124[19]);
assign inst_cellmath__125[15] = (N13952 & inst_cellmath__124[19]) | ((!N13952) & inst_cellmath__124[20]);
assign inst_cellmath__125[16] = (N13952 & inst_cellmath__124[20]) | ((!N13952) & inst_cellmath__124[21]);
assign inst_cellmath__125[17] = (N13952 & inst_cellmath__124[21]) | ((!N13952) & inst_cellmath__124[22]);
assign inst_cellmath__125[18] = (N13952 & inst_cellmath__124[22]) | ((!N13952) & inst_cellmath__124[23]);
assign inst_cellmath__125[19] = (N13952 & inst_cellmath__124[23]) | ((!N13952) & inst_cellmath__124[24]);
assign inst_cellmath__125[20] = (N13952 & inst_cellmath__124[24]) | ((!N13952) & inst_cellmath__124[25]);
assign inst_cellmath__125[21] = (N13952 & inst_cellmath__124[25]) | ((!N13952) & inst_cellmath__124[26]);
assign inst_cellmath__125[22] = !((N13952 & inst_cellmath__124[26]) | ((!N13952) & inst_cellmath__124[27]));
assign inst_cellmath__126 = (inst_cellmath__122 & inst_cellmath__124[3]) | ((!inst_cellmath__122) & inst_cellmath__124[4]);
assign {N14058, inst_cellmath__129[0]} = {1'B0, inst_cellmath__126} + {1'B0, inst_cellmath__125[0]};
assign {N14047, inst_cellmath__129[1]} = {1'B0, inst_cellmath__125[1]} + {1'B0, N14058};
assign {N14038, inst_cellmath__129[2]} = {1'B0, inst_cellmath__125[2]} + {1'B0, N14047};
assign {N14030, inst_cellmath__129[3]} = {1'B0, inst_cellmath__125[3]} + {1'B0, N14038};
assign {N14020, inst_cellmath__129[4]} = {1'B0, inst_cellmath__125[4]} + {1'B0, N14030};
assign {N14012, inst_cellmath__129[5]} = {1'B0, inst_cellmath__125[5]} + {1'B0, N14020};
assign {N14072, inst_cellmath__129[6]} = {1'B0, inst_cellmath__125[6]} + {1'B0, N14012};
assign {N14063, inst_cellmath__129[7]} = {1'B0, inst_cellmath__125[7]} + {1'B0, N14072};
assign {N14055, inst_cellmath__129[8]} = {1'B0, inst_cellmath__125[8]} + {1'B0, N14063};
assign {N14045, inst_cellmath__129[9]} = {1'B0, inst_cellmath__125[9]} + {1'B0, N14055};
assign {N14035, inst_cellmath__129[10]} = {1'B0, inst_cellmath__125[10]} + {1'B0, N14045};
assign {N14027, inst_cellmath__129[11]} = {1'B0, inst_cellmath__125[11]} + {1'B0, N14035};
assign {N14018, inst_cellmath__129[12]} = {1'B0, inst_cellmath__125[12]} + {1'B0, N14027};
assign {N14010, inst_cellmath__129[13]} = {1'B0, inst_cellmath__125[13]} + {1'B0, N14018};
assign {N14070, inst_cellmath__129[14]} = {1'B0, inst_cellmath__125[14]} + {1'B0, N14010};
assign {N14061, inst_cellmath__129[15]} = {1'B0, inst_cellmath__125[15]} + {1'B0, N14070};
assign {N14053, inst_cellmath__129[16]} = {1'B0, inst_cellmath__125[16]} + {1'B0, N14061};
assign {N14043, inst_cellmath__129[17]} = {1'B0, inst_cellmath__125[17]} + {1'B0, N14053};
assign {N14033, inst_cellmath__129[18]} = {1'B0, inst_cellmath__125[18]} + {1'B0, N14043};
assign {N14025, inst_cellmath__129[19]} = {1'B0, inst_cellmath__125[19]} + {1'B0, N14033};
assign {N14016, inst_cellmath__129[20]} = {1'B0, inst_cellmath__125[20]} + {1'B0, N14025};
assign {N14077, inst_cellmath__129[21]} = {1'B0, inst_cellmath__125[21]} + {1'B0, N14016};
assign inst_cellmath__129[22] = (!inst_cellmath__125[22]) ^ N14077;
assign N1682 = ((inst_cellmath__124[2] | inst_cellmath__124[1]) | inst_cellmath__124[3]) | inst_cellmath__124[0];
assign N1681 = (inst_cellmath__124[0] | inst_cellmath__124[1]) | inst_cellmath__124[2];
assign inst_cellmath__127 = (inst_cellmath__122 & N1681) | ((!inst_cellmath__122) & N1682);
assign N14181 = !((inst_cellmath__120[1] | inst_cellmath__120[2]) | inst_cellmath__120[6]);
assign N14169 = !((inst_cellmath__120[5] | inst_cellmath__120[11]) | inst_cellmath__120[15]);
assign N14179 = !(((!N14181) | inst_cellmath__120[14]) | inst_cellmath__120[12]);
assign N14153 = !((inst_cellmath__120[10] | inst_cellmath__120[8]) | inst_cellmath__120[9]);
assign N14173 = !((inst_cellmath__120[13] | inst_cellmath__120[16]) | inst_cellmath__120[19]);
assign N14185 = !(inst_cellmath__120[20] | inst_cellmath__120[18]);
assign N14149 = !(((inst_cellmath__120[4] | inst_cellmath__120[3]) | inst_cellmath__120[7]) | inst_cellmath__120[17]);
assign N14158 = !(inst_cellmath__120[22] | inst_cellmath__120[24]);
assign N14177 = !(N14179 & N14169);
assign N14146 = !(((N14153 & N14185) & N14149) & N14158);
assign N14165 = !((((!N14173) | inst_cellmath__120[21]) | N14146) | inst_cellmath__120[23]);
assign N14182 = !(inst_cellmath__120[25] | N14177);
assign N14160 = !((N14165 & N14182) & (!inst_cellmath__127));
assign N1922 = !(((!inst_cellmath__125[0]) & (!N14160)) | (!inst_cellmath__129[0]));
assign N1322 = !accept;
reg inst_cellmath__13_0_0__I260_QOUT;
always @ (posedge clk)
	if (N1322==1'b0)
		inst_cellmath__13_0_0__I260_QOUT <= 1'b0;
	else 
		inst_cellmath__13_0_0__I260_QOUT <= inst_cellmath__12[0];
assign inst_cellmath__13[0] = inst_cellmath__13_0_0__I260_QOUT;
reg inst_cellmath__13_0_1__I261_QOUT;
always @ (posedge clk)
	if (N1322==1'b0)
		inst_cellmath__13_0_1__I261_QOUT <= 1'b0;
	else 
		inst_cellmath__13_0_1__I261_QOUT <= inst_cellmath__12[1];
assign inst_cellmath__13[1] = inst_cellmath__13_0_1__I261_QOUT;
reg inst_cellmath__13_0_2__I262_QOUT;
always @ (posedge clk)
	if (N1322==1'b0)
		inst_cellmath__13_0_2__I262_QOUT <= 1'b0;
	else 
		inst_cellmath__13_0_2__I262_QOUT <= inst_cellmath__12[2];
assign inst_cellmath__13[2] = inst_cellmath__13_0_2__I262_QOUT;
reg inst_cellmath__13_0_3__I263_QOUT;
always @ (posedge clk)
	if (N1322==1'b0)
		inst_cellmath__13_0_3__I263_QOUT <= 1'b0;
	else 
		inst_cellmath__13_0_3__I263_QOUT <= inst_cellmath__12[3];
assign inst_cellmath__13[3] = inst_cellmath__13_0_3__I263_QOUT;
assign {N14214, N1324} = {1'B0, inst_cellmath__13[1]} + {1'B0, inst_cellmath__13[0]};
assign {N14213, N1325} = {1'B0, inst_cellmath__13[2]} + {1'B0, N14214};
assign N1326 = inst_cellmath__13[3] ^ N14213;
assign N1327 = ((inst_cellmath__13[3] & inst_cellmath__13[0]) & inst_cellmath__13[1]) & inst_cellmath__13[2];
assign inst_cellmath__12[0] = !(inst_cellmath__13[0] & (!N1327));
assign inst_cellmath__12[1] = N1327 | N1324;
assign inst_cellmath__12[2] = N1327 | N1325;
assign inst_cellmath__12[3] = N1327 | N1326;
assign inst_cellmath__46[0] = !(N12658 & (!inst_cellmath__44[0]));
assign inst_cellmath__46[1] = N12658 & inst_cellmath__44[1];
assign inst_cellmath__46[2] = N12658 & inst_cellmath__44[2];
assign inst_cellmath__46[3] = N12658 & inst_cellmath__44[3];
assign inst_cellmath__46[4] = N12658 & inst_cellmath__44[4];
assign inst_cellmath__46[5] = N12658 & inst_cellmath__44[5];
assign inst_cellmath__46[6] = N12658 & inst_cellmath__44[6];
assign inst_cellmath__46[7] = N12658 & inst_cellmath__44[7];
assign inst_cellmath__46[8] = N12658 & inst_cellmath__44[8];
assign inst_cellmath__46[9] = N12658 & inst_cellmath__44[9];
assign inst_cellmath__46[10] = N12658 & inst_cellmath__44[10];
assign inst_cellmath__46[11] = N12658 & inst_cellmath__44[11];
assign inst_cellmath__46[12] = N12658 & inst_cellmath__44[12];
assign inst_cellmath__46[13] = N12658 & inst_cellmath__44[13];
assign inst_cellmath__46[14] = N12658 & inst_cellmath__44[14];
assign inst_cellmath__46[15] = N12658 & inst_cellmath__44[15];
assign inst_cellmath__46[16] = N12658 & inst_cellmath__44[16];
assign inst_cellmath__46[17] = N12658 & inst_cellmath__44[17];
assign inst_cellmath__46[18] = N12658 & inst_cellmath__44[18];
assign inst_cellmath__46[19] = N12658 & inst_cellmath__44[19];
assign inst_cellmath__46[20] = N12658 & inst_cellmath__44[20];
assign inst_cellmath__46[21] = N12658 & inst_cellmath__44[21];
assign inst_cellmath__46[22] = N12658 & inst_cellmath__44[22];
assign inst_cellmath__46[23] = N12658 & inst_cellmath__44[23];
assign inst_cellmath__46[24] = N12658 & inst_cellmath__44[24];
assign inst_cellmath__47[0] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[0]));
assign inst_cellmath__47[1] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[1]));
assign inst_cellmath__47[2] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[2]));
assign inst_cellmath__47[3] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[3]));
assign inst_cellmath__47[4] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[4]));
assign inst_cellmath__47[5] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[5]));
assign inst_cellmath__47[6] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[6]));
assign inst_cellmath__47[7] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[7]));
assign inst_cellmath__47[8] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[8]));
assign inst_cellmath__47[9] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[9]));
assign inst_cellmath__47[10] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[10]));
assign inst_cellmath__47[11] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[11]));
assign inst_cellmath__47[12] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[12]));
assign inst_cellmath__47[13] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[13]));
assign inst_cellmath__47[14] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[14]));
assign inst_cellmath__47[15] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[15]));
assign inst_cellmath__47[16] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[16]));
assign inst_cellmath__47[17] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[17]));
assign inst_cellmath__47[18] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[18]));
assign inst_cellmath__47[19] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[19]));
assign inst_cellmath__47[20] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[20]));
assign inst_cellmath__47[21] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[21]));
assign inst_cellmath__47[22] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[22]));
assign inst_cellmath__47[23] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[23]));
assign inst_cellmath__47[24] = !(inst_cellmath__38__W0[2] | (!inst_cellmath__45[24]));
assign N1417 = !(inst_lookup0_cellmath__29[1] & inst_cellmath__42[0]);
assign inst_cellmath__42[1] = (inst_lookup0_cellmath__29[2] & N1417) | ((!inst_lookup0_cellmath__29[2]) & inst_lookup0_cellmath__29[1]);
assign inst_cellmath__42[2] = (inst_it2_cellmath__60[3] & inst_cellmath__46[0]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[0]);
assign inst_cellmath__42[3] = (inst_it2_cellmath__60[3] & inst_cellmath__46[1]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[1]);
assign inst_cellmath__42[4] = (inst_it2_cellmath__60[3] & inst_cellmath__46[2]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[2]);
assign inst_cellmath__42[5] = (inst_it2_cellmath__60[3] & inst_cellmath__46[3]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[3]);
assign inst_cellmath__42[6] = (inst_it2_cellmath__60[3] & inst_cellmath__46[4]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[4]);
assign inst_cellmath__42[7] = (inst_it2_cellmath__60[3] & inst_cellmath__46[5]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[5]);
assign inst_cellmath__42[8] = (inst_it2_cellmath__60[3] & inst_cellmath__46[6]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[6]);
assign inst_cellmath__42[9] = (inst_it2_cellmath__60[3] & inst_cellmath__46[7]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[7]);
assign inst_cellmath__42[10] = (inst_it2_cellmath__60[3] & inst_cellmath__46[8]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[8]);
assign inst_cellmath__42[11] = (inst_it2_cellmath__60[3] & inst_cellmath__46[9]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[9]);
assign inst_cellmath__42[12] = (inst_it2_cellmath__60[3] & inst_cellmath__46[10]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[10]);
assign inst_cellmath__42[13] = (inst_it2_cellmath__60[3] & inst_cellmath__46[11]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[11]);
assign inst_cellmath__42[14] = (inst_it2_cellmath__60[3] & inst_cellmath__46[12]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[12]);
assign inst_cellmath__42[15] = (inst_it2_cellmath__60[3] & inst_cellmath__46[13]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[13]);
assign inst_cellmath__42[16] = (inst_it2_cellmath__60[3] & inst_cellmath__46[14]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[14]);
assign inst_cellmath__42[17] = (inst_it2_cellmath__60[3] & inst_cellmath__46[15]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[15]);
assign inst_cellmath__42[18] = (inst_it2_cellmath__60[3] & inst_cellmath__46[16]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[16]);
assign inst_cellmath__42[19] = (inst_it2_cellmath__60[3] & inst_cellmath__46[17]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[17]);
assign inst_cellmath__42[20] = (inst_it2_cellmath__60[3] & inst_cellmath__46[18]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[18]);
assign inst_cellmath__42[21] = (inst_it2_cellmath__60[3] & inst_cellmath__46[19]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[19]);
assign inst_cellmath__42[22] = (inst_it2_cellmath__60[3] & inst_cellmath__46[20]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[20]);
assign inst_cellmath__42[23] = (inst_it2_cellmath__60[3] & inst_cellmath__46[21]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[21]);
assign inst_cellmath__42[24] = (inst_it2_cellmath__60[3] & inst_cellmath__46[22]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[22]);
assign inst_cellmath__42[25] = (inst_it2_cellmath__60[3] & inst_cellmath__46[23]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[23]);
assign inst_cellmath__42[26] = (inst_it2_cellmath__60[3] & inst_cellmath__46[24]) | ((!inst_it2_cellmath__60[3]) & inst_cellmath__47[24]);
assign inst_cellmath__43[1] = inst_cellmath__42[1] ^ inst_cellmath__43[0];
assign N14594 = !(((!inst_cellmath__42[1]) & (!inst_cellmath__42[0])) | (!inst_it2_cellmath__60[4]));
assign inst_cellmath__43[2] = (N14594 & inst_cellmath__46[0]) | ((!N14594) & inst_cellmath__47[0]);
assign inst_cellmath__43[3] = (N14594 & inst_cellmath__46[1]) | ((!N14594) & inst_cellmath__47[1]);
assign inst_cellmath__43[4] = (N14594 & inst_cellmath__46[2]) | ((!N14594) & inst_cellmath__47[2]);
assign inst_cellmath__43[5] = (N14594 & inst_cellmath__46[3]) | ((!N14594) & inst_cellmath__47[3]);
assign inst_cellmath__43[6] = (N14594 & inst_cellmath__46[4]) | ((!N14594) & inst_cellmath__47[4]);
assign inst_cellmath__43[7] = (N14594 & inst_cellmath__46[5]) | ((!N14594) & inst_cellmath__47[5]);
assign inst_cellmath__43[8] = (N14594 & inst_cellmath__46[6]) | ((!N14594) & inst_cellmath__47[6]);
assign inst_cellmath__43[9] = (N14594 & inst_cellmath__46[7]) | ((!N14594) & inst_cellmath__47[7]);
assign inst_cellmath__43[10] = (N14594 & inst_cellmath__46[8]) | ((!N14594) & inst_cellmath__47[8]);
assign inst_cellmath__43[11] = (N14594 & inst_cellmath__46[9]) | ((!N14594) & inst_cellmath__47[9]);
assign inst_cellmath__43[12] = (N14594 & inst_cellmath__46[10]) | ((!N14594) & inst_cellmath__47[10]);
assign inst_cellmath__43[13] = (N14594 & inst_cellmath__46[11]) | ((!N14594) & inst_cellmath__47[11]);
assign inst_cellmath__43[14] = (N14594 & inst_cellmath__46[12]) | ((!N14594) & inst_cellmath__47[12]);
assign inst_cellmath__43[15] = (N14594 & inst_cellmath__46[13]) | ((!N14594) & inst_cellmath__47[13]);
assign inst_cellmath__43[16] = (N14594 & inst_cellmath__46[14]) | ((!N14594) & inst_cellmath__47[14]);
assign inst_cellmath__43[17] = (N14594 & inst_cellmath__46[15]) | ((!N14594) & inst_cellmath__47[15]);
assign inst_cellmath__43[18] = (N14594 & inst_cellmath__46[16]) | ((!N14594) & inst_cellmath__47[16]);
assign inst_cellmath__43[19] = (N14594 & inst_cellmath__46[17]) | ((!N14594) & inst_cellmath__47[17]);
assign inst_cellmath__43[20] = (N14594 & inst_cellmath__46[18]) | ((!N14594) & inst_cellmath__47[18]);
assign inst_cellmath__43[21] = (N14594 & inst_cellmath__46[19]) | ((!N14594) & inst_cellmath__47[19]);
assign inst_cellmath__43[22] = (N14594 & inst_cellmath__46[20]) | ((!N14594) & inst_cellmath__47[20]);
assign inst_cellmath__43[23] = (N14594 & inst_cellmath__46[21]) | ((!N14594) & inst_cellmath__47[21]);
assign inst_cellmath__43[24] = (N14594 & inst_cellmath__46[22]) | ((!N14594) & inst_cellmath__47[22]);
assign inst_cellmath__43[25] = (N14594 & inst_cellmath__46[23]) | ((!N14594) & inst_cellmath__47[23]);
assign inst_cellmath__43[26] = (N14594 & inst_cellmath__46[24]) | ((!N14594) & inst_cellmath__47[24]);
assign inst_cellmath__14[2] = !inst_it2_lookup1_cellmath__55[2];
assign N14648 = !inst_cellmath__14[2];
assign inst_it2_cellmath__63__W1[1] = (!N2201) ^ N14648;
assign inst_it2_cellmath__56[2] = (!N2202) ^ N14648;
assign inst_it2_cellmath__56[3] = (!N2203) ^ N14648;
assign inst_it2_cellmath__56[4] = (!N2204) ^ N14648;
assign inst_it2_cellmath__56[5] = (!N2205) ^ N14648;
assign inst_it2_cellmath__56[6] = (!N2206) ^ N14648;
assign inst_it2_cellmath__56[7] = (!N2207) ^ N14648;
assign inst_it2_cellmath__56[8] = (!N2208) ^ N14648;
assign inst_it2_cellmath__56[9] = (!N2209) ^ N14648;
assign inst_it2_cellmath__56[10] = (!N2210) ^ N14648;
assign inst_it2_cellmath__56[11] = (!N2211) ^ N14648;
assign inst_it2_cellmath__56[12] = (!N2212) ^ N14648;
assign inst_it2_cellmath__56[13] = (!N2213) ^ N14648;
assign inst_it2_cellmath__56[14] = (!N2214) ^ N14648;
assign inst_it2_cellmath__56[15] = (!N2215) ^ N14648;
assign inst_it2_cellmath__56[16] = (!N2216) ^ N14648;
assign inst_it2_cellmath__56[17] = (!N2217) ^ N14648;
assign inst_it2_cellmath__56[18] = (!N2218) ^ N14648;
assign inst_it2_cellmath__56[19] = (!N2219) ^ N14648;
assign inst_it2_cellmath__56[20] = (!N2220) ^ N14648;
assign inst_it2_cellmath__56[21] = (!N2221) ^ N14648;
assign inst_it2_cellmath__56[22] = (!N2222) ^ N14648;
assign inst_it2_cellmath__56[23] = (!N2223) ^ N14648;
assign inst_it2_cellmath__56[24] = (!N2224) ^ N14648;
assign inst_it2_cellmath__57[1] = !N14648;
assign inst_it2_cellmath__57[2] = !((N2254 & N14648) | ((!N2254) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[3] = !((N2255 & N14648) | ((!N2255) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[4] = !((N2256 & N14648) | ((!N2256) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[5] = !((N2257 & N14648) | ((!N2257) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[6] = !((N2258 & N14648) | ((!N2258) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[7] = !((N2259 & N14648) | ((!N2259) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[8] = !((N2260 & N14648) | ((!N2260) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[9] = !((N2261 & N14648) | ((!N2261) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[10] = !((N2262 & N14648) | ((!N2262) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[11] = !((N2263 & N14648) | ((!N2263) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[12] = !((N2264 & N14648) | ((!N2264) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[13] = !((N2265 & N14648) | ((!N2265) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[14] = !((N2266 & N14648) | ((!N2266) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[15] = !((N2267 & N14648) | ((!N2267) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[16] = !((N2268 & N14648) | ((!N2268) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[17] = !((N2269 & N14648) | ((!N2269) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[18] = !((N2270 & N14648) | ((!N2270) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[19] = !((N2271 & N14648) | ((!N2271) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[20] = !((N2272 & N14648) | ((!N2272) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[21] = !((N2273 & N14648) | ((!N2273) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[22] = !((N2274 & N14648) | ((!N2274) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[23] = !((N2275 & N14648) | ((!N2275) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[24] = !((N2276 & N14648) | ((!N2276) & inst_it2_cellmath__57[1]));
assign inst_it2_cellmath__57[25] = !((N2277 & inst_it2_cellmath__57[1]) | ((!N2277) & N14648));
assign {inst_it2_cellmath__62__W0[3], inst_it2_cellmath__62__W1[3]} = {1'B0, inst_it2_cellmath__60[3]} + {1'B0, inst_it2_cellmath__61[3]} + {1'B0, inst_it2_cellmath__56[3]};
assign {inst_it2_cellmath__62__W0[4], inst_it2_cellmath__62__W1[4]} = {1'B0, inst_it2_cellmath__60[4]} + {1'B0, inst_it2_cellmath__61[4]} + {1'B0, inst_it2_cellmath__56[4]};
assign {inst_it2_cellmath__62__W0[5], inst_it2_cellmath__62__W1[5]} = {1'B0, inst_it2_cellmath__60[5]} + {1'B0, inst_it2_cellmath__61[5]} + {1'B0, inst_it2_cellmath__56[5]};
assign {inst_it2_cellmath__62__W0[6], inst_it2_cellmath__62__W1[6]} = {1'B0, inst_it2_cellmath__60[6]} + {1'B0, inst_it2_cellmath__61[6]} + {1'B0, inst_it2_cellmath__56[6]};
assign {inst_it2_cellmath__62__W0[7], inst_it2_cellmath__62__W1[7]} = {1'B0, inst_it2_cellmath__60[7]} + {1'B0, inst_it2_cellmath__61[7]} + {1'B0, inst_it2_cellmath__56[7]};
assign {inst_it2_cellmath__62__W0[8], inst_it2_cellmath__62__W1[8]} = {1'B0, inst_it2_cellmath__60[8]} + {1'B0, inst_it2_cellmath__61[8]} + {1'B0, inst_it2_cellmath__56[8]};
assign {inst_it2_cellmath__62__W0[9], inst_it2_cellmath__62__W1[9]} = {1'B0, inst_it2_cellmath__60[9]} + {1'B0, inst_it2_cellmath__61[9]} + {1'B0, inst_it2_cellmath__56[9]};
assign {inst_it2_cellmath__62__W0[10], inst_it2_cellmath__62__W1[10]} = {1'B0, inst_it2_cellmath__60[10]} + {1'B0, inst_it2_cellmath__61[10]} + {1'B0, inst_it2_cellmath__56[10]};
assign {inst_it2_cellmath__62__W0[11], inst_it2_cellmath__62__W1[11]} = {1'B0, inst_it2_cellmath__60[11]} + {1'B0, inst_it2_cellmath__61[11]} + {1'B0, inst_it2_cellmath__56[11]};
assign {inst_it2_cellmath__62__W0[12], inst_it2_cellmath__62__W1[12]} = {1'B0, inst_it2_cellmath__60[12]} + {1'B0, inst_it2_cellmath__61[12]} + {1'B0, inst_it2_cellmath__56[12]};
assign {inst_it2_cellmath__62__W0[13], inst_it2_cellmath__62__W1[13]} = {1'B0, inst_it2_cellmath__60[13]} + {1'B0, inst_it2_cellmath__61[13]} + {1'B0, inst_it2_cellmath__56[13]};
assign {inst_it2_cellmath__62__W0[14], inst_it2_cellmath__62__W1[14]} = {1'B0, inst_it2_cellmath__60[14]} + {1'B0, inst_it2_cellmath__61[14]} + {1'B0, inst_it2_cellmath__56[14]};
assign {inst_it2_cellmath__62__W0[15], inst_it2_cellmath__62__W1[15]} = {1'B0, inst_it2_cellmath__60[15]} + {1'B0, inst_it2_cellmath__61[15]} + {1'B0, inst_it2_cellmath__56[15]};
assign {inst_it2_cellmath__62__W0[16], inst_it2_cellmath__62__W1[16]} = {1'B0, inst_it2_cellmath__60[16]} + {1'B0, inst_it2_cellmath__61[16]} + {1'B0, inst_it2_cellmath__56[16]};
assign {inst_it2_cellmath__62__W0[17], inst_it2_cellmath__62__W1[17]} = {1'B0, inst_it2_cellmath__60[17]} + {1'B0, inst_it2_cellmath__61[17]} + {1'B0, inst_it2_cellmath__56[17]};
assign {inst_it2_cellmath__62__W0[18], inst_it2_cellmath__62__W1[18]} = {1'B0, inst_it2_cellmath__60[18]} + {1'B0, inst_it2_cellmath__61[18]} + {1'B0, inst_it2_cellmath__56[18]};
assign {inst_it2_cellmath__62__W0[19], inst_it2_cellmath__62__W1[19]} = {1'B0, inst_it2_cellmath__60[19]} + {1'B0, inst_it2_cellmath__61[19]} + {1'B0, inst_it2_cellmath__56[19]};
assign {inst_it2_cellmath__62__W0[20], inst_it2_cellmath__62__W1[20]} = {1'B0, inst_it2_cellmath__60[20]} + {1'B0, inst_it2_cellmath__61[20]} + {1'B0, inst_it2_cellmath__56[20]};
assign {inst_it2_cellmath__62__W0[21], inst_it2_cellmath__62__W1[21]} = {1'B0, inst_it2_cellmath__60[21]} + {1'B0, inst_it2_cellmath__61[21]} + {1'B0, inst_it2_cellmath__56[21]};
assign {inst_it2_cellmath__62__W0[22], inst_it2_cellmath__62__W1[22]} = {1'B0, inst_it2_cellmath__60[22]} + {1'B0, inst_it2_cellmath__61[22]} + {1'B0, inst_it2_cellmath__56[22]};
assign {inst_it2_cellmath__62__W0[23], inst_it2_cellmath__62__W1[23]} = {1'B0, inst_it2_cellmath__60[23]} + {1'B0, inst_it2_cellmath__61[23]} + {1'B0, inst_it2_cellmath__56[23]};
assign {inst_it2_cellmath__62__W0[24], inst_it2_cellmath__62__W1[24]} = {1'B0, inst_it2_cellmath__60[24]} + {1'B0, inst_it2_cellmath__61[24]} + {1'B0, inst_it2_cellmath__56[24]};
assign inst_it2_cellmath__62__W1[25] = (inst_it2_cellmath__60[25] ^ inst_it2_cellmath__61[25]) ^ inst_cellmath__14[2];
assign N28021 = !inst_cellmath__14[2];
assign inst_cellmath__14[1] = !N28021;
assign {inst_cellmath__14[3], inst_it2_cellmath__63__W1[2]} = {1'B0, inst_it2_cellmath__56[2]} + {1'B0, inst_it2_cellmath__57[2]};
assign {inst_cellmath__14[4], inst_it2_cellmath__63__W1[3]} = {1'B0, inst_it2_cellmath__62__W1[3]} + {1'B0, inst_it2_cellmath__57[3]};
assign {inst_cellmath__14[5], inst_it2_cellmath__63__W1[4]} = {1'B0, inst_it2_cellmath__62__W1[4]} + {1'B0, inst_it2_cellmath__62__W0[3]} + {1'B0, inst_it2_cellmath__57[4]};
assign {inst_cellmath__14[6], inst_it2_cellmath__63__W1[5]} = {1'B0, inst_it2_cellmath__62__W1[5]} + {1'B0, inst_it2_cellmath__62__W0[4]} + {1'B0, inst_it2_cellmath__57[5]};
assign {inst_cellmath__14[7], inst_it2_cellmath__63__W1[6]} = {1'B0, inst_it2_cellmath__62__W1[6]} + {1'B0, inst_it2_cellmath__62__W0[5]} + {1'B0, inst_it2_cellmath__57[6]};
assign {inst_cellmath__14[8], inst_it2_cellmath__63__W1[7]} = {1'B0, inst_it2_cellmath__62__W1[7]} + {1'B0, inst_it2_cellmath__62__W0[6]} + {1'B0, inst_it2_cellmath__57[7]};
assign {inst_cellmath__14[9], inst_it2_cellmath__63__W1[8]} = {1'B0, inst_it2_cellmath__62__W1[8]} + {1'B0, inst_it2_cellmath__62__W0[7]} + {1'B0, inst_it2_cellmath__57[8]};
assign {inst_cellmath__14[10], inst_it2_cellmath__63__W1[9]} = {1'B0, inst_it2_cellmath__62__W1[9]} + {1'B0, inst_it2_cellmath__62__W0[8]} + {1'B0, inst_it2_cellmath__57[9]};
assign {inst_cellmath__14[11], inst_it2_cellmath__63__W1[10]} = {1'B0, inst_it2_cellmath__62__W1[10]} + {1'B0, inst_it2_cellmath__62__W0[9]} + {1'B0, inst_it2_cellmath__57[10]};
assign {inst_cellmath__14[12], inst_it2_cellmath__63__W1[11]} = {1'B0, inst_it2_cellmath__62__W1[11]} + {1'B0, inst_it2_cellmath__62__W0[10]} + {1'B0, inst_it2_cellmath__57[11]};
assign {inst_cellmath__14[13], inst_it2_cellmath__63__W1[12]} = {1'B0, inst_it2_cellmath__62__W1[12]} + {1'B0, inst_it2_cellmath__62__W0[11]} + {1'B0, inst_it2_cellmath__57[12]};
assign {inst_cellmath__14[14], inst_it2_cellmath__63__W1[13]} = {1'B0, inst_it2_cellmath__62__W1[13]} + {1'B0, inst_it2_cellmath__62__W0[12]} + {1'B0, inst_it2_cellmath__57[13]};
assign {inst_cellmath__14[15], inst_it2_cellmath__63__W1[14]} = {1'B0, inst_it2_cellmath__62__W1[14]} + {1'B0, inst_it2_cellmath__62__W0[13]} + {1'B0, inst_it2_cellmath__57[14]};
assign {inst_cellmath__14[16], inst_it2_cellmath__63__W1[15]} = {1'B0, inst_it2_cellmath__62__W1[15]} + {1'B0, inst_it2_cellmath__62__W0[14]} + {1'B0, inst_it2_cellmath__57[15]};
assign {inst_cellmath__14[17], inst_it2_cellmath__63__W1[16]} = {1'B0, inst_it2_cellmath__62__W1[16]} + {1'B0, inst_it2_cellmath__62__W0[15]} + {1'B0, inst_it2_cellmath__57[16]};
assign {inst_cellmath__14[18], inst_it2_cellmath__63__W1[17]} = {1'B0, inst_it2_cellmath__62__W1[17]} + {1'B0, inst_it2_cellmath__62__W0[16]} + {1'B0, inst_it2_cellmath__57[17]};
assign {inst_cellmath__14[19], inst_it2_cellmath__63__W1[18]} = {1'B0, inst_it2_cellmath__62__W1[18]} + {1'B0, inst_it2_cellmath__62__W0[17]} + {1'B0, inst_it2_cellmath__57[18]};
assign {inst_cellmath__14[20], inst_it2_cellmath__63__W1[19]} = {1'B0, inst_it2_cellmath__62__W1[19]} + {1'B0, inst_it2_cellmath__62__W0[18]} + {1'B0, inst_it2_cellmath__57[19]};
assign {inst_cellmath__14[21], inst_it2_cellmath__63__W1[20]} = {1'B0, inst_it2_cellmath__62__W1[20]} + {1'B0, inst_it2_cellmath__62__W0[19]} + {1'B0, inst_it2_cellmath__57[20]};
assign {inst_cellmath__14[22], inst_it2_cellmath__63__W1[21]} = {1'B0, inst_it2_cellmath__62__W1[21]} + {1'B0, inst_it2_cellmath__62__W0[20]} + {1'B0, inst_it2_cellmath__57[21]};
assign {inst_cellmath__14[23], inst_it2_cellmath__63__W1[22]} = {1'B0, inst_it2_cellmath__62__W1[22]} + {1'B0, inst_it2_cellmath__62__W0[21]} + {1'B0, inst_it2_cellmath__57[22]};
assign {inst_cellmath__14[24], inst_it2_cellmath__63__W1[23]} = {1'B0, inst_it2_cellmath__62__W1[23]} + {1'B0, inst_it2_cellmath__62__W0[22]} + {1'B0, inst_it2_cellmath__57[23]};
assign {inst_cellmath__14[25], inst_it2_cellmath__63__W1[24]} = {1'B0, inst_it2_cellmath__62__W1[24]} + {1'B0, inst_it2_cellmath__62__W0[23]} + {1'B0, inst_it2_cellmath__57[24]};
assign {N14981, inst_it2_cellmath__63__W1[25]} = {1'B0, inst_it2_cellmath__62__W1[25]} + {1'B0, inst_it2_cellmath__62__W0[24]} + {1'B0, inst_it2_cellmath__57[25]};
assign N1555 = !(inst_it2_lookup1_cellmath__55[1] & inst_cellmath__40[0]);
assign inst_cellmath__40[1] = (inst_it2_lookup1_cellmath__55[2] & N1555) | ((!inst_it2_lookup1_cellmath__55[2]) & inst_it2_lookup1_cellmath__55[1]);
assign inst_cellmath__40[2] = (inst_cellmath__14[1] & inst_cellmath__42[0]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[0]);
assign inst_cellmath__40[3] = (inst_cellmath__14[1] & inst_cellmath__42[1]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[1]);
assign inst_cellmath__40[4] = (inst_cellmath__14[1] & inst_cellmath__42[2]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[2]);
assign inst_cellmath__40[5] = (inst_cellmath__14[1] & inst_cellmath__42[3]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[3]);
assign inst_cellmath__40[6] = (inst_cellmath__14[1] & inst_cellmath__42[4]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[4]);
assign inst_cellmath__40[7] = (inst_cellmath__14[1] & inst_cellmath__42[5]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[5]);
assign inst_cellmath__40[8] = (inst_cellmath__14[1] & inst_cellmath__42[6]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[6]);
assign inst_cellmath__40[9] = (inst_cellmath__14[1] & inst_cellmath__42[7]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[7]);
assign inst_cellmath__40[10] = (inst_cellmath__14[1] & inst_cellmath__42[8]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[8]);
assign inst_cellmath__40[11] = (inst_cellmath__14[1] & inst_cellmath__42[9]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[9]);
assign inst_cellmath__40[12] = (inst_cellmath__14[1] & inst_cellmath__42[10]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[10]);
assign inst_cellmath__40[13] = (inst_cellmath__14[1] & inst_cellmath__42[11]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[11]);
assign inst_cellmath__40[14] = (inst_cellmath__14[1] & inst_cellmath__42[12]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[12]);
assign inst_cellmath__40[15] = (inst_cellmath__14[1] & inst_cellmath__42[13]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[13]);
assign inst_cellmath__40[16] = (inst_cellmath__14[1] & inst_cellmath__42[14]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[14]);
assign inst_cellmath__40[17] = (inst_cellmath__14[1] & inst_cellmath__42[15]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[15]);
assign inst_cellmath__40[18] = (inst_cellmath__14[1] & inst_cellmath__42[16]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[16]);
assign inst_cellmath__40[19] = (inst_cellmath__14[1] & inst_cellmath__42[17]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[17]);
assign inst_cellmath__40[20] = (inst_cellmath__14[1] & inst_cellmath__42[18]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[18]);
assign inst_cellmath__40[21] = (inst_cellmath__14[1] & inst_cellmath__42[19]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[19]);
assign inst_cellmath__40[22] = (inst_cellmath__14[1] & inst_cellmath__42[20]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[20]);
assign inst_cellmath__40[23] = (inst_cellmath__14[1] & inst_cellmath__42[21]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[21]);
assign inst_cellmath__40[24] = (inst_cellmath__14[1] & inst_cellmath__42[22]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[22]);
assign inst_cellmath__40[25] = (inst_cellmath__14[1] & inst_cellmath__42[23]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[23]);
assign inst_cellmath__40[26] = (inst_cellmath__14[1] & inst_cellmath__42[24]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[24]);
assign inst_cellmath__40[27] = (inst_cellmath__14[1] & inst_cellmath__42[25]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[25]);
assign inst_cellmath__40[28] = (inst_cellmath__14[1] & inst_cellmath__42[26]) | ((!inst_cellmath__14[1]) & inst_cellmath__43[26]);
assign inst_cellmath__41[1] = inst_cellmath__40[1] ^ inst_cellmath__41[0];
assign N15334 = !(((!inst_cellmath__40[1]) & (!inst_cellmath__40[0])) | (!inst_cellmath__14[2]));
assign inst_cellmath__41[2] = (N15334 & inst_cellmath__42[0]) | ((!N15334) & inst_cellmath__43[0]);
assign inst_cellmath__41[3] = (N15334 & inst_cellmath__42[1]) | ((!N15334) & inst_cellmath__43[1]);
assign inst_cellmath__41[4] = (N15334 & inst_cellmath__42[2]) | ((!N15334) & inst_cellmath__43[2]);
assign inst_cellmath__41[5] = (N15334 & inst_cellmath__42[3]) | ((!N15334) & inst_cellmath__43[3]);
assign inst_cellmath__41[6] = (N15334 & inst_cellmath__42[4]) | ((!N15334) & inst_cellmath__43[4]);
assign inst_cellmath__41[7] = (N15334 & inst_cellmath__42[5]) | ((!N15334) & inst_cellmath__43[5]);
assign inst_cellmath__41[8] = (N15334 & inst_cellmath__42[6]) | ((!N15334) & inst_cellmath__43[6]);
assign inst_cellmath__41[9] = (N15334 & inst_cellmath__42[7]) | ((!N15334) & inst_cellmath__43[7]);
assign inst_cellmath__41[10] = (N15334 & inst_cellmath__42[8]) | ((!N15334) & inst_cellmath__43[8]);
assign inst_cellmath__41[11] = (N15334 & inst_cellmath__42[9]) | ((!N15334) & inst_cellmath__43[9]);
assign inst_cellmath__41[12] = (N15334 & inst_cellmath__42[10]) | ((!N15334) & inst_cellmath__43[10]);
assign inst_cellmath__41[13] = (N15334 & inst_cellmath__42[11]) | ((!N15334) & inst_cellmath__43[11]);
assign inst_cellmath__41[14] = (N15334 & inst_cellmath__42[12]) | ((!N15334) & inst_cellmath__43[12]);
assign inst_cellmath__41[15] = (N15334 & inst_cellmath__42[13]) | ((!N15334) & inst_cellmath__43[13]);
assign inst_cellmath__41[16] = (N15334 & inst_cellmath__42[14]) | ((!N15334) & inst_cellmath__43[14]);
assign inst_cellmath__41[17] = (N15334 & inst_cellmath__42[15]) | ((!N15334) & inst_cellmath__43[15]);
assign inst_cellmath__41[18] = (N15334 & inst_cellmath__42[16]) | ((!N15334) & inst_cellmath__43[16]);
assign inst_cellmath__41[19] = (N15334 & inst_cellmath__42[17]) | ((!N15334) & inst_cellmath__43[17]);
assign inst_cellmath__41[20] = (N15334 & inst_cellmath__42[18]) | ((!N15334) & inst_cellmath__43[18]);
assign inst_cellmath__41[21] = (N15334 & inst_cellmath__42[19]) | ((!N15334) & inst_cellmath__43[19]);
assign inst_cellmath__41[22] = (N15334 & inst_cellmath__42[20]) | ((!N15334) & inst_cellmath__43[20]);
assign inst_cellmath__41[23] = (N15334 & inst_cellmath__42[21]) | ((!N15334) & inst_cellmath__43[21]);
assign inst_cellmath__41[24] = (N15334 & inst_cellmath__42[22]) | ((!N15334) & inst_cellmath__43[22]);
assign inst_cellmath__41[25] = (N15334 & inst_cellmath__42[23]) | ((!N15334) & inst_cellmath__43[23]);
assign inst_cellmath__41[26] = (N15334 & inst_cellmath__42[24]) | ((!N15334) & inst_cellmath__43[24]);
assign inst_cellmath__41[27] = (N15334 & inst_cellmath__42[25]) | ((!N15334) & inst_cellmath__43[25]);
assign inst_cellmath__41[28] = (N15334 & inst_cellmath__42[26]) | ((!N15334) & inst_cellmath__43[26]);
assign N15444 = !inst_cellmath__9[23];
assign N15413 = !inst_cellmath__9[24];
assign N15436 = !inst_cellmath__9[25];
assign N15406 = !inst_cellmath__9[26];
assign N15431 = !inst_cellmath__9[27];
assign N15401 = !inst_cellmath__9[28];
assign N15423 = !inst_cellmath__9[29];
assign N15432 = !inst_cellmath__8[24];
assign N15424 = (!inst_cellmath__8[24]) ^ N15436;
assign N15435 = inst_cellmath__8[24] | N15436;
assign N15417 = (!inst_cellmath__8[26]) ^ N15406;
assign N15430 = inst_cellmath__8[26] | N15406;
assign N15411 = (!inst_cellmath__8[27]) ^ N15431;
assign N15421 = inst_cellmath__8[27] | N15431;
assign N15403 = (!inst_cellmath__8[28]) ^ N15401;
assign N15415 = inst_cellmath__8[28] | N15401;
assign N15398 = (!inst_cellmath__8[29]) ^ N15423;
assign N15409 = inst_cellmath__8[29] | N15423;
assign N15443 = (!inst_cellmath__8[30]) ^ inst_cellmath__9[30];
assign inst_cellmath__67[0] = (!N15444) ^ inst_cellmath__8[23];
assign N15426 = N15444 | inst_cellmath__8[23];
assign {N15418, inst_cellmath__67[1]} = {1'B0, N15413} + {1'B0, N15432} + {1'B0, N15426};
assign {N15440, inst_cellmath__67[2]} = {1'B0, inst_cellmath__8[25]} + {1'B0, N15424} + {1'B0, N15418};
assign {N15412, inst_cellmath__67[3]} = {1'B0, N15435} + {1'B0, N15417} + {1'B0, N15440};
assign {N15434, inst_cellmath__67[4]} = {1'B0, N15430} + {1'B0, N15411} + {1'B0, N15412};
assign {N15404, inst_cellmath__67[5]} = {1'B0, N15421} + {1'B0, N15403} + {1'B0, N15434};
assign {N15429, inst_cellmath__67[6]} = {1'B0, N15415} + {1'B0, N15398} + {1'B0, N15404};
assign {N15400, inst_cellmath__67[7]} = {1'B0, N15409} + {1'B0, N15443} + {1'B0, N15429};
assign N15503 = !inst_cellmath__9[30];
assign N15497 = !inst_cellmath__8[30];
assign {N15504, inst_cellmath__68[0]} = {1'B0, inst_cellmath__8[23]} + {1'B0, N15444};
assign {N15495, inst_cellmath__68[1]} = {1'B0, inst_cellmath__8[24]} + {1'B0, N15413} + {1'B0, N15504};
assign {N15518, inst_cellmath__68[2]} = {1'B0, inst_cellmath__8[25]} + {1'B0, N15436} + {1'B0, N15495};
assign {N15491, inst_cellmath__68[3]} = {1'B0, inst_cellmath__8[26]} + {1'B0, N15406} + {1'B0, N15518};
assign {N15511, inst_cellmath__68[4]} = {1'B0, inst_cellmath__8[27]} + {1'B0, N15431} + {1'B0, N15491};
assign {N15486, inst_cellmath__68[5]} = {1'B0, inst_cellmath__8[28]} + {1'B0, N15401} + {1'B0, N15511};
assign {N15506, inst_cellmath__68[6]} = {1'B0, inst_cellmath__8[29]} + {1'B0, N15423} + {1'B0, N15486};
assign {N15523, inst_cellmath__68[7]} = {1'B0, N15497} + {1'B0, N15503} + {1'B0, N15506};
assign inst_cellmath__68[8] = (!inst_cellmath__8[30]) ^ N15523;
assign inst_cellmath__68[9] = !(inst_cellmath__8[30] | N15523);
assign N15554 = inst_cellmath__68[0] & inst_cellmath__68[1];
assign N15560 = !((inst_cellmath__68[3] & inst_cellmath__68[4]) & inst_cellmath__68[7]);
assign N15552 = !(((inst_cellmath__68[2] & N15554) & inst_cellmath__68[6]) & inst_cellmath__68[5]);
assign N1675 = !(N15560 | N15552);
assign N18408 = !(inst_cellmath__68[8] | N1675);
assign inst_cellmath__69 = !(N18408 | inst_cellmath__68[9]);
assign N15585 = !(inst_cellmath__68[0] | inst_cellmath__68[1]);
assign N15589 = !(inst_cellmath__68[2] | inst_cellmath__68[3]);
assign N15582 = !(inst_cellmath__68[6] | inst_cellmath__68[7]);
assign N15583 = !inst_cellmath__68[8];
assign N15579 = !((((!N15583) | (!N15585)) | inst_cellmath__68[4]) | inst_cellmath__68[5]);
assign N1677 = !((N15589 & N15582) & N15579);
assign inst_cellmath__70 = !(N1677 & (!inst_cellmath__68[9]));
assign N15608 = !((inst_cellmath__68[1] & inst_cellmath__68[0]) & (!inst_cellmath__68[9]));
assign N15618 = ((inst_cellmath__68[2] & inst_cellmath__68[3]) & inst_cellmath__68[4]) & inst_cellmath__68[6];
assign N15605 = !((N15618 & inst_cellmath__68[7]) & (!inst_cellmath__68[8]));
assign inst_cellmath__71 = !(((!inst_cellmath__68[5]) | N15608) | N15605);
assign N15631 = !(inst_cellmath__68[4] | inst_cellmath__68[6]);
assign N15640 = !inst_cellmath__68[7];
assign N15636 = !(((N15640 & N15583) & N15589) & N15631);
assign inst_cellmath__72 = !((((!inst_cellmath__68[0]) | inst_cellmath__68[1]) | inst_cellmath__68[5]) | N15636);
assign inst_cellmath__73 = !(inst_cellmath__71 | (!inst_cellmath__69));
assign inst_cellmath__74 = inst_cellmath__72 | inst_cellmath__70;
assign N15660 = !(inst_cellmath__8[30] & inst_cellmath__8[24]);
assign N15663 = !(inst_cellmath__8[29] & inst_cellmath__8[25]);
assign N15666 = !(inst_cellmath__8[27] & inst_cellmath__8[28]);
assign N15656 = !(inst_cellmath__8[26] & inst_cellmath__8[23]);
assign inst_cellmath__75 = !(((N15663 | N15660) | N15666) | N15656);
assign N15679 = !(inst_cellmath__9[25] & inst_cellmath__9[27]);
assign N15681 = ((inst_cellmath__9[26] & inst_cellmath__9[24]) & inst_cellmath__9[29]) & inst_cellmath__9[30];
assign N18417 = !((inst_cellmath__9[28] & inst_cellmath__9[23]) & N15681);
assign inst_cellmath__76 = !(N15679 | N18417);
assign N15722 = !(inst_cellmath__8[1] | inst_cellmath__8[2]);
assign N15732 = !(inst_cellmath__8[18] | inst_cellmath__8[16]);
assign N15699 = !(inst_cellmath__8[14] | inst_cellmath__8[12]);
assign N15726 = !(inst_cellmath__8[19] | inst_cellmath__8[17]);
assign N15736 = !(inst_cellmath__8[15] | inst_cellmath__8[13]);
assign N15702 = !(inst_cellmath__8[11] | inst_cellmath__8[9]);
assign N15711 = !(inst_cellmath__8[7] | inst_cellmath__8[5]);
assign N15720 = !(inst_cellmath__8[3] | inst_cellmath__8[0]);
assign N15730 = !(inst_cellmath__8[22] | inst_cellmath__8[21]);
assign N15724 = ((inst_cellmath__8[4] | inst_cellmath__8[8]) | inst_cellmath__8[6]) | inst_cellmath__8[10];
assign N15728 = ((N15736 & N15711) & N15702) & N15726;
assign N15710 = !((N15722 & N15720) & N15730);
assign N15733 = !((N15732 & N15699) & N15728);
assign inst_cellmath__77 = ((inst_cellmath__8[20] | N15710) | N15724) | N15733;
assign N15782 = !(inst_cellmath__9[1] | inst_cellmath__9[2]);
assign N15792 = !(inst_cellmath__9[18] | inst_cellmath__9[16]);
assign N15758 = !(inst_cellmath__9[14] | inst_cellmath__9[12]);
assign N15786 = !(inst_cellmath__9[19] | inst_cellmath__9[17]);
assign N15795 = !(inst_cellmath__9[15] | inst_cellmath__9[13]);
assign N15762 = !(inst_cellmath__9[11] | inst_cellmath__9[9]);
assign N15770 = !(inst_cellmath__9[7] | inst_cellmath__9[5]);
assign N15779 = !(inst_cellmath__9[3] | inst_cellmath__9[0]);
assign N15790 = !(inst_cellmath__9[20] | inst_it2_lookup1_cellmath__53[1]);
assign N15784 = ((inst_cellmath__9[4] | inst_cellmath__9[8]) | inst_cellmath__9[6]) | inst_cellmath__9[10];
assign N15788 = ((N15795 & N15770) & N15762) & N15786;
assign N15759 = !((N15779 & N15782) & N15790);
assign N15780 = !((N15792 & N15758) & N15788);
assign inst_cellmath__78 = ((inst_it2_lookup1_cellmath__53[0] | N15759) | N15784) | N15780;
assign inst_cellmath__79 = inst_cellmath__75 & inst_cellmath__77;
assign inst_cellmath__80 = inst_cellmath__76 & inst_cellmath__78;
assign inst_cellmath__83 = !(inst_cellmath__77 | (!inst_cellmath__75));
assign inst_cellmath__84 = !(inst_cellmath__78 | (!inst_cellmath__76));
assign N15834 = !(inst_cellmath__8[30] | inst_cellmath__8[24]);
assign N15837 = !(inst_cellmath__8[29] | inst_cellmath__8[25]);
assign N15840 = !(inst_cellmath__8[27] | inst_cellmath__8[28]);
assign N15830 = !(inst_cellmath__8[26] | inst_cellmath__8[23]);
assign inst_cellmath__85 = ((N15834 & N15837) & N15840) & N15830;
assign N15852 = !(inst_cellmath__9[25] | inst_cellmath__9[27]);
assign N15855 = !(inst_cellmath__9[28] | inst_cellmath__9[23]);
assign N15858 = !(inst_cellmath__9[29] | inst_cellmath__9[24]);
assign N15848 = !(inst_cellmath__9[30] | inst_cellmath__9[26]);
assign inst_cellmath__86 = ((N15852 & N15858) & N15855) & N15848;
assign N1678 = inst_cellmath__83 & inst_cellmath__84;
assign N1679 = inst_cellmath__86 & inst_cellmath__85;
assign inst_cellmath__87 = ((N1679 | inst_cellmath__79) | inst_cellmath__80) | N1678;
assign inst_cellmath__88 = inst_cellmath__86 | inst_cellmath__83;
assign inst_cellmath__89 = inst_cellmath__85 | inst_cellmath__84;
assign inst_cellmath__91 = inst_cellmath__9[31] ^ inst_cellmath__8[31];
assign N1680 = inst_cellmath__91 | inst_cellmath__87;
assign N15943 = !(inst_cellmath__79 | (!inst_cellmath__80));
assign N15898 = !(inst_cellmath__80 | inst_cellmath__79);
assign N15964 = !((inst_cellmath__79 & inst_cellmath__8[31]) | (N15943 & inst_cellmath__9[31]));
assign N1751 = (inst_cellmath__79 & inst_cellmath__8[0]) | (N15943 & inst_cellmath__9[0]);
assign N1752 = (inst_cellmath__79 & inst_cellmath__8[1]) | (N15943 & inst_cellmath__9[1]);
assign N1753 = (inst_cellmath__79 & inst_cellmath__8[2]) | (N15943 & inst_cellmath__9[2]);
assign N1754 = (inst_cellmath__79 & inst_cellmath__8[3]) | (N15943 & inst_cellmath__9[3]);
assign N1755 = (inst_cellmath__79 & inst_cellmath__8[4]) | (N15943 & inst_cellmath__9[4]);
assign N1756 = (inst_cellmath__79 & inst_cellmath__8[5]) | (N15943 & inst_cellmath__9[5]);
assign N1757 = (inst_cellmath__79 & inst_cellmath__8[6]) | (N15943 & inst_cellmath__9[6]);
assign N1758 = (inst_cellmath__79 & inst_cellmath__8[7]) | (N15943 & inst_cellmath__9[7]);
assign N1759 = (inst_cellmath__79 & inst_cellmath__8[8]) | (N15943 & inst_cellmath__9[8]);
assign N1760 = (inst_cellmath__79 & inst_cellmath__8[9]) | (N15943 & inst_cellmath__9[9]);
assign N1761 = (inst_cellmath__79 & inst_cellmath__8[10]) | (N15943 & inst_cellmath__9[10]);
assign N1762 = (inst_cellmath__79 & inst_cellmath__8[11]) | (N15943 & inst_cellmath__9[11]);
assign N1763 = (inst_cellmath__79 & inst_cellmath__8[12]) | (N15943 & inst_cellmath__9[12]);
assign N1764 = (inst_cellmath__79 & inst_cellmath__8[13]) | (N15943 & inst_cellmath__9[13]);
assign N1765 = (inst_cellmath__79 & inst_cellmath__8[14]) | (N15943 & inst_cellmath__9[14]);
assign N1766 = (inst_cellmath__79 & inst_cellmath__8[15]) | (N15943 & inst_cellmath__9[15]);
assign N1767 = (inst_cellmath__79 & inst_cellmath__8[16]) | (N15943 & inst_cellmath__9[16]);
assign N1768 = (inst_cellmath__79 & inst_cellmath__8[17]) | (N15943 & inst_cellmath__9[17]);
assign N1769 = (inst_cellmath__79 & inst_cellmath__8[18]) | (N15943 & inst_cellmath__9[18]);
assign N1770 = (inst_cellmath__79 & inst_cellmath__8[19]) | (N15943 & inst_cellmath__9[19]);
assign N1771 = (inst_cellmath__79 & inst_cellmath__8[20]) | (N15943 & inst_cellmath__9[20]);
assign N1772 = (inst_cellmath__79 & inst_cellmath__8[21]) | (N15943 & inst_it2_lookup1_cellmath__53[0]);
assign N1750 = (!N15964) | (N15898 & N1680);
assign N28027 = !((inst_cellmath__12[0] & inst_cellmath__12[2]) & inst_cellmath__12[1]);
assign inst_cellmath__96 = !(inst_cellmath__12[3] | N28027);
reg inst_cellmath__98_0_I318_QOUT;
always @ (posedge clk)
	inst_cellmath__98_0_I318_QOUT <= N1750;
assign inst_cellmath__113[31] = inst_cellmath__98_0_I318_QOUT;
reg inst_cellmath__100_0_I319_QOUT;
always @ (posedge clk)
	inst_cellmath__100_0_I319_QOUT <= inst_cellmath__87;
assign inst_cellmath__100 = inst_cellmath__100_0_I319_QOUT;
reg inst_cellmath__101_0_I320_QOUT;
always @ (posedge clk)
	inst_cellmath__101_0_I320_QOUT <= inst_cellmath__88;
assign inst_cellmath__101 = inst_cellmath__101_0_I320_QOUT;
reg inst_cellmath__102_0_I321_QOUT;
always @ (posedge clk)
	inst_cellmath__102_0_I321_QOUT <= inst_cellmath__89;
assign inst_cellmath__102 = inst_cellmath__102_0_I321_QOUT;
reg inst_cellmath__103_0_I322_QOUT;
always @ (posedge clk)
	inst_cellmath__103_0_I322_QOUT <= inst_cellmath__69;
assign inst_cellmath__103 = inst_cellmath__103_0_I322_QOUT;
reg inst_cellmath__104_0_I323_QOUT;
always @ (posedge clk)
	inst_cellmath__104_0_I323_QOUT <= inst_cellmath__73;
assign inst_cellmath__104 = inst_cellmath__104_0_I323_QOUT;
reg inst_cellmath__105_0_I324_QOUT;
always @ (posedge clk)
	inst_cellmath__105_0_I324_QOUT <= inst_cellmath__70;
assign inst_cellmath__105 = inst_cellmath__105_0_I324_QOUT;
reg inst_cellmath__106_0_I325_QOUT;
always @ (posedge clk)
	inst_cellmath__106_0_I325_QOUT <= inst_cellmath__74;
assign inst_cellmath__106 = inst_cellmath__106_0_I325_QOUT;
reg inst_cellmath__110_0_0__I326_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_0__I326_QOUT <= inst_cellmath__67[0];
assign inst_cellmath__110[0] = inst_cellmath__110_0_0__I326_QOUT;
reg inst_cellmath__110_0_1__I327_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_1__I327_QOUT <= inst_cellmath__67[1];
assign inst_cellmath__110[1] = inst_cellmath__110_0_1__I327_QOUT;
reg inst_cellmath__110_0_2__I328_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_2__I328_QOUT <= inst_cellmath__67[2];
assign inst_cellmath__110[2] = inst_cellmath__110_0_2__I328_QOUT;
reg inst_cellmath__110_0_3__I329_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_3__I329_QOUT <= inst_cellmath__67[3];
assign inst_cellmath__110[3] = inst_cellmath__110_0_3__I329_QOUT;
reg inst_cellmath__110_0_4__I330_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_4__I330_QOUT <= inst_cellmath__67[4];
assign inst_cellmath__110[4] = inst_cellmath__110_0_4__I330_QOUT;
reg inst_cellmath__110_0_5__I331_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_5__I331_QOUT <= inst_cellmath__67[5];
assign inst_cellmath__110[5] = inst_cellmath__110_0_5__I331_QOUT;
reg inst_cellmath__110_0_6__I332_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_6__I332_QOUT <= inst_cellmath__67[6];
assign inst_cellmath__110[6] = inst_cellmath__110_0_6__I332_QOUT;
reg inst_cellmath__110_0_7__I333_QOUT;
always @ (posedge clk)
	inst_cellmath__110_0_7__I333_QOUT <= inst_cellmath__67[7];
assign inst_cellmath__110[7] = inst_cellmath__110_0_7__I333_QOUT;
reg inst_cellmath__111_0_0__I334_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_0__I334_QOUT <= inst_cellmath__68[0];
assign inst_cellmath__111[0] = inst_cellmath__111_0_0__I334_QOUT;
reg inst_cellmath__111_0_1__I335_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_1__I335_QOUT <= inst_cellmath__68[1];
assign inst_cellmath__111[1] = inst_cellmath__111_0_1__I335_QOUT;
reg inst_cellmath__111_0_2__I336_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_2__I336_QOUT <= inst_cellmath__68[2];
assign inst_cellmath__111[2] = inst_cellmath__111_0_2__I336_QOUT;
reg inst_cellmath__111_0_3__I337_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_3__I337_QOUT <= inst_cellmath__68[3];
assign inst_cellmath__111[3] = inst_cellmath__111_0_3__I337_QOUT;
reg inst_cellmath__111_0_4__I338_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_4__I338_QOUT <= inst_cellmath__68[4];
assign inst_cellmath__111[4] = inst_cellmath__111_0_4__I338_QOUT;
reg inst_cellmath__111_0_5__I339_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_5__I339_QOUT <= inst_cellmath__68[5];
assign inst_cellmath__111[5] = inst_cellmath__111_0_5__I339_QOUT;
reg inst_cellmath__111_0_6__I340_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_6__I340_QOUT <= inst_cellmath__68[6];
assign inst_cellmath__111[6] = inst_cellmath__111_0_6__I340_QOUT;
reg inst_cellmath__111_0_7__I341_QOUT;
always @ (posedge clk)
	inst_cellmath__111_0_7__I341_QOUT <= inst_cellmath__68[7];
assign inst_cellmath__111[7] = inst_cellmath__111_0_7__I341_QOUT;
reg inst_cellmath__109_0_I342_QOUT;
always @ (posedge clk)
	inst_cellmath__109_0_I342_QOUT <= inst_cellmath__96;
assign inst_cellmath__109 = inst_cellmath__109_0_I342_QOUT;
assign N4587 = !inst_cellmath__109;
assign N4594 = !N4587;
assign N16019 = !(inst_cellmath__103 | inst_cellmath__101);
assign N16014 = !inst_cellmath__100;
assign N16016 = !(((!N16014) | inst_cellmath__105) | inst_cellmath__102);
assign inst_cellmath__135 = !(N16019 & N16016);
assign N16033 = !(inst_cellmath__102 | inst_cellmath__101);
assign N16030 = !(((!N16014) | inst_cellmath__106) | inst_cellmath__104);
assign inst_cellmath__136 = !(N16033 & N16030);
assign inst_cellmath__137 = (inst_cellmath__122 & inst_cellmath__136) | ((!inst_cellmath__122) & inst_cellmath__135);
assign N16067 = !(inst_cellmath__122 | inst_cellmath__137);
assign N16083 = !(inst_cellmath__137 | (!inst_cellmath__122));
assign N16052 = !((N16083 & inst_cellmath__110[0]) | (N16067 & inst_cellmath__111[0]));
assign N16070 = !((N16083 & inst_cellmath__110[1]) | (N16067 & inst_cellmath__111[1]));
assign N16086 = !((N16083 & inst_cellmath__110[2]) | (N16067 & inst_cellmath__111[2]));
assign N16064 = !((N16083 & inst_cellmath__110[3]) | (N16067 & inst_cellmath__111[3]));
assign N16080 = !((N16083 & inst_cellmath__110[4]) | (N16067 & inst_cellmath__111[4]));
assign N16059 = !((N16083 & inst_cellmath__110[5]) | (N16067 & inst_cellmath__111[5]));
assign N16076 = !((N16083 & inst_cellmath__110[6]) | (N16067 & inst_cellmath__111[6]));
assign N16055 = !((N16083 & inst_cellmath__110[7]) | (N16067 & inst_cellmath__111[7]));
assign N16051 = !(((inst_cellmath__101 | inst_cellmath__103) | inst_cellmath__100) & inst_cellmath__137);
assign inst_cellmath__113[23] = !(N16051 & N16052);
assign inst_cellmath__113[24] = !(N16051 & N16070);
assign inst_cellmath__113[25] = !(N16051 & N16086);
assign inst_cellmath__113[26] = !(N16051 & N16064);
assign inst_cellmath__113[27] = !(N16051 & N16080);
assign inst_cellmath__113[28] = !(N16051 & N16059);
assign inst_cellmath__113[29] = !(N16051 & N16076);
assign inst_cellmath__113[30] = !(N16051 & N16055);
assign N16178 = inst_cellmath__100 & inst_cellmath__137;
assign N16122 = !inst_cellmath__137;
assign inst_cellmath__113[0] = (N16178 & inst_cellmath__112[0]) | (N16122 & N1922);
assign inst_cellmath__113[1] = (N16178 & inst_cellmath__112[1]) | (N16122 & inst_cellmath__129[1]);
assign inst_cellmath__113[2] = (N16178 & inst_cellmath__112[2]) | (N16122 & inst_cellmath__129[2]);
assign inst_cellmath__113[3] = (N16178 & inst_cellmath__112[3]) | (N16122 & inst_cellmath__129[3]);
assign inst_cellmath__113[4] = (N16178 & inst_cellmath__112[4]) | (N16122 & inst_cellmath__129[4]);
assign inst_cellmath__113[5] = (N16178 & inst_cellmath__112[5]) | (N16122 & inst_cellmath__129[5]);
assign inst_cellmath__113[6] = (N16178 & inst_cellmath__112[6]) | (N16122 & inst_cellmath__129[6]);
assign inst_cellmath__113[7] = (N16178 & inst_cellmath__112[7]) | (N16122 & inst_cellmath__129[7]);
assign inst_cellmath__113[8] = (N16178 & inst_cellmath__112[8]) | (N16122 & inst_cellmath__129[8]);
assign inst_cellmath__113[9] = (N16178 & inst_cellmath__112[9]) | (N16122 & inst_cellmath__129[9]);
assign inst_cellmath__113[10] = (N16178 & inst_cellmath__112[10]) | (N16122 & inst_cellmath__129[10]);
assign inst_cellmath__113[11] = (N16178 & inst_cellmath__112[11]) | (N16122 & inst_cellmath__129[11]);
assign inst_cellmath__113[12] = (N16178 & inst_cellmath__112[12]) | (N16122 & inst_cellmath__129[12]);
assign inst_cellmath__113[13] = (N16178 & inst_cellmath__112[13]) | (N16122 & inst_cellmath__129[13]);
assign inst_cellmath__113[14] = (N16178 & inst_cellmath__112[14]) | (N16122 & inst_cellmath__129[14]);
assign inst_cellmath__113[15] = (N16178 & inst_cellmath__112[15]) | (N16122 & inst_cellmath__129[15]);
assign inst_cellmath__113[16] = (N16178 & inst_cellmath__112[16]) | (N16122 & inst_cellmath__129[16]);
assign inst_cellmath__113[17] = (N16178 & inst_cellmath__112[17]) | (N16122 & inst_cellmath__129[17]);
assign inst_cellmath__113[18] = (N16178 & inst_cellmath__112[18]) | (N16122 & inst_cellmath__129[18]);
assign inst_cellmath__113[19] = (N16178 & inst_cellmath__112[19]) | (N16122 & inst_cellmath__129[19]);
assign inst_cellmath__113[20] = (N16178 & inst_cellmath__112[20]) | (N16122 & inst_cellmath__129[20]);
assign inst_cellmath__113[21] = (N16178 & inst_cellmath__112[21]) | (N16122 & inst_cellmath__129[21]);
assign inst_cellmath__113[22] = (inst_cellmath__129[22] & N16122) | N16178;
assign inst_cellmath__9[21] = inst_it2_lookup1_cellmath__53[0];
assign inst_cellmath__9[22] = inst_it2_lookup1_cellmath__53[1];
assign inst_cellmath__14[0] = 1'B0;
assign inst_cellmath__16[0] = 1'B0;
assign inst_cellmath__17[0] = 1'B0;
assign inst_cellmath__22[3] = inst_cellmath__22[4];
assign inst_lookup0_cellmath__27[0] = inst_it2_lookup1_cellmath__53[0];
assign inst_lookup0_cellmath__27[1] = inst_it2_lookup1_cellmath__53[1];
assign inst_lookup0_cellmath__29[0] = inst_cellmath__42[0];
assign inst_cellmath__30[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__30[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__30[2] = inst_cellmath__38__W1[2];
assign inst_cellmath__30[25] = inst_it2_cellmath__60[4];
assign inst_cellmath__31[0] = inst_cellmath__31[1];
assign inst_cellmath__34[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__34[1] = 1'B0;
assign inst_cellmath__34[2] = 1'B0;
assign inst_cellmath__35[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__35[1] = 1'B0;
assign inst_cellmath__35[2] = 1'B0;
assign inst_cellmath__38__W0[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__38__W0[1] = 1'B0;
assign inst_cellmath__38__W0[25] = 1'B0;
assign inst_cellmath__38__W1[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__38__W1[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__39__W0[0] = inst_it2_cellmath__60[3];
assign inst_cellmath__39__W0[1] = inst_it2_cellmath__60[4];
assign inst_cellmath__39__W0[2] = inst_it2_cellmath__60[5];
assign inst_cellmath__39__W0[3] = inst_it2_cellmath__60[6];
assign inst_cellmath__39__W0[4] = inst_it2_cellmath__60[7];
assign inst_cellmath__39__W0[5] = inst_it2_cellmath__60[8];
assign inst_cellmath__39__W0[6] = inst_it2_cellmath__60[9];
assign inst_cellmath__39__W0[7] = inst_it2_cellmath__60[10];
assign inst_cellmath__39__W0[8] = inst_it2_cellmath__60[11];
assign inst_cellmath__39__W0[9] = inst_it2_cellmath__60[12];
assign inst_cellmath__39__W0[10] = inst_it2_cellmath__60[13];
assign inst_cellmath__39__W0[11] = inst_it2_cellmath__60[14];
assign inst_cellmath__39__W0[12] = inst_it2_cellmath__60[15];
assign inst_cellmath__39__W0[13] = inst_it2_cellmath__60[16];
assign inst_cellmath__39__W0[14] = inst_it2_cellmath__60[17];
assign inst_cellmath__39__W0[15] = inst_it2_cellmath__60[18];
assign inst_cellmath__39__W0[16] = inst_it2_cellmath__60[19];
assign inst_cellmath__39__W0[17] = inst_it2_cellmath__60[20];
assign inst_cellmath__39__W0[18] = inst_it2_cellmath__60[21];
assign inst_cellmath__39__W0[19] = inst_it2_cellmath__60[22];
assign inst_cellmath__39__W0[20] = inst_it2_cellmath__60[23];
assign inst_cellmath__39__W0[21] = inst_it2_cellmath__60[24];
assign inst_cellmath__39__W0[22] = inst_it2_cellmath__60[25];
assign inst_cellmath__39__W0[25] = 1'B0;
assign inst_cellmath__39__W1[0] = 1'B0;
assign inst_cellmath__39__W1[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__39__W1[2] = inst_it2_cellmath__61[4];
assign inst_cellmath__39__W1[3] = inst_it2_cellmath__61[5];
assign inst_cellmath__39__W1[4] = inst_it2_cellmath__61[6];
assign inst_cellmath__39__W1[5] = inst_it2_cellmath__61[7];
assign inst_cellmath__39__W1[6] = inst_it2_cellmath__61[8];
assign inst_cellmath__39__W1[7] = inst_it2_cellmath__61[9];
assign inst_cellmath__39__W1[8] = inst_it2_cellmath__61[10];
assign inst_cellmath__39__W1[9] = inst_it2_cellmath__61[11];
assign inst_cellmath__39__W1[10] = inst_it2_cellmath__61[12];
assign inst_cellmath__39__W1[11] = inst_it2_cellmath__61[13];
assign inst_cellmath__39__W1[12] = inst_it2_cellmath__61[14];
assign inst_cellmath__39__W1[13] = inst_it2_cellmath__61[15];
assign inst_cellmath__39__W1[14] = inst_it2_cellmath__61[16];
assign inst_cellmath__39__W1[15] = inst_it2_cellmath__61[17];
assign inst_cellmath__39__W1[16] = inst_it2_cellmath__61[18];
assign inst_cellmath__39__W1[17] = inst_it2_cellmath__61[19];
assign inst_cellmath__39__W1[18] = inst_it2_cellmath__61[20];
assign inst_cellmath__39__W1[19] = inst_it2_cellmath__61[21];
assign inst_cellmath__39__W1[20] = inst_it2_cellmath__61[22];
assign inst_cellmath__39__W1[21] = inst_it2_cellmath__61[23];
assign inst_cellmath__39__W1[22] = inst_it2_cellmath__61[24];
assign inst_cellmath__39__W1[23] = inst_it2_cellmath__61[25];
assign inst_cellmath__42[27] = 1'B0;
assign inst_cellmath__42[28] = 1'B0;
assign inst_cellmath__43[27] = 1'B0;
assign inst_cellmath__43[28] = 1'B0;
assign inst_cellmath__46[25] = 1'B0;
assign inst_cellmath__46[26] = 1'B0;
assign inst_cellmath__46[27] = 1'B0;
assign inst_cellmath__46[28] = 1'B0;
assign inst_cellmath__47[25] = 1'B0;
assign inst_cellmath__47[26] = 1'B0;
assign inst_cellmath__47[27] = 1'B0;
assign inst_cellmath__47[28] = 1'B0;
assign inst_it2_lookup1_cellmath__55[0] = inst_cellmath__40[0];
assign inst_it2_cellmath__56[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__56[1] = inst_it2_cellmath__63__W1[1];
assign inst_it2_cellmath__56[25] = inst_cellmath__14[2];
assign inst_it2_cellmath__57[0] = inst_it2_cellmath__57[1];
assign inst_it2_cellmath__60[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__60[1] = 1'B0;
assign inst_it2_cellmath__60[2] = 1'B0;
assign inst_it2_cellmath__61[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__61[1] = 1'B0;
assign inst_it2_cellmath__61[2] = 1'B0;
assign inst_it2_cellmath__62__W0[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__62__W0[1] = 1'B0;
assign inst_it2_cellmath__62__W0[2] = 1'B0;
assign inst_it2_cellmath__62__W0[25] = 1'B0;
assign inst_it2_cellmath__62__W1[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__62__W1[1] = inst_it2_cellmath__63__W1[1];
assign inst_it2_cellmath__62__W1[2] = 1'B0;
assign inst_it2_cellmath__63__W1[0] = 1'B0;
assign inst_cellmath__67[8] = 1'B0;
assign inst_cellmath__67[9] = 1'B0;
assign inst_cellmath__120[0] = 1'B0;
assign inst_cellmath__124[28] = 1'B0;
endmodule

/* CADENCE  urfwQw7cqRA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



