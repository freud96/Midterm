/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:38 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_add2_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
wire  inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__23,
	inst_cellmath__24,
	inst_cellmath__27,
	inst_cellmath__28,
	inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__32;
wire [24:0] inst_cellmath__39;
wire [7:0] inst_cellmath__40;
wire [8:0] inst_cellmath__44;
wire [7:0] inst_cellmath__47;
wire [24:0] inst_cellmath__48,
	inst_cellmath__49;
wire [25:0] inst_cellmath__51;
wire  inst_cellmath__52;
wire [5:0] inst_delta;
wire [24:0] inst_cellmath__55;
wire [25:0] inst_cellmath__56;
wire  inst_cellmath__62;
wire [24:0] inst_cellmath__63;
wire [7:0] inst_cellmath__66;
wire  inst_cellmath__69,
	inst_cellmath__72,
	inst_cellmath__73,
	inst_cellmath__77;
wire N417,N418,N420,N421,N422,N423,N424 
	,N425,N426,N427,N428,N429,N430,N431,N432 
	,N433,N434,N435,N436,N437,N438,N439,N440 
	,N441,N442,N443,N444,N445,N446,N447,N448 
	,N449,N450,N451,N452,N453,N454,N455,N456 
	,N457,N458,N459,N460,N461,N462,N463,N464 
	,N465,N466,N467,N468,N469,N470,N471,N473 
	,N474,N475,N477,N478,N479,N482,N483,N485 
	,N488,N493,N495,N496,N498,N499,N500,N501 
	,N502,N504,N505,N506,N507,N509,N510,N513 
	,N514,N515,N516,N522,N539,N575,N576,N577 
	,N578,N579,N580,N581,N582,N583,N584,N585 
	,N586,N587,N588,N589,N590,N591,N592,N593 
	,N594,N595,N596,N597,N2804,N2806,N2809,N2811 
	,N2815,N2817,N2822,N2827,N2838,N2842,N2844,N2851 
	,N2888,N2914,N2988,N2992,N3010,N3014,N3131,N3133 
	,N3154,N3162,N3165,N3167,N3171,N3173,N3176,N3182 
	,N3186,N3220,N3222,N3243,N3251,N3254,N3256,N3260 
	,N3262,N3265,N3271,N3275,N3328,N3337,N3341,N3345 
	,N3350,N3353,N3376,N3378,N3379,N3380,N3381,N3383 
	,N3385,N3386,N3387,N3391,N3392,N3393,N3394,N3397 
	,N3398,N3399,N3400,N3402,N3405,N3406,N3408,N3410 
	,N3412,N3413,N3414,N3415,N3418,N3419,N3420,N3422 
	,N3423,N3425,N3426,N3428,N3429,N3432,N3433,N3434 
	,N3435,N3437,N3438,N3440,N3441,N3445,N3446,N3447 
	,N3448,N3450,N3452,N3453,N3454,N3455,N3458,N3459 
	,N3461,N3462,N3465,N3466,N3467,N3468,N3470,N3471 
	,N3472,N3474,N3475,N3476,N3479,N3480,N3481,N3482 
	,N3484,N3485,N3487,N3488,N3489,N3490,N3492,N3494 
	,N3495,N3496,N3498,N3501,N3502,N3503,N3504,N3507 
	,N3508,N3509,N3511,N3513,N3515,N3516,N3517,N3518 
	,N3520,N3521,N3523,N3525,N3526,N3531,N3533,N3534 
	,N3535,N3704,N3772,N3900,N3905,N3908,N3911,N3913 
	,N3917,N3919,N3924,N3927,N3930,N3932,N3938,N3941 
	,N3944,N3947,N3951,N3954,N3957,N3959,N3963,N3966 
	,N3971,N3974,N3977,N3980,N3983,N3985,N3990,N3993 
	,N3996,N3999,N4002,N4004,N4009,N4012,N4015,N4017 
	,N4023,N4026,N4029,N4032,N4035,N4037,N4040,N4043 
	,N4046,N4049,N4159,N4164,N4177,N4180,N4184,N4188 
	,N4193,N4197,N4200,N4206,N4210,N4216,N4220,N4224 
	,N4226,N4230,N4234,N4239,N4242,N4247,N4252,N4256 
	,N4259,N4263,N4267,N4271,N4276,N4280,N4335,N4336 
	,N4338,N4339,N4341,N4342,N4345,N4347,N4348,N4349 
	,N4351,N4352,N4354,N4355,N4359,N4360,N4362,N4364 
	,N4366,N4367,N4368,N4370,N4371,N4372,N4374,N4375 
	,N4376,N4378,N4380,N4382,N4383,N4384,N4388,N4389 
	,N4390,N4392,N4393,N4395,N4398,N4400,N4401,N4402 
	,N4404,N4405,N4407,N4408,N4411,N4412,N4414,N4415 
	,N4417,N4418,N4420,N4421,N4423,N4426,N4428,N4552 
	,N4554,N4557,N4561,N4565,N4566,N4567,N4569,N4570 
	,N4571,N4573,N4575,N4578,N4593,N4603,N4632,N4635 
	,N4636,N4639,N4640,N4641,N4644,N4645,N4646,N4650 
	,N4652,N4653,N4654,N4655,N4657,N4660,N4662,N4668 
	,N4670,N4728,N4729,N4731,N4733,N4734,N4736,N4739 
	,N4740,N4741,N4742,N4744,N4746,N4748,N4749,N4750 
	,N4752,N4753,N4755,N4758,N4759,N4760,N4762,N4763 
	,N4765,N4766,N4767,N4769,N4770,N4772,N4773,N4775 
	,N4778,N4779,N4781,N4783,N4784,N4786,N4787,N4788 
	,N4790,N4793,N4794,N4796,N4798,N4799,N4801,N4803 
	,N4804,N4806,N4807,N4809,N4811,N4812,N4814,N4816 
	,N4817,N4818,N4820,N4822,N4823,N4825,N4826,N4828 
	,N4830,N4831,N4833,N4835,N4836,N4837,N4840,N4842 
	,N4844,N4845,N4846,N4847,N4849,N4851,N4852,N4853 
	,N4855,N4856,N4858,N4859,N4861,N4863,N4864,N4866 
	,N4867,N4869,N4870,N4871,N4875,N4876,N4878,N4880 
	,N4881,N4883,N4884,N4885,N4887,N4888,N4890,N4893 
	,N4895,N4897,N4898,N6142,N6143,N6144,N6145,N6146 
	,N6147,N6148,N6149,N6150,N6152,N6154,N6161,N6165 
	,N6173,N6178,N6187,N6195,N6205,N6212,N6216,N10018 
	,N10019,N10111,N10124,N10128,N10133,N10141,N10144,N10152 
	,N10157,N10162,N10167,N10197,N10202,N10208,N10209,N10211 
	,N10216,N10217,N10220,N10221,N10223,N10290,N10297,N10324 
	,N10327,N10339,N10346,N10347,N10362,N10363,N10367,N10369 
	,N10374,N10377,N10417,N10423;
CLKINVX4 cynw_cm_float_add2_I0 (.Y(N500), .A(a_exp[0]));
INVX1 cynw_cm_float_add2_I1 (.Y(N501), .A(a_exp[1]));
INVXL cynw_cm_float_add2_I2 (.Y(N502), .A(a_exp[2]));
INVXL cynw_cm_float_add2_I4 (.Y(N504), .A(a_exp[4]));
INVXL cynw_cm_float_add2_I5 (.Y(N505), .A(a_exp[5]));
ADDHX1 inst_cellmath__43_1_I388 (.CO(N2817), .S(N509), .A(b_exp[0]), .B(N500));
ADDFHXL inst_cellmath__43_1_I389 (.CO(N2811), .S(N510), .A(N501), .B(b_exp[1]), .CI(N2817));
INVXL inst_cellmath__49_0_I5375 (.Y(N10362), .A(a_exp[3]));
ADDFHXL inst_cellmath__49_0_I5376 (.CO(N10327), .S(N10377), .A(N502), .B(b_exp[2]), .CI(N2811));
ADDFHXL inst_cellmath__49_0_I5377 (.CO(N2804), .S(N10339), .A(N10362), .B(b_exp[3]), .CI(N10327));
ADDFHXL inst_cellmath__43_1_I392 (.CO(N2827), .S(N513), .A(N504), .B(b_exp[4]), .CI(N2804));
XOR2XL inst_cellmath__43_1_I397 (.Y(inst_cellmath__44[0]), .A(N500), .B(b_exp[0]));
NOR2X1 or2_A_I2177 (.Y(N6178), .A(N500), .B(b_exp[0]));
INVXL or2_A_I2178 (.Y(N2806), .A(N6178));
ADDFXL inst_cellmath__43_1_I399 (.CO(N2851), .S(inst_cellmath__44[1]), .A(N501), .B(b_exp[1]), .CI(N2806));
ADDFXL inst_cellmath__43_1_I400 (.CO(N2822), .S(inst_cellmath__44[2]), .A(N502), .B(b_exp[2]), .CI(N2851));
ADDFX1 inst_cellmath__49_0_I5378 (.CO(N2844), .S(N10367), .A(N10362), .B(b_exp[3]), .CI(N2822));
ADDFXL inst_cellmath__43_1_I402 (.CO(N2815), .S(inst_cellmath__44[4]), .A(N504), .B(b_exp[4]), .CI(N2844));
ADDFXL inst_cellmath__43_1_I403 (.CO(N2838), .S(inst_cellmath__44[5]), .A(N505), .B(b_exp[5]), .CI(N2815));
INVXL cynw_cm_float_add2_I5368 (.Y(N506), .A(a_exp[6]));
ADDFXL inst_cellmath__43_1_I404 (.CO(N2809), .S(inst_cellmath__44[6]), .A(N506), .B(b_exp[6]), .CI(N2838));
INVXL cynw_cm_float_add2_I5369 (.Y(N507), .A(a_exp[7]));
ADDFHXL cynw_cm_float_add2_I5370 (.CO(N10290), .S(N514), .A(N505), .B(b_exp[5]), .CI(N2827));
ADDFHXL cynw_cm_float_add2_I5371 (.CO(N10297), .S(N515), .A(N506), .B(b_exp[6]), .CI(N10290));
ADDFHX1 cynw_cm_float_add2_I5372 (.CO(N2842), .S(N516), .A(N507), .B(b_exp[7]), .CI(N10297));
INVX3 cynw_cm_float_add2_I5373 (.Y(N10111), .A(N2842));
CLKINVX16 cynw_cm_float_add2_I5269 (.Y(N2914), .A(N10111));
MX2XL cynw_cm_float_add2_I409 (.Y(inst_cellmath__48[1]), .A(b_man[0]), .B(a_man[0]), .S0(N2914));
MX2XL cynw_cm_float_add2_I410 (.Y(inst_cellmath__48[2]), .A(b_man[1]), .B(a_man[1]), .S0(N2914));
MX2XL cynw_cm_float_add2_I411 (.Y(inst_cellmath__48[3]), .A(b_man[2]), .B(a_man[2]), .S0(N2914));
MX2XL cynw_cm_float_add2_I412 (.Y(inst_cellmath__48[4]), .A(b_man[3]), .B(a_man[3]), .S0(N2914));
MX2XL cynw_cm_float_add2_I413 (.Y(inst_cellmath__48[5]), .A(b_man[4]), .B(a_man[4]), .S0(N2914));
MX2XL cynw_cm_float_add2_I414 (.Y(inst_cellmath__48[6]), .A(b_man[5]), .B(a_man[5]), .S0(N2914));
MX2XL cynw_cm_float_add2_I415 (.Y(inst_cellmath__48[7]), .A(b_man[6]), .B(a_man[6]), .S0(N2914));
MX2XL cynw_cm_float_add2_I416 (.Y(inst_cellmath__48[8]), .A(b_man[7]), .B(a_man[7]), .S0(N2914));
MX2XL cynw_cm_float_add2_I417 (.Y(inst_cellmath__48[9]), .A(b_man[8]), .B(a_man[8]), .S0(N2914));
MX2XL cynw_cm_float_add2_I418 (.Y(inst_cellmath__48[10]), .A(b_man[9]), .B(a_man[9]), .S0(N2914));
MX2XL cynw_cm_float_add2_I5409 (.Y(inst_cellmath__48[11]), .A(b_man[10]), .B(a_man[10]), .S0(N2842));
INVXL buf1_A_I5472 (.Y(N10417), .A(N10111));
INVXL buf1_A_I5473 (.Y(N2888), .A(N10417));
MX2XL cynw_cm_float_add2_I2067 (.Y(inst_cellmath__48[12]), .A(b_man[11]), .B(a_man[11]), .S0(N2914));
MX2XL cynw_cm_float_add2_I421 (.Y(inst_cellmath__48[13]), .A(b_man[12]), .B(a_man[12]), .S0(N2914));
MX2XL cynw_cm_float_add2_I422 (.Y(inst_cellmath__48[14]), .A(b_man[13]), .B(a_man[13]), .S0(N2914));
MX2XL cynw_cm_float_add2_I423 (.Y(inst_cellmath__48[15]), .A(b_man[14]), .B(a_man[14]), .S0(N2914));
MX2XL cynw_cm_float_add2_I424 (.Y(inst_cellmath__48[16]), .A(b_man[15]), .B(a_man[15]), .S0(N2914));
MX2XL cynw_cm_float_add2_I425 (.Y(inst_cellmath__48[17]), .A(b_man[16]), .B(a_man[16]), .S0(N2914));
MX2XL cynw_cm_float_add2_I426 (.Y(inst_cellmath__48[18]), .A(b_man[17]), .B(a_man[17]), .S0(N2914));
MX2XL cynw_cm_float_add2_I427 (.Y(inst_cellmath__48[19]), .A(b_man[18]), .B(a_man[18]), .S0(N2914));
MX2XL cynw_cm_float_add2_I428 (.Y(inst_cellmath__48[20]), .A(b_man[19]), .B(a_man[19]), .S0(N2914));
MX2XL cynw_cm_float_add2_I429 (.Y(inst_cellmath__48[21]), .A(b_man[20]), .B(a_man[20]), .S0(N2914));
MX2XL cynw_cm_float_add2_I430 (.Y(inst_cellmath__48[22]), .A(b_man[21]), .B(a_man[21]), .S0(N2914));
MX2XL cynw_cm_float_add2_I431 (.Y(inst_cellmath__48[23]), .A(b_man[22]), .B(a_man[22]), .S0(N2914));
INVXL cynw_cm_float_add2_I5180 (.Y(N10018), .A(a_exp[0]));
INVX1 cynw_cm_float_add2_I5181 (.Y(N10019), .A(N10018));
OR4X1 inst_cellmath__28__5__I5410 (.Y(N2988), .A(a_exp[7]), .B(a_exp[1]), .C(a_exp[6]), .D(N10019));
OR4X1 inst_cellmath__28__5__I5411 (.Y(N2992), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
OR4X1 inst_cellmath__31__7__I5412 (.Y(N3010), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 inst_cellmath__31__7__I5413 (.Y(N3014), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
MX2XL cynw_cm_float_add2_I448 (.Y(N575), .A(a_man[0]), .B(b_man[0]), .S0(N2914));
MX2XL cynw_cm_float_add2_I449 (.Y(N576), .A(a_man[1]), .B(b_man[1]), .S0(N2914));
MX2XL cynw_cm_float_add2_I450 (.Y(N577), .A(a_man[2]), .B(b_man[2]), .S0(N2914));
MX2XL cynw_cm_float_add2_I451 (.Y(N578), .A(a_man[3]), .B(b_man[3]), .S0(N2914));
MX2XL cynw_cm_float_add2_I452 (.Y(N579), .A(a_man[4]), .B(b_man[4]), .S0(N2914));
MX2XL cynw_cm_float_add2_I453 (.Y(N580), .A(a_man[5]), .B(b_man[5]), .S0(N2914));
MX2XL cynw_cm_float_add2_I454 (.Y(N581), .A(a_man[6]), .B(b_man[6]), .S0(N2914));
MX2XL cynw_cm_float_add2_I455 (.Y(N582), .A(a_man[7]), .B(b_man[7]), .S0(N2914));
MX2XL cynw_cm_float_add2_I456 (.Y(N583), .A(a_man[8]), .B(b_man[8]), .S0(N2914));
MX2XL cynw_cm_float_add2_I457 (.Y(N584), .A(a_man[9]), .B(b_man[9]), .S0(N2914));
MX2XL cynw_cm_float_add2_I458 (.Y(N585), .A(a_man[10]), .B(b_man[10]), .S0(N2914));
MX2XL cynw_cm_float_add2_I459 (.Y(N586), .A(a_man[11]), .B(b_man[11]), .S0(N2914));
MX2XL cynw_cm_float_add2_I460 (.Y(N587), .A(a_man[12]), .B(b_man[12]), .S0(N2914));
MX2XL cynw_cm_float_add2_I461 (.Y(N588), .A(a_man[13]), .B(b_man[13]), .S0(N2914));
MX2XL cynw_cm_float_add2_I462 (.Y(N589), .A(a_man[14]), .B(b_man[14]), .S0(N2914));
MX2XL cynw_cm_float_add2_I463 (.Y(N590), .A(a_man[15]), .B(b_man[15]), .S0(N2914));
MX2XL cynw_cm_float_add2_I464 (.Y(N591), .A(a_man[16]), .B(b_man[16]), .S0(N2914));
MX2XL cynw_cm_float_add2_I465 (.Y(N592), .A(a_man[17]), .B(b_man[17]), .S0(N2914));
MX2XL cynw_cm_float_add2_I466 (.Y(N593), .A(a_man[18]), .B(b_man[18]), .S0(N2914));
MX2XL cynw_cm_float_add2_I467 (.Y(N594), .A(a_man[19]), .B(b_man[19]), .S0(N2914));
MX2XL cynw_cm_float_add2_I468 (.Y(N595), .A(a_man[20]), .B(b_man[20]), .S0(N2914));
MX2XL cynw_cm_float_add2_I469 (.Y(N596), .A(a_man[21]), .B(b_man[21]), .S0(N2914));
MX2XL cynw_cm_float_add2_I470 (.Y(N597), .A(a_man[22]), .B(b_man[22]), .S0(N2914));
NAND2XL inst_cellmath__30_0_I471 (.Y(N3131), .A(b_exp[0]), .B(b_exp[1]));
AND4XL inst_cellmath__30_0_I5414 (.Y(N3133), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I2179 (.Y(N6187), .A(b_exp[7]), .B(b_exp[6]), .C(N3133));
NOR2XL hyperpropagate_4_1_A_I2180 (.Y(inst_cellmath__30), .A(N3131), .B(N6187));
NOR2XL inst_cellmath__32__8__I484 (.Y(N3154), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__32__8__I485 (.Y(N3162), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__32__8__I486 (.Y(N3173), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__32__8__I487 (.Y(N3182), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__32__8__I5415 (.Y(N3167), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__32__8__I5416 (.Y(N3176), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__32__8__I5417 (.Y(N3186), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__32__8__I491 (.Y(N3171), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N3167));
NAND4XL inst_cellmath__32__8__I493 (.Y(N3165), .A(N3154), .B(N3173), .C(N3162), .D(N3182));
NOR4BX1 inst_cellmath__32__8__I5418 (.Y(inst_cellmath__32), .AN(N3171), .B(N3165), .C(N3176), .D(N3186));
AND2XL cynw_cm_float_add2_I496 (.Y(inst_cellmath__24), .A(inst_cellmath__30), .B(inst_cellmath__32));
XOR2XL cynw_cm_float_add2_I497 (.Y(inst_cellmath__55[0]), .A(a_sign), .B(b_sign));
NAND2XL inst_cellmath__27_0_I498 (.Y(N3220), .A(N10019), .B(a_exp[1]));
AND4XL inst_cellmath__27_0_I5419 (.Y(N3222), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I2181 (.Y(N6195), .A(a_exp[7]), .B(a_exp[6]), .C(N3222));
NOR2XL hyperpropagate_4_1_A_I2182 (.Y(inst_cellmath__27), .A(N3220), .B(N6195));
NOR2XL inst_cellmath__29__6__I511 (.Y(N3243), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__29__6__I512 (.Y(N3251), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__29__6__I513 (.Y(N3262), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__29__6__I514 (.Y(N3271), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__29__6__I5420 (.Y(N3256), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__29__6__I5421 (.Y(N3265), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__29__6__I5422 (.Y(N3275), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__29__6__I518 (.Y(N3260), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N3256));
NAND4XL inst_cellmath__29__6__I520 (.Y(N3254), .A(N3243), .B(N3262), .C(N3251), .D(N3271));
NOR4BX1 inst_cellmath__29__6__I5423 (.Y(inst_cellmath__29), .AN(N3260), .B(N3254), .C(N3265), .D(N3275));
AND2XL cynw_cm_float_add2_I523 (.Y(inst_cellmath__21), .A(inst_cellmath__27), .B(inst_cellmath__29));
AND3XL cynw_cm_float_add2_I524 (.Y(N495), .A(inst_cellmath__24), .B(inst_cellmath__21), .C(inst_cellmath__55[0]));
NOR2BX1 cynw_cm_float_add2_I525 (.Y(inst_cellmath__20), .AN(inst_cellmath__27), .B(inst_cellmath__29));
NOR2BX1 cynw_cm_float_add2_I526 (.Y(inst_cellmath__23), .AN(inst_cellmath__30), .B(inst_cellmath__32));
OR3XL cynw_cm_float_add2_I527 (.Y(inst_cellmath__62), .A(inst_cellmath__23), .B(inst_cellmath__20), .C(N495));
INVXL inst_cellmath__47_0_I529 (.Y(N3341), .A(inst_cellmath__44[1]));
INVXL inst_cellmath__47_0_I532 (.Y(N3328), .A(inst_cellmath__44[4]));
INVXL inst_cellmath__47_0_I533 (.Y(N3337), .A(inst_cellmath__44[5]));
INVXL inst_cellmath__47_0_I534 (.Y(N3345), .A(inst_cellmath__44[6]));
ADDFX1 inst_cellmath__49_0_I5379 (.CO(N10347), .S(inst_cellmath__44[7]), .A(N507), .B(b_exp[7]), .CI(N2809));
INVXL inst_cellmath__47_0_I535 (.Y(N3353), .A(inst_cellmath__44[7]));
INVX3 inst_cellmath__49_0_I5380 (.Y(inst_cellmath__44[8]), .A(N10347));
CLKINVX4 inst_cellmath__49_0_I5383 (.Y(N3350), .A(inst_cellmath__44[8]));
AOI22X4 inst_cellmath__47_0_I2008 (.Y(inst_cellmath__47[0]), .A0(N509), .A1(inst_cellmath__44[8]), .B0(inst_cellmath__44[0]), .B1(N3350));
AOI22X2 inst_cellmath__47_0_I538 (.Y(inst_cellmath__47[1]), .A0(N3341), .A1(N3350), .B0(N510), .B1(inst_cellmath__44[8]));
INVX8 inst_cellmath__49_0_I548 (.Y(N3455), .A(inst_cellmath__47[0]));
NOR2BX1 inst_cellmath__49_0_I549 (.Y(N3513), .AN(inst_cellmath__48[1]), .B(N3455));
MX2XL inst_cellmath__49_0_I550 (.Y(N3425), .A(inst_cellmath__48[2]), .B(inst_cellmath__48[1]), .S0(N3455));
MX2XL inst_cellmath__49_0_I552 (.Y(N3496), .A(inst_cellmath__48[4]), .B(inst_cellmath__48[3]), .S0(N3455));
MX2XL inst_cellmath__49_0_I554 (.Y(N3406), .A(inst_cellmath__48[6]), .B(inst_cellmath__48[5]), .S0(N3455));
MX2XL inst_cellmath__49_0_I556 (.Y(N3475), .A(inst_cellmath__48[8]), .B(inst_cellmath__48[7]), .S0(N3455));
MX2XL inst_cellmath__49_0_I558 (.Y(N3387), .A(inst_cellmath__48[10]), .B(inst_cellmath__48[9]), .S0(N3455));
MX2XL inst_cellmath__49_0_I560 (.Y(N3454), .A(inst_cellmath__48[12]), .B(inst_cellmath__48[11]), .S0(N3455));
MX2XL inst_cellmath__49_0_I562 (.Y(N3525), .A(inst_cellmath__48[14]), .B(inst_cellmath__48[13]), .S0(N3455));
MX2XL inst_cellmath__49_0_I564 (.Y(N3434), .A(inst_cellmath__48[16]), .B(inst_cellmath__48[15]), .S0(N3455));
MX2XL inst_cellmath__49_0_I566 (.Y(N3503), .A(inst_cellmath__48[18]), .B(inst_cellmath__48[17]), .S0(N3455));
MX2XL inst_cellmath__49_0_I567 (.Y(N3380), .A(inst_cellmath__48[19]), .B(inst_cellmath__48[18]), .S0(N3455));
MX2XL inst_cellmath__49_0_I568 (.Y(N3414), .A(inst_cellmath__48[20]), .B(inst_cellmath__48[19]), .S0(N3455));
MX2XL inst_cellmath__49_0_I569 (.Y(N3447), .A(inst_cellmath__48[21]), .B(inst_cellmath__48[20]), .S0(N3455));
MX2XL inst_cellmath__49_0_I570 (.Y(N3481), .A(inst_cellmath__48[22]), .B(inst_cellmath__48[21]), .S0(N3455));
MX2XL inst_cellmath__49_0_I571 (.Y(N3517), .A(inst_cellmath__48[23]), .B(inst_cellmath__48[22]), .S0(N3455));
NAND2BXL inst_cellmath__49_0_I572 (.Y(N3393), .AN(inst_cellmath__48[23]), .B(N3455));
INVX3 inst_cellmath__49_0_I5392 (.Y(N3490), .A(inst_cellmath__47[1]));
INVX3 inst_cellmath__49_0_I5393 (.Y(N3526), .A(N3490));
MX2X1 inst_cellmath__49_0_I5384 (.Y(N3459), .A(inst_cellmath__48[3]), .B(inst_cellmath__48[2]), .S0(N3455));
AOI22XL inst_cellmath__49_0_I575 (.Y(N3458), .A0(N3526), .A1(N3459), .B0(N3513), .B1(N3490));
AOI22XL inst_cellmath__49_0_I576 (.Y(N3495), .A0(N3526), .A1(N3496), .B0(N3425), .B1(N3490));
AOI22XL inst_cellmath__49_0_I578 (.Y(N3405), .A0(N3526), .A1(N3406), .B0(N3496), .B1(N3490));
MX2XL inst_cellmath__49_0_I5386 (.Y(N3441), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[6]), .S0(N3455));
MX2XL inst_cellmath__49_0_I5385 (.Y(N3531), .A(inst_cellmath__48[5]), .B(inst_cellmath__48[4]), .S0(N3455));
AOI22XL inst_cellmath__49_0_I579 (.Y(N3440), .A0(N3526), .A1(N3441), .B0(N3531), .B1(N3490));
AOI22XL inst_cellmath__49_0_I580 (.Y(N3474), .A0(N3526), .A1(N3475), .B0(N3406), .B1(N3490));
AOI22XL inst_cellmath__49_0_I582 (.Y(N3386), .A0(N3526), .A1(N3387), .B0(N3475), .B1(N3490));
MX2XL inst_cellmath__49_0_I5388 (.Y(N3420), .A(inst_cellmath__48[11]), .B(inst_cellmath__48[10]), .S0(N3455));
MX2X1 inst_cellmath__49_0_I5387 (.Y(N3509), .A(inst_cellmath__48[9]), .B(inst_cellmath__48[8]), .S0(N3455));
AOI22X2 inst_cellmath__49_0_I583 (.Y(N3419), .A0(N3526), .A1(N3420), .B0(N3509), .B1(N3490));
AOI22X1 inst_cellmath__49_0_I584 (.Y(N3453), .A0(N3526), .A1(N3454), .B0(N3387), .B1(N3490));
AOI22XL inst_cellmath__49_0_I586 (.Y(N3523), .A0(N3526), .A1(N3525), .B0(N3454), .B1(N3490));
MX2X1 inst_cellmath__49_0_I5390 (.Y(N3399), .A(inst_cellmath__48[15]), .B(inst_cellmath__48[14]), .S0(N3455));
MX2XL inst_cellmath__49_0_I5389 (.Y(N3489), .A(inst_cellmath__48[13]), .B(inst_cellmath__48[12]), .S0(N3455));
AOI22X2 inst_cellmath__49_0_I587 (.Y(N3398), .A0(N3526), .A1(N3399), .B0(N3489), .B1(N3490));
AOI22X1 inst_cellmath__49_0_I588 (.Y(N3433), .A0(N3526), .A1(N3434), .B0(N3525), .B1(N3490));
AOI22XL inst_cellmath__49_0_I590 (.Y(N3502), .A0(N3526), .A1(N3503), .B0(N3434), .B1(N3490));
MX2X1 inst_cellmath__49_0_I5391 (.Y(N3467), .A(inst_cellmath__48[17]), .B(inst_cellmath__48[16]), .S0(N3455));
AOI22X1 inst_cellmath__49_0_I591 (.Y(N3378), .A0(N3526), .A1(N3380), .B0(N3467), .B1(N3490));
AOI22XL inst_cellmath__49_0_I592 (.Y(N3412), .A0(N3526), .A1(N3414), .B0(N3503), .B1(N3490));
AOI22XL inst_cellmath__49_0_I593 (.Y(N3446), .A0(N3526), .A1(N3447), .B0(N3380), .B1(N3490));
AOI22XL inst_cellmath__49_0_I594 (.Y(N3480), .A0(N3526), .A1(N3481), .B0(N3414), .B1(N3490));
AOI22X1 inst_cellmath__49_0_I595 (.Y(N3516), .A0(N3526), .A1(N3517), .B0(N3447), .B1(N3490));
AOI22XL inst_cellmath__49_0_I596 (.Y(N3392), .A0(N3526), .A1(N3393), .B0(N3481), .B1(N3490));
AOI22XL inst_cellmath__49_0_I597 (.Y(N3428), .A0(N3526), .A1(N3455), .B0(N3517), .B1(N3490));
NAND2XL inst_cellmath__49_0_I598 (.Y(N3461), .A(N3393), .B(N3490));
NAND2XL inst_cellmath__49_0_I599 (.Y(N3534), .A(N3455), .B(N3490));
INVXL inst_cellmath__49_0_I5381 (.Y(N10374), .A(inst_cellmath__44[2]));
AO22X1 inst_cellmath__49_0_I5401 (.Y(N3437), .A0(N10377), .A1(inst_cellmath__44[8]), .B0(N10374), .B1(N3350));
INVX2 inst_cellmath__49_0_I5402 (.Y(N3470), .A(N3437));
AOI22X1 inst_cellmath__49_0_I602 (.Y(N3494), .A0(N3437), .A1(N3458), .B0(N3440), .B1(N3470));
AOI22XL inst_cellmath__49_0_I605 (.Y(N3438), .A0(N3437), .A1(N3405), .B0(N3386), .B1(N3470));
AOI22XL inst_cellmath__49_0_I606 (.Y(N3472), .A0(N3437), .A1(N3440), .B0(N3419), .B1(N3470));
AOI22XL inst_cellmath__49_0_I607 (.Y(N3507), .A0(N3437), .A1(N3474), .B0(N3453), .B1(N3470));
INVX1 inst_cellmath__49_0_I5394 (.Y(N10346), .A(N3526));
AOI22XL inst_cellmath__49_0_I5426 (.Y(N3508), .A0(N3526), .A1(N3509), .B0(N3441), .B1(N10346));
AOI22XL inst_cellmath__49_0_I5427 (.Y(N3487), .A0(N3489), .A1(N3526), .B0(N3420), .B1(N10346));
AOI22XL inst_cellmath__49_0_I608 (.Y(N3385), .A0(N3437), .A1(N3508), .B0(N3487), .B1(N3470));
AOI22XL inst_cellmath__49_0_I609 (.Y(N3418), .A0(N3437), .A1(N3386), .B0(N3523), .B1(N3470));
AOI22X2 inst_cellmath__49_0_I610 (.Y(N3452), .A0(N3437), .A1(N3419), .B0(N3398), .B1(N3470));
AOI22XL inst_cellmath__49_0_I613 (.Y(N3397), .A0(N3437), .A1(N3523), .B0(N3502), .B1(N3470));
AOI22XL inst_cellmath__49_0_I614 (.Y(N3432), .A0(N3437), .A1(N3398), .B0(N3378), .B1(N3470));
AOI22XL inst_cellmath__49_0_I615 (.Y(N3465), .A0(N3437), .A1(N3433), .B0(N3412), .B1(N3470));
AOI22X1 inst_cellmath__49_0_I5400 (.Y(N3466), .A0(N3526), .A1(N3467), .B0(N3399), .B1(N10346));
AOI22XL inst_cellmath__49_0_I616 (.Y(N3501), .A0(N3437), .A1(N3466), .B0(N3446), .B1(N3470));
AOI22XL inst_cellmath__49_0_I617 (.Y(N3376), .A0(N3437), .A1(N3502), .B0(N3480), .B1(N3470));
AOI22X1 inst_cellmath__49_0_I618 (.Y(N3410), .A0(N3437), .A1(N3378), .B0(N3516), .B1(N3470));
AOI22XL inst_cellmath__49_0_I620 (.Y(N3479), .A0(N3437), .A1(N3446), .B0(N3428), .B1(N3470));
AOI22XL inst_cellmath__49_0_I621 (.Y(N3515), .A0(N3437), .A1(N3480), .B0(N3461), .B1(N3470));
AOI22XL inst_cellmath__49_0_I622 (.Y(N3391), .A0(N3437), .A1(N3516), .B0(N3534), .B1(N3470));
NOR2XL inst_cellmath__49_0_I623 (.Y(N3426), .A(N3470), .B(N3392));
NOR2XL inst_cellmath__49_0_I624 (.Y(N3533), .A(N3470), .B(N3428));
NOR2XL inst_cellmath__49_0_I625 (.Y(N3476), .A(N3470), .B(N3461));
NOR2XL inst_cellmath__49_0_I626 (.Y(N3422), .A(N3470), .B(N3534));
NOR2XL inst_cellmath__49_0_I5275 (.Y(inst_cellmath__28), .A(N2988), .B(N2992));
NOR2XL inst_cellmath__49_0_I5276 (.Y(inst_cellmath__31), .A(N3010), .B(N3014));
AOI22XL inst_cellmath__49_0_I5277 (.Y(N10167), .A0(N3328), .A1(N3350), .B0(N513), .B1(inst_cellmath__44[8]));
AOI22XL inst_cellmath__49_0_I5278 (.Y(N10128), .A0(inst_cellmath__44[8]), .A1(N514), .B0(N3350), .B1(N3337));
AOI22XL inst_cellmath__49_0_I5279 (.Y(N10141), .A0(inst_cellmath__44[8]), .A1(N515), .B0(N3350), .B1(N3345));
AOI22XL inst_cellmath__49_0_I5280 (.Y(N10152), .A0(inst_cellmath__44[8]), .A1(N516), .B0(N3350), .B1(N3353));
AOI22XL inst_cellmath__49_0_I5281 (.Y(N10162), .A0(N3437), .A1(N3495), .B0(N3470), .B1(N3474));
AOI22XL inst_cellmath__49_0_I5282 (.Y(N3485), .A0(N3437), .A1(N3453), .B0(N3433), .B1(N3470));
AOI22X1 inst_cellmath__49_0_I5283 (.Y(N3445), .A0(N3437), .A1(N3412), .B0(N3392), .B1(N3470));
INVXL inst_cellmath__49_0_I5382 (.Y(N10324), .A(N10367));
AOI22XL inst_cellmath__49_0_I5395 (.Y(N10363), .A0(N3526), .A1(N3531), .B0(N3459), .B1(N10346));
AOI22X1 inst_cellmath__49_0_I5403 (.Y(N10369), .A0(N3437), .A1(N10363), .B0(N3508), .B1(N3470));
AOI22X1 inst_cellmath__49_0_I5404 (.Y(N3521), .A0(N3466), .A1(N3470), .B0(N3437), .B1(N3487));
AO22X1 inst_cellmath__49_0_I5405 (.Y(N3381), .A0(N10339), .A1(inst_cellmath__44[8]), .B0(N10324), .B1(N3350));
INVX1 inst_cellmath__49_0_I5406 (.Y(N3415), .A(N3381));
AOI22XL inst_cellmath__49_0_I5407 (.Y(N3400), .A0(N3381), .A1(N10369), .B0(N3521), .B1(N3415));
AND2XL inst_cellmath__49_0_I5428 (.Y(N10157), .A(N3415), .B(N3485));
INVXL inst_cellmath__49_0_I5291 (.Y(N3484), .A(N10167));
INVX1 inst_cellmath__49_0_I5292 (.Y(N3520), .A(N3484));
AOI211X1 inst_cellmath__49_0_I5430 (.Y(N10144), .A0(N3381), .A1(N10162), .B0(N10167), .C0(N10157));
AOI21X1 inst_cellmath__49_0_I5294 (.Y(N10124), .A0(N3381), .A1(N3445), .B0(N3484));
NOR3X1 inst_cellmath__49_0_I5295 (.Y(N3704), .A(N10141), .B(N10128), .C(N10152));
NOR2X1 inst_cellmath__49_0_I5296 (.Y(N3772), .A(inst_cellmath__31), .B(inst_cellmath__28));
AND2XL inst_cellmath__49_0_I5297 (.Y(N522), .A(N3772), .B(N3704));
NAND2X1 inst_cellmath__49_0_I5298 (.Y(N10133), .A(N3772), .B(N3704));
NOR3X1 inst_cellmath__49_0_I5299 (.Y(inst_cellmath__39[1]), .A(N10133), .B(N10124), .C(N10144));
AOI22X1 inst_cellmath__49_0_I629 (.Y(N3488), .A0(N3415), .A1(N3452), .B0(N3494), .B1(N3381));
AOI22XL inst_cellmath__49_0_I632 (.Y(N3435), .A0(N3415), .A1(N3397), .B0(N3438), .B1(N3381));
AOI22XL inst_cellmath__49_0_I633 (.Y(N3468), .A0(N3415), .A1(N3432), .B0(N3472), .B1(N3381));
AOI22XL inst_cellmath__49_0_I634 (.Y(N3504), .A0(N3415), .A1(N3465), .B0(N3507), .B1(N3381));
AOI22XL inst_cellmath__49_0_I635 (.Y(N3379), .A0(N3415), .A1(N3501), .B0(N3385), .B1(N3381));
AOI22XL inst_cellmath__49_0_I636 (.Y(N3413), .A0(N3415), .A1(N3376), .B0(N3418), .B1(N3381));
AOI22XL inst_cellmath__49_0_I637 (.Y(N3448), .A0(N3415), .A1(N3410), .B0(N3452), .B1(N3381));
AOI22XL inst_cellmath__49_0_I638 (.Y(N3482), .A0(N3415), .A1(N3445), .B0(N3485), .B1(N3381));
AOI22XL inst_cellmath__49_0_I639 (.Y(N3518), .A0(N3415), .A1(N3479), .B0(N3521), .B1(N3381));
AOI22XL inst_cellmath__49_0_I640 (.Y(N3394), .A0(N3415), .A1(N3515), .B0(N3397), .B1(N3381));
AOI22XL inst_cellmath__49_0_I641 (.Y(N3429), .A0(N3415), .A1(N3391), .B0(N3432), .B1(N3381));
AOI22XL inst_cellmath__49_0_I642 (.Y(N3462), .A0(N3415), .A1(N3426), .B0(N3465), .B1(N3381));
AOI22XL inst_cellmath__49_0_I643 (.Y(N3498), .A0(N3415), .A1(N3533), .B0(N3501), .B1(N3381));
AOI22XL inst_cellmath__49_0_I644 (.Y(N3535), .A0(N3415), .A1(N3476), .B0(N3376), .B1(N3381));
AOI22X1 inst_cellmath__49_0_I645 (.Y(N3408), .A0(N3415), .A1(N3422), .B0(N3410), .B1(N3381));
NAND2XL inst_cellmath__49_0_I647 (.Y(N3511), .A(N3479), .B(N3381));
NAND2XL inst_cellmath__49_0_I648 (.Y(N3423), .A(N3515), .B(N3381));
NAND2XL inst_cellmath__49_0_I649 (.Y(N3492), .A(N3391), .B(N3381));
NAND2XL inst_cellmath__49_0_I650 (.Y(N3402), .A(N3426), .B(N3381));
NAND2XL inst_cellmath__49_0_I651 (.Y(N3471), .A(N3533), .B(N3381));
NAND2XL inst_cellmath__49_0_I652 (.Y(N3383), .A(N3476), .B(N3381));
NAND2XL inst_cellmath__49_0_I653 (.Y(N3450), .A(N3422), .B(N3381));
AOI22X1 inst_cellmath__49_0_I656 (.Y(inst_cellmath__49[0]), .A0(N3484), .A1(N3488), .B0(N3408), .B1(N3520));
AOI22XL inst_cellmath__49_0_I658 (.Y(inst_cellmath__49[2]), .A0(N3484), .A1(N3400), .B0(N3511), .B1(N3520));
AOI22XL inst_cellmath__49_0_I659 (.Y(inst_cellmath__49[3]), .A0(N3484), .A1(N3435), .B0(N3423), .B1(N3520));
AOI22XL inst_cellmath__49_0_I660 (.Y(inst_cellmath__49[4]), .A0(N3484), .A1(N3468), .B0(N3492), .B1(N3520));
AOI22XL inst_cellmath__49_0_I661 (.Y(inst_cellmath__49[5]), .A0(N3484), .A1(N3504), .B0(N3402), .B1(N3520));
AOI22XL inst_cellmath__49_0_I662 (.Y(inst_cellmath__49[6]), .A0(N3484), .A1(N3379), .B0(N3471), .B1(N3520));
AOI22XL inst_cellmath__49_0_I663 (.Y(inst_cellmath__49[7]), .A0(N3484), .A1(N3413), .B0(N3383), .B1(N3520));
AOI22XL inst_cellmath__49_0_I664 (.Y(inst_cellmath__49[8]), .A0(N3484), .A1(N3448), .B0(N3450), .B1(N3520));
NAND3XL hyperpropagate_4_1_A_I5474 (.Y(N10423), .A(N3381), .B(N3704), .C(N3445));
NOR2XL hyperpropagate_4_1_A_I5475 (.Y(N539), .A(N3520), .B(N10423));
AND2X1 cynw_cm_float_add2_I708 (.Y(inst_cellmath__39[0]), .A(N522), .B(inst_cellmath__49[0]));
AND3XL cynw_cm_float_add2_I2090 (.Y(inst_cellmath__39[2]), .A(N3772), .B(N3704), .C(inst_cellmath__49[2]));
AND3XL cynw_cm_float_add2_I2091 (.Y(inst_cellmath__39[3]), .A(N3772), .B(N3704), .C(inst_cellmath__49[3]));
AND3XL cynw_cm_float_add2_I2092 (.Y(inst_cellmath__39[4]), .A(N3772), .B(N3704), .C(inst_cellmath__49[4]));
AND3XL cynw_cm_float_add2_I2093 (.Y(inst_cellmath__39[5]), .A(N3772), .B(inst_cellmath__49[5]), .C(N3704));
AND3XL cynw_cm_float_add2_I2094 (.Y(inst_cellmath__39[6]), .A(N3772), .B(inst_cellmath__49[6]), .C(N3704));
AND3XL cynw_cm_float_add2_I2095 (.Y(inst_cellmath__39[7]), .A(N3772), .B(inst_cellmath__49[7]), .C(N3704));
AND3XL cynw_cm_float_add2_I2096 (.Y(inst_cellmath__39[8]), .A(N3772), .B(inst_cellmath__49[8]), .C(N3704));
NOR4BBX1 cynw_cm_float_add2_I2097 (.Y(inst_cellmath__39[9]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3482));
NOR4BBX1 cynw_cm_float_add2_I2098 (.Y(inst_cellmath__39[10]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3518));
NOR4BBX1 cynw_cm_float_add2_I2099 (.Y(inst_cellmath__39[11]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3394));
NOR4BBX1 cynw_cm_float_add2_I2100 (.Y(inst_cellmath__39[12]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3429));
NOR4BBX1 cynw_cm_float_add2_I2101 (.Y(inst_cellmath__39[13]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3462));
NOR4BBX1 cynw_cm_float_add2_I2102 (.Y(inst_cellmath__39[14]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3498));
NOR4BBX1 cynw_cm_float_add2_I2103 (.Y(inst_cellmath__39[15]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3535));
NOR4BBX1 cynw_cm_float_add2_I2104 (.Y(inst_cellmath__39[16]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3408));
AND2XL cynw_cm_float_add2_I725 (.Y(inst_cellmath__39[17]), .A(N3772), .B(N539));
NOR4BBX1 cynw_cm_float_add2_I2106 (.Y(inst_cellmath__39[18]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3511));
NOR4BBX1 cynw_cm_float_add2_I2107 (.Y(inst_cellmath__39[19]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3423));
NOR4BBX1 cynw_cm_float_add2_I2108 (.Y(inst_cellmath__39[20]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3492));
NOR4BBX1 cynw_cm_float_add2_I2109 (.Y(inst_cellmath__39[21]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3402));
NOR4BBX1 cynw_cm_float_add2_I2110 (.Y(inst_cellmath__39[22]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3471));
NOR4BBX1 cynw_cm_float_add2_I2111 (.Y(inst_cellmath__39[23]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3383));
NOR4BBX1 cynw_cm_float_add2_I2112 (.Y(inst_cellmath__39[24]), .AN(N3704), .BN(N3772), .C(N3520), .D(N3450));
INVX1 inst_cellmath__55_2mx_I733 (.Y(inst_cellmath__55[24]), .A(inst_cellmath__55[0]));
XNOR2X1 inst_cellmath__55_2mx_I734 (.Y(inst_cellmath__55[1]), .A(N575), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I735 (.Y(inst_cellmath__55[2]), .A(N576), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I736 (.Y(inst_cellmath__55[3]), .A(N577), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I737 (.Y(inst_cellmath__55[4]), .A(N578), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I738 (.Y(inst_cellmath__55[5]), .A(N579), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I739 (.Y(inst_cellmath__55[6]), .A(N580), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I740 (.Y(inst_cellmath__55[7]), .A(N581), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I741 (.Y(inst_cellmath__55[8]), .A(N582), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I742 (.Y(inst_cellmath__55[9]), .A(N583), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I743 (.Y(inst_cellmath__55[10]), .A(N584), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I744 (.Y(inst_cellmath__55[11]), .A(N585), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I745 (.Y(inst_cellmath__55[12]), .A(N586), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I746 (.Y(inst_cellmath__55[13]), .A(N587), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I747 (.Y(inst_cellmath__55[14]), .A(N588), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I748 (.Y(inst_cellmath__55[15]), .A(N589), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I749 (.Y(inst_cellmath__55[16]), .A(N590), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I750 (.Y(inst_cellmath__55[17]), .A(N591), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I751 (.Y(inst_cellmath__55[18]), .A(N592), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I752 (.Y(inst_cellmath__55[19]), .A(N593), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I753 (.Y(inst_cellmath__55[20]), .A(N594), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I754 (.Y(inst_cellmath__55[21]), .A(N595), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I755 (.Y(inst_cellmath__55[22]), .A(N596), .B(inst_cellmath__55[24]));
XNOR2X1 inst_cellmath__55_2mx_I756 (.Y(inst_cellmath__55[23]), .A(N597), .B(inst_cellmath__55[24]));
ADDHX1 inst_cellmath__57__22__I757 (.CO(N4035), .S(N445), .A(inst_cellmath__55[0]), .B(inst_cellmath__39[0]));
ADDFXL inst_cellmath__57__22__I758 (.CO(N4015), .S(N446), .A(inst_cellmath__39[1]), .B(inst_cellmath__55[1]), .CI(N4035));
ADDFXL inst_cellmath__57__22__I759 (.CO(N3930), .S(N447), .A(inst_cellmath__39[2]), .B(inst_cellmath__55[2]), .CI(N4015));
ADDFXL inst_cellmath__57__22__I760 (.CO(N3996), .S(N448), .A(inst_cellmath__39[3]), .B(inst_cellmath__55[3]), .CI(N3930));
ADDFHXL inst_cellmath__57__22__I761 (.CO(N3911), .S(N449), .A(inst_cellmath__39[4]), .B(inst_cellmath__55[4]), .CI(N3996));
ADDFHXL inst_cellmath__57__22__I762 (.CO(N3977), .S(N450), .A(inst_cellmath__39[5]), .B(inst_cellmath__55[5]), .CI(N3911));
ADDFHXL inst_cellmath__57__22__I763 (.CO(N4043), .S(N451), .A(inst_cellmath__39[6]), .B(inst_cellmath__55[6]), .CI(N3977));
ADDFHXL inst_cellmath__57__22__I764 (.CO(N3957), .S(N452), .A(inst_cellmath__39[7]), .B(inst_cellmath__55[7]), .CI(N4043));
ADDFHXL inst_cellmath__57__22__I765 (.CO(N4023), .S(N453), .A(inst_cellmath__39[8]), .B(inst_cellmath__55[8]), .CI(N3957));
ADDFHXL inst_cellmath__57__22__I766 (.CO(N3938), .S(N454), .A(inst_cellmath__39[9]), .B(inst_cellmath__55[9]), .CI(N4023));
ADDFHXL inst_cellmath__57__22__I767 (.CO(N4004), .S(N455), .A(inst_cellmath__39[10]), .B(inst_cellmath__55[10]), .CI(N3938));
ADDFHXL inst_cellmath__57__22__I768 (.CO(N3919), .S(N456), .A(inst_cellmath__39[11]), .B(inst_cellmath__55[11]), .CI(N4004));
ADDFHXL inst_cellmath__57__22__I769 (.CO(N3985), .S(N457), .A(inst_cellmath__39[12]), .B(inst_cellmath__55[12]), .CI(N3919));
ADDFHXL inst_cellmath__57__22__I770 (.CO(N3900), .S(N458), .A(inst_cellmath__39[13]), .B(inst_cellmath__55[13]), .CI(N3985));
ADDFHXL inst_cellmath__57__22__I771 (.CO(N3966), .S(N459), .A(inst_cellmath__39[14]), .B(inst_cellmath__55[14]), .CI(N3900));
ADDFHXL inst_cellmath__57__22__I772 (.CO(N4032), .S(N460), .A(inst_cellmath__39[15]), .B(inst_cellmath__55[15]), .CI(N3966));
ADDFHXL inst_cellmath__57__22__I773 (.CO(N3947), .S(N461), .A(inst_cellmath__39[16]), .B(inst_cellmath__55[16]), .CI(N4032));
ADDFHXL inst_cellmath__57__22__I774 (.CO(N4012), .S(N462), .A(inst_cellmath__39[17]), .B(inst_cellmath__55[17]), .CI(N3947));
ADDFHXL inst_cellmath__57__22__I775 (.CO(N3927), .S(N463), .A(inst_cellmath__39[18]), .B(inst_cellmath__55[18]), .CI(N4012));
ADDFHXL inst_cellmath__57__22__I776 (.CO(N3993), .S(N464), .A(inst_cellmath__39[19]), .B(inst_cellmath__55[19]), .CI(N3927));
ADDFHXL inst_cellmath__57__22__I777 (.CO(N3908), .S(N465), .A(inst_cellmath__39[20]), .B(inst_cellmath__55[20]), .CI(N3993));
ADDFHXL inst_cellmath__57__22__I778 (.CO(N3974), .S(N466), .A(inst_cellmath__39[21]), .B(inst_cellmath__55[21]), .CI(N3908));
ADDFHXL inst_cellmath__57__22__I779 (.CO(N4040), .S(N467), .A(inst_cellmath__39[22]), .B(inst_cellmath__55[22]), .CI(N3974));
ADDFXL inst_cellmath__57__22__I780 (.CO(N3954), .S(N468), .A(inst_cellmath__39[23]), .B(inst_cellmath__55[23]), .CI(N4040));
XOR3XL inst_cellmath__57__22__I1984 (.Y(N469), .A(inst_cellmath__55[24]), .B(inst_cellmath__39[24]), .C(N3954));
ADDFXL inst_cellmath__57__22__I783 (.CO(N4002), .S(N420), .A(inst_cellmath__55[1]), .B(inst_cellmath__55[0]), .CI(inst_cellmath__39[1]));
ADDFXL inst_cellmath__57__22__I784 (.CO(N3917), .S(N421), .A(inst_cellmath__39[2]), .B(inst_cellmath__55[2]), .CI(N4002));
ADDFXL inst_cellmath__57__22__I785 (.CO(N3983), .S(N422), .A(inst_cellmath__39[3]), .B(inst_cellmath__55[3]), .CI(N3917));
ADDFXL inst_cellmath__57__22__I786 (.CO(N4049), .S(N423), .A(inst_cellmath__39[4]), .B(inst_cellmath__55[4]), .CI(N3983));
ADDFXL inst_cellmath__57__22__I787 (.CO(N3963), .S(N424), .A(inst_cellmath__39[5]), .B(inst_cellmath__55[5]), .CI(N4049));
ADDFXL inst_cellmath__57__22__I788 (.CO(N4029), .S(N425), .A(inst_cellmath__39[6]), .B(inst_cellmath__55[6]), .CI(N3963));
ADDFXL inst_cellmath__57__22__I789 (.CO(N3944), .S(N426), .A(inst_cellmath__39[7]), .B(inst_cellmath__55[7]), .CI(N4029));
ADDFXL inst_cellmath__57__22__I790 (.CO(N4009), .S(N427), .A(inst_cellmath__39[8]), .B(inst_cellmath__55[8]), .CI(N3944));
ADDFXL inst_cellmath__57__22__I791 (.CO(N3924), .S(N428), .A(inst_cellmath__39[9]), .B(inst_cellmath__55[9]), .CI(N4009));
ADDFXL inst_cellmath__57__22__I792 (.CO(N3990), .S(N429), .A(inst_cellmath__39[10]), .B(inst_cellmath__55[10]), .CI(N3924));
ADDFXL inst_cellmath__57__22__I793 (.CO(N3905), .S(N430), .A(inst_cellmath__39[11]), .B(inst_cellmath__55[11]), .CI(N3990));
ADDFXL inst_cellmath__57__22__I794 (.CO(N3971), .S(N431), .A(inst_cellmath__39[12]), .B(inst_cellmath__55[12]), .CI(N3905));
ADDFXL inst_cellmath__57__22__I795 (.CO(N4037), .S(N432), .A(inst_cellmath__39[13]), .B(inst_cellmath__55[13]), .CI(N3971));
ADDFXL inst_cellmath__57__22__I796 (.CO(N3951), .S(N433), .A(inst_cellmath__39[14]), .B(inst_cellmath__55[14]), .CI(N4037));
ADDFXL inst_cellmath__57__22__I797 (.CO(N4017), .S(N434), .A(inst_cellmath__39[15]), .B(inst_cellmath__55[15]), .CI(N3951));
ADDFXL inst_cellmath__57__22__I798 (.CO(N3932), .S(N435), .A(inst_cellmath__39[16]), .B(inst_cellmath__55[16]), .CI(N4017));
ADDFXL inst_cellmath__57__22__I799 (.CO(N3999), .S(N436), .A(inst_cellmath__39[17]), .B(inst_cellmath__55[17]), .CI(N3932));
ADDFXL inst_cellmath__57__22__I800 (.CO(N3913), .S(N437), .A(inst_cellmath__39[18]), .B(inst_cellmath__55[18]), .CI(N3999));
ADDFXL inst_cellmath__57__22__I801 (.CO(N3980), .S(N438), .A(inst_cellmath__39[19]), .B(inst_cellmath__55[19]), .CI(N3913));
ADDFXL inst_cellmath__57__22__I802 (.CO(N4046), .S(N439), .A(inst_cellmath__39[20]), .B(inst_cellmath__55[20]), .CI(N3980));
ADDFXL inst_cellmath__57__22__I803 (.CO(N3959), .S(N440), .A(inst_cellmath__39[21]), .B(inst_cellmath__55[21]), .CI(N4046));
ADDFXL inst_cellmath__57__22__I804 (.CO(N4026), .S(N441), .A(inst_cellmath__39[22]), .B(inst_cellmath__55[22]), .CI(N3959));
ADDFXL inst_cellmath__57__22__I805 (.CO(N3941), .S(N442), .A(inst_cellmath__39[23]), .B(inst_cellmath__55[23]), .CI(N4026));
ADDFXL inst_cellmath__57__22__I806 (.CO(N444), .S(N443), .A(inst_cellmath__39[24]), .B(inst_cellmath__55[24]), .CI(N3941));
INVX2 cynw_cm_float_add2_I32 (.Y(inst_cellmath__56[25]), .A(N444));
INVX2 cynw_cm_float_add2_I2034 (.Y(N6142), .A(inst_cellmath__56[25]));
INVXL cynw_cm_float_add2_I2040 (.Y(N6148), .A(N6142));
INVXL cynw_cm_float_add2_I2039 (.Y(N6147), .A(N6142));
INVX2 cynw_cm_float_add2_I2038 (.Y(N6146), .A(N6142));
INVXL cynw_cm_float_add2_I2037 (.Y(N6145), .A(N6142));
INVX1 cynw_cm_float_add2_I2036 (.Y(N6144), .A(N6142));
INVX1 cynw_cm_float_add2_I2035 (.Y(N6143), .A(N6142));
NOR2BX1 cynw_cm_float_add2_I807 (.Y(N418), .AN(a_sign), .B(inst_cellmath__28));
NOR2BX1 cynw_cm_float_add2_I808 (.Y(N417), .AN(b_sign), .B(inst_cellmath__31));
AOI22XL inst_cellmath__52_0_I810 (.Y(N4164), .A0(N2888), .A1(N418), .B0(N417), .B1(N2842));
AOI22XL inst_cellmath__52_0_I811 (.Y(N4159), .A0(N2888), .A1(b_sign), .B0(a_sign), .B1(N2842));
MXI2XL inst_cellmath__52_0_I812 (.Y(inst_cellmath__52), .A(N4159), .B(N4164), .S0(N6148));
NOR2XL cynw_cm_float_add2_I813 (.Y(inst_cellmath__51[25]), .A(inst_cellmath__55[0]), .B(N6148));
MXI2XL inst_cellmath__51__24__I815 (.Y(N4259), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N445));
MXI2XL inst_cellmath__51__24__I816 (.Y(N4177), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N446));
MXI2XL inst_cellmath__51__24__I817 (.Y(N4200), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N447));
MXI2XL inst_cellmath__51__24__I818 (.Y(N4224), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N448));
MXI2XL inst_cellmath__51__24__I819 (.Y(N4247), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N449));
MXI2XL inst_cellmath__51__24__I820 (.Y(N4271), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N450));
MXI2XL inst_cellmath__51__24__I821 (.Y(N4188), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N451));
MXI2XL inst_cellmath__51__24__I822 (.Y(N4210), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N452));
MXI2XL inst_cellmath__51__24__I823 (.Y(N4234), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N453));
MXI2XL inst_cellmath__51__24__I824 (.Y(N4256), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N454));
MXI2XL inst_cellmath__51__24__I825 (.Y(N4280), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N455));
MXI2XL inst_cellmath__51__24__I826 (.Y(N4197), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N456));
MXI2XL inst_cellmath__51__24__I827 (.Y(N4220), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N457));
MXI2XL inst_cellmath__51__24__I828 (.Y(N4242), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N458));
MXI2XL inst_cellmath__51__24__I829 (.Y(N4267), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N459));
MXI2XL inst_cellmath__51__24__I830 (.Y(N4184), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N460));
MXI2XL inst_cellmath__51__24__I831 (.Y(N4206), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N461));
MXI2XL inst_cellmath__51__24__I832 (.Y(N4230), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N462));
MXI2XL inst_cellmath__51__24__I833 (.Y(N4252), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N463));
MXI2XL inst_cellmath__51__24__I834 (.Y(N4276), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N464));
MXI2XL inst_cellmath__51__24__I835 (.Y(N4193), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N465));
MXI2XL inst_cellmath__51__24__I836 (.Y(N4216), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N466));
MXI2XL inst_cellmath__51__24__I837 (.Y(N4239), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N467));
MXI2XL inst_cellmath__51__24__I838 (.Y(N4263), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N468));
MXI2XL inst_cellmath__51__24__I839 (.Y(N4180), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N469));
INVX2 inst_cellmath__51__24__I840 (.Y(N4226), .A(inst_cellmath__56[25]));
INVX2 inst_cellmath__51__24__I2041 (.Y(N6149), .A(N4226));
INVX2 inst_cellmath__51__24__I2042 (.Y(N6150), .A(N6149));
BUFX3 inst_cellmath__51__24__I5450 (.Y(N6152), .A(N4226));
AOI22XL inst_cellmath__51__24__I841 (.Y(N470), .A0(N6152), .A1(inst_cellmath__39[0]), .B0(N4259), .B1(N6147));
AOI22XL inst_cellmath__51__24__I842 (.Y(N471), .A0(N6152), .A1(N420), .B0(N4177), .B1(N6147));
AOI22X1 inst_cellmath__51__24__I844 (.Y(N473), .A0(N422), .A1(N6152), .B0(N4224), .B1(N6147));
AOI22XL inst_cellmath__51__24__I845 (.Y(N474), .A0(N6152), .A1(N423), .B0(N4247), .B1(N6147));
AOI22X1 inst_cellmath__51__24__I846 (.Y(N475), .A0(N6152), .A1(N424), .B0(N4271), .B1(N6147));
AOI22X1 inst_cellmath__51__24__I848 (.Y(N477), .A0(N426), .A1(N6150), .B0(N4210), .B1(N6146));
AOI22X1 inst_cellmath__51__24__I849 (.Y(N478), .A0(N427), .A1(N6150), .B0(N4234), .B1(N6146));
AOI22X1 inst_cellmath__51__24__I850 (.Y(N479), .A0(N428), .A1(N6150), .B0(N4256), .B1(N6146));
AOI22XL inst_cellmath__51__24__I853 (.Y(N482), .A0(N6152), .A1(N431), .B0(N4220), .B1(N6145));
AOI22X1 inst_cellmath__51__24__I854 (.Y(N483), .A0(N6152), .A1(N432), .B0(N4242), .B1(N6145));
AOI22X1 inst_cellmath__51__24__I856 (.Y(N485), .A0(N434), .A1(N6150), .B0(N4184), .B1(N6145));
AOI22X1 inst_cellmath__51__24__I859 (.Y(N488), .A0(N6152), .A1(N437), .B0(N4252), .B1(N6145));
AOI22X1 inst_cellmath__51__24__I864 (.Y(N493), .A0(N442), .A1(N6150), .B0(N4263), .B1(N6144));
INVXL cynw_cm_float_add2_I38 (.Y(inst_cellmath__51[0]), .A(N470));
INVXL cynw_cm_float_add2_I39 (.Y(inst_cellmath__51[1]), .A(N471));
AO22XL cynw_cm_float_add2_I2024 (.Y(inst_cellmath__51[2]), .A0(N4200), .A1(N6143), .B0(N6152), .B1(N421));
INVX1 cynw_cm_float_add2_I41 (.Y(inst_cellmath__51[3]), .A(N473));
INVX1 cynw_cm_float_add2_I42 (.Y(inst_cellmath__51[4]), .A(N474));
INVX1 cynw_cm_float_add2_I43 (.Y(inst_cellmath__51[5]), .A(N475));
AO22X1 cynw_cm_float_add2_I2063 (.Y(inst_cellmath__51[6]), .A0(N4188), .A1(N6146), .B0(N425), .B1(N6152));
INVX1 cynw_cm_float_add2_I45 (.Y(inst_cellmath__51[7]), .A(N477));
INVX1 cynw_cm_float_add2_I46 (.Y(inst_cellmath__51[8]), .A(N478));
INVX1 cynw_cm_float_add2_I47 (.Y(inst_cellmath__51[9]), .A(N479));
AOI22X1 cynw_cm_float_add2_I2054 (.Y(N6165), .A0(N4267), .A1(N6143), .B0(N6150), .B1(N433));
INVX1 cynw_cm_float_add2_I56 (.Y(inst_cellmath__51[18]), .A(N488));
AO22XL cynw_cm_float_add2_I1998 (.Y(inst_cellmath__51[19]), .A0(N4276), .A1(N6144), .B0(N6150), .B1(N438));
AO22XL cynw_cm_float_add2_I2058 (.Y(inst_cellmath__51[20]), .A0(N4193), .A1(N6145), .B0(N6152), .B1(N439));
AO22XL cynw_cm_float_add2_I2026 (.Y(inst_cellmath__51[21]), .A0(N4216), .A1(N6143), .B0(N6150), .B1(N440));
AOI22X1 cynw_cm_float_add2_I2059 (.Y(N6173), .A0(N4239), .A1(N6143), .B0(N6150), .B1(N441));
INVX1 cynw_cm_float_add2_I2060 (.Y(inst_cellmath__51[22]), .A(N6173));
INVX1 cynw_cm_float_add2_I61 (.Y(inst_cellmath__51[23]), .A(N493));
AO22X1 cynw_cm_float_add2_I1985 (.Y(inst_cellmath__51[24]), .A0(N4180), .A1(N6144), .B0(N443), .B1(N6150));
NOR2XL inst_delta_0_I867 (.Y(N4402), .A(inst_cellmath__51[1]), .B(inst_cellmath__51[0]));
NOR2BX1 inst_delta_0_I868 (.Y(N4349), .AN(inst_cellmath__51[2]), .B(inst_cellmath__51[3]));
INVXL inst_delta_0_I869 (.Y(N4368), .A(inst_cellmath__51[5]));
OAI21XL inst_delta_0_I870 (.Y(N4390), .A0(inst_cellmath__51[4]), .A1(N4349), .B0(N4368));
NOR2X1 inst_delta_0_I871 (.Y(N4412), .A(inst_cellmath__51[3]), .B(inst_cellmath__51[2]));
NOR2X1 inst_delta_0_I872 (.Y(N4336), .A(inst_cellmath__51[5]), .B(inst_cellmath__51[4]));
NOR2BX1 inst_delta_0_I873 (.Y(N4378), .AN(inst_cellmath__51[6]), .B(inst_cellmath__51[7]));
INVXL inst_delta_0_I874 (.Y(N4398), .A(inst_cellmath__51[9]));
OAI21X1 inst_delta_0_I875 (.Y(N4421), .A0(inst_cellmath__51[8]), .A1(N4378), .B0(N4398));
NOR2X1 inst_delta_0_I876 (.Y(N4345), .A(inst_cellmath__51[7]), .B(inst_cellmath__51[6]));
NOR2X1 inst_delta_0_I877 (.Y(N4364), .A(inst_cellmath__51[9]), .B(inst_cellmath__51[8]));
AO22XL inst_cellmath__66_0_I5435 (.Y(inst_cellmath__51[10]), .A0(N4280), .A1(N6146), .B0(N429), .B1(N6152));
AO22X1 inst_cellmath__66_0_I5356 (.Y(inst_cellmath__51[11]), .A0(N4197), .A1(N6143), .B0(N430), .B1(N6152));
NOR2BX1 inst_delta_0_I878 (.Y(N4408), .AN(inst_cellmath__51[10]), .B(inst_cellmath__51[11]));
INVX1 inst_cellmath__66_0_I5354 (.Y(inst_cellmath__51[13]), .A(N483));
INVXL inst_delta_0_I879 (.Y(N4428), .A(inst_cellmath__51[13]));
INVX1 inst_cellmath__66_0_I5353 (.Y(inst_cellmath__51[12]), .A(N482));
OAI21X1 inst_delta_0_I880 (.Y(N4355), .A0(inst_cellmath__51[12]), .A1(N4408), .B0(N4428));
INVX1 inst_cellmath__66_0_I5359 (.Y(inst_cellmath__51[14]), .A(N6165));
INVX1 inst_cellmath__66_0_I5355 (.Y(inst_cellmath__51[15]), .A(N485));
NOR2BX1 inst_delta_0_I883 (.Y(N4341), .AN(inst_cellmath__51[14]), .B(inst_cellmath__51[15]));
AO22X1 inst_cellmath__66_0_I5361 (.Y(inst_cellmath__51[17]), .A0(N4230), .A1(N6144), .B0(N6150), .B1(N436));
INVXL inst_delta_0_I884 (.Y(N4362), .A(inst_cellmath__51[17]));
AO22X1 inst_cellmath__66_0_I5362 (.Y(inst_cellmath__51[16]), .A0(N4206), .A1(N6144), .B0(N6150), .B1(N435));
OAI21X1 inst_delta_0_I885 (.Y(N4383), .A0(inst_cellmath__51[16]), .A1(N4341), .B0(N4362));
NOR2BX1 inst_delta_0_I888 (.Y(N4370), .AN(inst_cellmath__51[18]), .B(inst_cellmath__51[19]));
INVXL inst_delta_0_I889 (.Y(N4392), .A(inst_cellmath__51[21]));
OAI21XL inst_delta_0_I890 (.Y(N4414), .A0(inst_cellmath__51[20]), .A1(N4370), .B0(N4392));
NOR2XL inst_delta_0_I891 (.Y(N4338), .A(inst_cellmath__51[19]), .B(inst_cellmath__51[18]));
NOR2X1 inst_delta_0_I892 (.Y(N4359), .A(inst_cellmath__51[21]), .B(inst_cellmath__51[20]));
NOR2BX1 inst_delta_0_I893 (.Y(N4400), .AN(inst_cellmath__51[22]), .B(inst_cellmath__51[23]));
INVXL inst_delta_0_I894 (.Y(N4423), .A(inst_cellmath__51[25]));
OAI21XL inst_delta_0_I895 (.Y(N4347), .A0(inst_cellmath__51[24]), .A1(N4400), .B0(N4423));
NOR2X1 inst_delta_0_I896 (.Y(N4366), .A(inst_cellmath__51[23]), .B(inst_cellmath__51[22]));
NOR2X2 inst_delta_0_I897 (.Y(N4388), .A(inst_cellmath__51[25]), .B(inst_cellmath__51[24]));
NAND2BXL inst_delta_0_I898 (.Y(N4384), .AN(N4412), .B(N4336));
NAND2X1 inst_delta_0_I899 (.Y(N4352), .A(N4336), .B(N4412));
NAND2X1 inst_delta_0_I900 (.Y(N4371), .A(N4364), .B(N4345));
NOR2X1 inst_cellmath__66_0_I5357 (.Y(N4375), .A(inst_cellmath__51[11]), .B(inst_cellmath__51[10]));
NOR2X1 inst_cellmath__66_0_I5358 (.Y(N4395), .A(inst_cellmath__51[13]), .B(inst_cellmath__51[12]));
NAND2BXL inst_delta_0_I901 (.Y(N4415), .AN(N4375), .B(N4395));
NOR2X1 inst_cellmath__66_0_I5363 (.Y(N4426), .A(inst_cellmath__51[17]), .B(inst_cellmath__51[16]));
INVXL inst_delta_0_I902 (.Y(N4339), .A(N4426));
NOR2X1 inst_cellmath__66_0_I5360 (.Y(N4405), .A(inst_cellmath__51[14]), .B(inst_cellmath__51[15]));
AOI21XL inst_delta_0_I903 (.Y(N4360), .A0(N4405), .A1(N4415), .B0(N4339));
NAND2BXL inst_delta_0_I906 (.Y(N4348), .AN(N4338), .B(N4359));
INVXL inst_delta_0_I907 (.Y(N4367), .A(N4388));
AOI21XL inst_delta_0_I908 (.Y(N4389), .A0(N4366), .A1(N4348), .B0(N4367));
NAND2X1 inst_delta_0_I909 (.Y(N4411), .A(N4359), .B(N4338));
NAND2X2 inst_delta_0_I910 (.Y(N4335), .A(N4388), .B(N4366));
NAND2BXL inst_delta_0_I911 (.Y(N4420), .AN(N4371), .B(N4352));
NAND2X1 inst_cellmath__66_0_I5364 (.Y(N4380), .A(N4375), .B(N4395));
NAND2X1 inst_cellmath__66_0_I5365 (.Y(N4401), .A(N4426), .B(N4405));
NOR2BX1 inst_delta_0_I913 (.Y(N4354), .AN(N4380), .B(N4401));
INVXL inst_delta_0_I914 (.Y(N4374), .A(N4335));
OAI21XL inst_delta_0_I915 (.Y(N4393), .A0(N4411), .A1(N4354), .B0(N4374));
NOR2X1 inst_cellmath__66_0_I5302 (.Y(N4407), .A(N4371), .B(N4352));
NAND2BXL inst_delta_0_I918 (.Y(N4382), .AN(N4402), .B(N4407));
NOR2X2 inst_cellmath__66_0_I5304 (.Y(N4372), .A(N4335), .B(N4411));
INVXL inst_delta_0_I919 (.Y(N4404), .A(N4372));
NOR2X1 inst_cellmath__66_0_I5366 (.Y(N4418), .A(N4401), .B(N4380));
AOI21XL inst_delta_0_I920 (.Y(inst_delta[3]), .A0(N4418), .A1(N4382), .B0(N4404));
NAND2XL inst_delta_0_I921 (.Y(N4351), .A(N4407), .B(N4402));
NAND2X2 inst_cellmath__66_0_I5305 (.Y(N4417), .A(N4418), .B(N4372));
NOR2BX1 inst_delta_0_I923 (.Y(inst_delta[4]), .AN(N4351), .B(N4417));
NOR2XL inst_delta_0_I924 (.Y(inst_delta[5]), .A(N4417), .B(N4351));
OAI21XL inst_delta_0_I925 (.Y(inst_delta[2]), .A0(N4417), .A1(N4420), .B0(N4393));
OAI2BB1X1 inst_delta_0_I926 (.Y(N4376), .A0N(N4345), .A1N(N4384), .B0(N4364));
AOI21XL inst_delta_0_I927 (.Y(N4342), .A0(N4372), .A1(N4360), .B0(N4389));
NOR2BX1 cynw_cm_float_add2_I935 (.Y(N496), .AN(inst_cellmath__52), .B(inst_delta[5]));
AO21XL cynw_cm_float_add2_I2128 (.Y(inst_cellmath__69), .A0(a_sign), .A1(b_sign), .B0(N496));
NOR2BX1 cynw_cm_float_add2_I938 (.Y(x[31]), .AN(inst_cellmath__69), .B(inst_cellmath__62));
MX2XL cynw_cm_float_add2_I941 (.Y(inst_cellmath__40[0]), .A(N10019), .B(b_exp[0]), .S0(N2914));
MX2XL cynw_cm_float_add2_I942 (.Y(inst_cellmath__40[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(N2914));
MX2XL cynw_cm_float_add2_I943 (.Y(inst_cellmath__40[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(N2914));
MX2XL cynw_cm_float_add2_I944 (.Y(inst_cellmath__40[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(N2914));
MX2XL cynw_cm_float_add2_I945 (.Y(inst_cellmath__40[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(N2914));
MX2XL cynw_cm_float_add2_I946 (.Y(inst_cellmath__40[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(N2914));
MX2XL cynw_cm_float_add2_I947 (.Y(inst_cellmath__40[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(N2914));
MX2XL cynw_cm_float_add2_I948 (.Y(inst_cellmath__40[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(N2914));
INVXL inst_cellmath__73_0_I949 (.Y(N4571), .A(inst_cellmath__40[2]));
INVXL inst_cellmath__73_0_I950 (.Y(N4566), .A(inst_cellmath__40[4]));
NOR2BX1 inst_cellmath__66_0_I5301 (.Y(N10217), .AN(inst_cellmath__51[0]), .B(inst_cellmath__51[1]));
OAI21X1 inst_cellmath__66_0_I5306 (.Y(N10220), .A0(N4371), .A1(N4390), .B0(N4421));
AOI21X1 inst_cellmath__66_0_I5309 (.Y(N10209), .A0(N10217), .A1(N4407), .B0(N10220));
OAI21X1 inst_cellmath__66_0_I5307 (.Y(N10197), .A0(N4355), .A1(N4401), .B0(N4383));
OAI21X1 inst_cellmath__66_0_I5308 (.Y(N10202), .A0(N4335), .A1(N4414), .B0(N4347));
AOI21XL inst_cellmath__66_0_I5312 (.Y(N10216), .A0(N10197), .A1(N4372), .B0(N10202));
OAI21XL inst_cellmath__66_0_I5436 (.Y(inst_delta[0]), .A0(N4417), .A1(N10209), .B0(N10216));
NAND2BXL inst_cellmath__73_0_I951 (.Y(N4578), .AN(inst_cellmath__40[0]), .B(inst_delta[0]));
OA21X1 inst_cellmath__73_0_I1988 (.Y(N4569), .A0(N4376), .A1(N4417), .B0(N4342));
BUFX6 inst_cellmath__73_0_I2129 (.Y(N6154), .A(N4569));
AND2XL inst_cellmath__73_0_I953 (.Y(N4573), .A(inst_cellmath__40[1]), .B(N6154));
OAI22XL inst_cellmath__73_0_I954 (.Y(N4561), .A0(N4573), .A1(N4578), .B0(inst_cellmath__40[1]), .B1(N6154));
OR2XL inst_cellmath__73_0_I955 (.Y(N4557), .A(N4571), .B(inst_delta[2]));
AOI22XL inst_cellmath__73_0_I956 (.Y(N4567), .A0(N4561), .A1(N4557), .B0(N4571), .B1(inst_delta[2]));
INVXL inst_cellmath__73_0_I957 (.Y(N4565), .A(inst_delta[3]));
AND2XL inst_cellmath__73_0_I958 (.Y(N4570), .A(inst_cellmath__40[3]), .B(N4565));
OAI22XL inst_cellmath__73_0_I959 (.Y(N4575), .A0(N4570), .A1(N4567), .B0(inst_cellmath__40[3]), .B1(N4565));
OR2XL inst_cellmath__73_0_I960 (.Y(N4554), .A(N4566), .B(inst_delta[4]));
AOI22X1 inst_cellmath__73_0_I961 (.Y(N4552), .A0(N4575), .A1(N4554), .B0(N4566), .B1(inst_delta[4]));
NOR4X1 inst_cellmath__73_0_I962 (.Y(inst_cellmath__73), .A(inst_cellmath__40[7]), .B(inst_cellmath__40[6]), .C(inst_cellmath__40[5]), .D(N4552));
AND4XL inst_cellmath__75__32__I963 (.Y(N4603), .A(inst_cellmath__40[7]), .B(inst_cellmath__40[4]), .C(inst_cellmath__40[2]), .D(inst_cellmath__40[3]));
NAND2XL inst_cellmath__75__32__I964 (.Y(N4593), .A(N4603), .B(inst_cellmath__40[6]));
NAND3XL hyperpropagate_4_1_A_I2183 (.Y(N6205), .A(inst_cellmath__40[5]), .B(inst_cellmath__40[1]), .C(inst_cellmath__51[25]));
NOR2XL hyperpropagate_4_1_A_I2184 (.Y(N499), .A(N4593), .B(N6205));
OR4X1 cynw_cm_float_add2_I968 (.Y(inst_cellmath__77), .A(inst_cellmath__24), .B(inst_cellmath__21), .C(inst_cellmath__62), .D(N499));
AND2XL cynw_cm_float_add2_I969 (.Y(N498), .A(inst_cellmath__31), .B(inst_cellmath__28));
NOR4X6 cynw_cm_float_add2_I970 (.Y(inst_cellmath__72), .A(N498), .B(inst_cellmath__77), .C(inst_delta[5]), .D(inst_cellmath__73));
INVX1 inst_cellmath__66_0_I5310 (.Y(N10223), .A(N10202));
NAND2X1 inst_cellmath__66_0_I5311 (.Y(N10211), .A(N10197), .B(N4372));
NOR2X2 inst_cellmath__66_0_I5313 (.Y(N10208), .A(N10209), .B(N4417));
NAND2X2 inst_cellmath__66_0_I5316 (.Y(N10221), .A(N10223), .B(N10211));
NOR2X2 inst_cellmath__66_0_I5317 (.Y(N4645), .A(N10221), .B(N10208));
INVXL inst_cellmath__66_0_I973 (.Y(N4640), .A(inst_delta[2]));
INVXL buf1_A_I2185 (.Y(N6212), .A(N4640));
INVXL buf1_A_I2186 (.Y(N6161), .A(N6212));
INVXL inst_cellmath__66_0_I975 (.Y(N4635), .A(inst_delta[4]));
INVXL inst_cellmath__66_0_I976 (.Y(N4652), .A(inst_cellmath__40[1]));
ADDHX1 inst_cellmath__66_0_I977 (.CO(N4657), .S(N4644), .A(inst_cellmath__40[2]), .B(inst_cellmath__40[1]));
ADDHX1 inst_cellmath__66_0_I978 (.CO(N4632), .S(N4668), .A(inst_cellmath__40[3]), .B(N4657));
ADDHX1 inst_cellmath__66_0_I979 (.CO(N4650), .S(N4639), .A(inst_cellmath__40[4]), .B(N4632));
INVXL inst_cellmath__66_0_I980 (.Y(N4660), .A(inst_cellmath__40[5]));
INVXL inst_cellmath__66_0_I981 (.Y(N4654), .A(inst_cellmath__40[6]));
ADDHX1 inst_cellmath__66_0_I983 (.CO(N4653), .S(inst_cellmath__66[0]), .A(inst_cellmath__40[0]), .B(N4645));
ADDFXL inst_cellmath__66_0_I984 (.CO(N4646), .S(inst_cellmath__66[1]), .A(N4569), .B(N4652), .CI(N4653));
ADDFXL inst_cellmath__66_0_I985 (.CO(N4670), .S(inst_cellmath__66[2]), .A(N4640), .B(N4644), .CI(N4646));
ADDFXL inst_cellmath__66_0_I986 (.CO(N4641), .S(inst_cellmath__66[3]), .A(N4565), .B(N4668), .CI(N4670));
ADDFXL inst_cellmath__66_0_I987 (.CO(N4662), .S(inst_cellmath__66[4]), .A(N4635), .B(N4639), .CI(N4641));
ADDFXL inst_cellmath__66_0_I988 (.CO(N4636), .S(inst_cellmath__66[5]), .A(N4650), .B(N4660), .CI(N4662));
ADDFXL inst_cellmath__66_0_I989 (.CO(N4655), .S(inst_cellmath__66[6]), .A(N4654), .B(inst_cellmath__40[5]), .CI(N4636));
XNOR3XL inst_cellmath__66_0_I2022 (.Y(inst_cellmath__66[7]), .A(inst_cellmath__40[7]), .B(inst_cellmath__40[6]), .C(N4655));
MX2XL inst_cellmath__60_0_I991 (.Y(x[23]), .A(inst_cellmath__77), .B(inst_cellmath__66[0]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__60_0_I992 (.Y(x[24]), .A(inst_cellmath__77), .B(inst_cellmath__66[1]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__60_0_I993 (.Y(x[25]), .A(inst_cellmath__77), .B(inst_cellmath__66[2]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__60_0_I994 (.Y(x[26]), .A(inst_cellmath__77), .B(inst_cellmath__66[3]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__60_0_I995 (.Y(x[27]), .A(inst_cellmath__77), .B(inst_cellmath__66[4]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__60_0_I996 (.Y(x[28]), .A(inst_cellmath__77), .B(inst_cellmath__66[5]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__60_0_I997 (.Y(x[29]), .A(inst_cellmath__77), .B(inst_cellmath__66[6]), .S0(inst_cellmath__72));
INVXL mx2_A_I2187 (.Y(N6216), .A(inst_cellmath__72));
AO22XL mx2_A_I2188 (.Y(x[30]), .A0(inst_cellmath__77), .A1(N6216), .B0(inst_cellmath__66[7]), .B1(inst_cellmath__72));
INVXL inst_cellmath__63_0_I1000 (.Y(N4867), .A(inst_delta[3]));
AND2XL inst_cellmath__63_0_I1002 (.Y(N4856), .A(N4867), .B(inst_cellmath__51[0]));
AND2XL inst_cellmath__63_0_I1003 (.Y(N4760), .A(N4867), .B(inst_cellmath__51[1]));
AND2XL inst_cellmath__63_0_I1004 (.Y(N4833), .A(N4867), .B(inst_cellmath__51[2]));
AND2XL inst_cellmath__63_0_I1005 (.Y(N4736), .A(N4867), .B(inst_cellmath__51[3]));
AND2XL inst_cellmath__63_0_I1006 (.Y(N4814), .A(N4867), .B(inst_cellmath__51[4]));
AND2XL inst_cellmath__63_0_I1007 (.Y(N4887), .A(N4867), .B(inst_cellmath__51[5]));
AND2XL inst_cellmath__63_0_I1008 (.Y(N4790), .A(N4867), .B(inst_cellmath__51[6]));
AND2XL inst_cellmath__63_0_I1009 (.Y(N4866), .A(N4867), .B(inst_cellmath__51[7]));
MX2XL inst_cellmath__63_0_I1010 (.Y(N4769), .A(inst_cellmath__51[0]), .B(inst_cellmath__51[8]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1011 (.Y(N4807), .A(inst_cellmath__51[1]), .B(inst_cellmath__51[9]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1012 (.Y(N4842), .A(inst_cellmath__51[2]), .B(inst_cellmath__51[10]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1013 (.Y(N4881), .A(inst_cellmath__51[3]), .B(inst_cellmath__51[11]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1014 (.Y(N4746), .A(inst_cellmath__51[4]), .B(inst_cellmath__51[12]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1015 (.Y(N4784), .A(inst_cellmath__51[5]), .B(inst_cellmath__51[13]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1016 (.Y(N4822), .A(inst_cellmath__51[6]), .B(inst_cellmath__51[14]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1017 (.Y(N4859), .A(inst_cellmath__51[7]), .B(inst_cellmath__51[15]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1018 (.Y(N4895), .A(inst_cellmath__51[8]), .B(inst_cellmath__51[16]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1019 (.Y(N4763), .A(inst_cellmath__51[9]), .B(inst_cellmath__51[17]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1020 (.Y(N4799), .A(inst_cellmath__51[10]), .B(inst_cellmath__51[18]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1021 (.Y(N4836), .A(inst_cellmath__51[11]), .B(inst_cellmath__51[19]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1022 (.Y(N4875), .A(inst_cellmath__51[12]), .B(inst_cellmath__51[20]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1023 (.Y(N4741), .A(inst_cellmath__51[13]), .B(inst_cellmath__51[21]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1024 (.Y(N4779), .A(inst_cellmath__51[14]), .B(inst_cellmath__51[22]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1025 (.Y(N4818), .A(inst_cellmath__51[15]), .B(inst_cellmath__51[23]), .S0(N4867));
MX2XL inst_cellmath__63_0_I1026 (.Y(N4852), .A(inst_cellmath__51[16]), .B(inst_cellmath__51[24]), .S0(N4867));
NAND2XL inst_cellmath__63_0_I1029 (.Y(N4849), .A(N4856), .B(N4635));
NAND2XL inst_cellmath__63_0_I1030 (.Y(N4752), .A(N4760), .B(N4635));
NAND2XL inst_cellmath__63_0_I1031 (.Y(N4828), .A(N4833), .B(N4635));
NAND2XL inst_cellmath__63_0_I1032 (.Y(N4731), .A(N4736), .B(N4635));
NAND2XL inst_cellmath__63_0_I1033 (.Y(N4806), .A(N4814), .B(N4635));
NAND2XL inst_cellmath__63_0_I1034 (.Y(N4880), .A(N4887), .B(N4635));
NAND2XL inst_cellmath__63_0_I1035 (.Y(N4783), .A(N4790), .B(N4635));
NAND2XL inst_cellmath__63_0_I1036 (.Y(N4858), .A(N4866), .B(N4635));
NAND2XL inst_cellmath__63_0_I1037 (.Y(N4762), .A(N4769), .B(N4635));
NAND2XL inst_cellmath__63_0_I1038 (.Y(N4835), .A(N4807), .B(N4635));
NAND2XL inst_cellmath__63_0_I1039 (.Y(N4740), .A(N4842), .B(N4635));
NAND2XL inst_cellmath__63_0_I1040 (.Y(N4817), .A(N4881), .B(N4635));
NAND2XL inst_cellmath__63_0_I1041 (.Y(N4890), .A(N4746), .B(N4635));
NAND2XL inst_cellmath__63_0_I1042 (.Y(N4794), .A(N4784), .B(N4635));
NAND2XL inst_cellmath__63_0_I1043 (.Y(N4870), .A(N4822), .B(N4635));
NAND2XL inst_cellmath__63_0_I1044 (.Y(N4772), .A(N4859), .B(N4635));
AOI22XL inst_cellmath__63_0_I1045 (.Y(N4846), .A0(inst_delta[4]), .A1(N4856), .B0(N4895), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1046 (.Y(N4884), .A0(inst_delta[4]), .A1(N4760), .B0(N4763), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1047 (.Y(N4749), .A0(inst_delta[4]), .A1(N4833), .B0(N4799), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1048 (.Y(N4787), .A0(inst_delta[4]), .A1(N4736), .B0(N4836), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1049 (.Y(N4825), .A0(inst_delta[4]), .A1(N4814), .B0(N4875), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1050 (.Y(N4863), .A0(inst_delta[4]), .A1(N4887), .B0(N4741), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1051 (.Y(N4728), .A0(inst_delta[4]), .A1(N4790), .B0(N4779), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1052 (.Y(N4766), .A0(inst_delta[4]), .A1(N4866), .B0(N4818), .B1(N4635));
AOI22XL inst_cellmath__63_0_I1053 (.Y(N4803), .A0(inst_delta[4]), .A1(N4769), .B0(N4852), .B1(N4635));
INVXL inst_cellmath__63_0_I1055 (.Y(N4775), .A(N4645));
INVXL inst_cellmath__63_0_I1056 (.Y(N4844), .A(N4775));
INVXL inst_cellmath__63_0_I1057 (.Y(N4897), .A(N4844));
NOR2BX1 inst_cellmath__63_0_I1060 (.Y(N4798), .AN(N4844), .B(N4849));
AOI22XL inst_cellmath__63_0_I1061 (.Y(N4739), .A0(N4844), .A1(N4752), .B0(N4849), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1062 (.Y(N4778), .A0(N4844), .A1(N4828), .B0(N4752), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1063 (.Y(N4816), .A0(N4844), .A1(N4731), .B0(N4828), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1064 (.Y(N4851), .A0(N4844), .A1(N4806), .B0(N4731), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1065 (.Y(N4888), .A0(N4844), .A1(N4880), .B0(N4806), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1066 (.Y(N4753), .A0(N4844), .A1(N4783), .B0(N4880), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1067 (.Y(N4793), .A0(N4844), .A1(N4858), .B0(N4783), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1068 (.Y(N4830), .A0(N4844), .A1(N4762), .B0(N4858), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1069 (.Y(N4869), .A0(N4844), .A1(N4835), .B0(N4762), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1070 (.Y(N4733), .A0(N4844), .A1(N4740), .B0(N4835), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1071 (.Y(N4770), .A0(N4844), .A1(N4817), .B0(N4740), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1072 (.Y(N4809), .A0(N4844), .A1(N4890), .B0(N4817), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1073 (.Y(N4845), .A0(N4844), .A1(N4794), .B0(N4890), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1074 (.Y(N4883), .A0(N4844), .A1(N4870), .B0(N4794), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1075 (.Y(N4748), .A0(N4844), .A1(N4772), .B0(N4870), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1076 (.Y(N4786), .A0(N4844), .A1(N4846), .B0(N4772), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1077 (.Y(N4823), .A0(N4844), .A1(N4884), .B0(N4846), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1078 (.Y(N4861), .A0(N4844), .A1(N4749), .B0(N4884), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1079 (.Y(N4898), .A0(N4844), .A1(N4787), .B0(N4749), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1080 (.Y(N4765), .A0(N4844), .A1(N4825), .B0(N4787), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1081 (.Y(N4801), .A0(N4844), .A1(N4863), .B0(N4825), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1082 (.Y(N4837), .A0(N4844), .A1(N4728), .B0(N4863), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1083 (.Y(N4876), .A0(N4844), .A1(N4766), .B0(N4728), .B1(N4897));
AOI22XL inst_cellmath__63_0_I1084 (.Y(N4742), .A0(N4844), .A1(N4803), .B0(N4766), .B1(N4897));
INVXL inst_cellmath__63_0_I1086 (.Y(N4812), .A(N6154));
NAND2XL inst_cellmath__63_0_I1087 (.Y(N4853), .A(N4798), .B(N6154));
NAND2XL inst_cellmath__63_0_I1088 (.Y(N4755), .A(N4739), .B(N6154));
AOI22XL inst_cellmath__63_0_I1089 (.Y(N4831), .A0(N4812), .A1(N4798), .B0(N4778), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1090 (.Y(N4871), .A0(N4812), .A1(N4739), .B0(N4816), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1091 (.Y(N4734), .A0(N4812), .A1(N4778), .B0(N4851), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1092 (.Y(N4773), .A0(N4812), .A1(N4816), .B0(N4888), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1093 (.Y(N4811), .A0(N4812), .A1(N4851), .B0(N4753), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1094 (.Y(N4847), .A0(N4812), .A1(N4888), .B0(N4793), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1095 (.Y(N4885), .A0(N4812), .A1(N4753), .B0(N4830), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1096 (.Y(N4750), .A0(N4812), .A1(N4793), .B0(N4869), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1097 (.Y(N4788), .A0(N4812), .A1(N4830), .B0(N4733), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1098 (.Y(N4826), .A0(N4812), .A1(N4869), .B0(N4770), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1099 (.Y(N4864), .A0(N4812), .A1(N4733), .B0(N4809), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1100 (.Y(N4729), .A0(N4812), .A1(N4770), .B0(N4845), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1101 (.Y(N4767), .A0(N4812), .A1(N4809), .B0(N4883), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1102 (.Y(N4804), .A0(N4812), .A1(N4845), .B0(N4748), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1103 (.Y(N4840), .A0(N4812), .A1(N4883), .B0(N4786), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1104 (.Y(N4878), .A0(N4812), .A1(N4748), .B0(N4823), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1105 (.Y(N4744), .A0(N4812), .A1(N4786), .B0(N4861), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1106 (.Y(N4781), .A0(N4812), .A1(N4823), .B0(N4898), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1107 (.Y(N4820), .A0(N4812), .A1(N4861), .B0(N4765), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1108 (.Y(N4855), .A0(N4812), .A1(N4898), .B0(N4801), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1109 (.Y(N4893), .A0(N4812), .A1(N4765), .B0(N4837), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1110 (.Y(N4759), .A0(N4812), .A1(N4801), .B0(N4876), .B1(N6154));
AOI22XL inst_cellmath__63_0_I1111 (.Y(N4796), .A0(N4812), .A1(N4837), .B0(N4742), .B1(N6154));
INVXL inst_cellmath__63_0_I1113 (.Y(N4758), .A(N6161));
NOR2XL inst_cellmath__63_0_I1116 (.Y(inst_cellmath__63[2]), .A(N4758), .B(N4831));
NOR2XL inst_cellmath__63_0_I1117 (.Y(inst_cellmath__63[3]), .A(N4758), .B(N4871));
AOI22XL inst_cellmath__63_0_I1118 (.Y(inst_cellmath__63[4]), .A0(N6161), .A1(N4734), .B0(N4853), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1119 (.Y(inst_cellmath__63[5]), .A0(N6161), .A1(N4773), .B0(N4755), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1120 (.Y(inst_cellmath__63[6]), .A0(N6161), .A1(N4811), .B0(N4831), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1121 (.Y(inst_cellmath__63[7]), .A0(N6161), .A1(N4847), .B0(N4871), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1122 (.Y(inst_cellmath__63[8]), .A0(N6161), .A1(N4885), .B0(N4734), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1123 (.Y(inst_cellmath__63[9]), .A0(N6161), .A1(N4750), .B0(N4773), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1124 (.Y(inst_cellmath__63[10]), .A0(N6161), .A1(N4788), .B0(N4811), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1125 (.Y(inst_cellmath__63[11]), .A0(N6161), .A1(N4826), .B0(N4847), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1126 (.Y(inst_cellmath__63[12]), .A0(N6161), .A1(N4864), .B0(N4885), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1127 (.Y(inst_cellmath__63[13]), .A0(N6161), .A1(N4729), .B0(N4750), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1128 (.Y(inst_cellmath__63[14]), .A0(N6161), .A1(N4767), .B0(N4788), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1129 (.Y(inst_cellmath__63[15]), .A0(N6161), .A1(N4804), .B0(N4826), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1130 (.Y(inst_cellmath__63[16]), .A0(N6161), .A1(N4840), .B0(N4864), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1131 (.Y(inst_cellmath__63[17]), .A0(N6161), .A1(N4878), .B0(N4729), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1132 (.Y(inst_cellmath__63[18]), .A0(N6161), .A1(N4744), .B0(N4767), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1133 (.Y(inst_cellmath__63[19]), .A0(N6161), .A1(N4781), .B0(N4804), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1134 (.Y(inst_cellmath__63[20]), .A0(N6161), .A1(N4820), .B0(N4840), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1135 (.Y(inst_cellmath__63[21]), .A0(N6161), .A1(N4855), .B0(N4878), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1136 (.Y(inst_cellmath__63[22]), .A0(N6161), .A1(N4893), .B0(N4744), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1137 (.Y(inst_cellmath__63[23]), .A0(N6161), .A1(N4759), .B0(N4781), .B1(N4758));
AOI22XL inst_cellmath__63_0_I1138 (.Y(inst_cellmath__63[24]), .A0(N6161), .A1(N4796), .B0(N4820), .B1(N4758));
MX2XL inst_cellmath__61_0_I1139 (.Y(x[0]), .A(inst_cellmath__62), .B(inst_cellmath__63[2]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1140 (.Y(x[1]), .A(inst_cellmath__62), .B(inst_cellmath__63[3]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1141 (.Y(x[2]), .A(inst_cellmath__62), .B(inst_cellmath__63[4]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1142 (.Y(x[3]), .A(inst_cellmath__62), .B(inst_cellmath__63[5]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1143 (.Y(x[4]), .A(inst_cellmath__62), .B(inst_cellmath__63[6]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1144 (.Y(x[5]), .A(inst_cellmath__62), .B(inst_cellmath__63[7]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1145 (.Y(x[6]), .A(inst_cellmath__62), .B(inst_cellmath__63[8]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1146 (.Y(x[7]), .A(inst_cellmath__62), .B(inst_cellmath__63[9]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1147 (.Y(x[8]), .A(inst_cellmath__62), .B(inst_cellmath__63[10]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1148 (.Y(x[9]), .A(inst_cellmath__62), .B(inst_cellmath__63[11]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1149 (.Y(x[10]), .A(inst_cellmath__62), .B(inst_cellmath__63[12]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1150 (.Y(x[11]), .A(inst_cellmath__62), .B(inst_cellmath__63[13]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1151 (.Y(x[12]), .A(inst_cellmath__62), .B(inst_cellmath__63[14]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1152 (.Y(x[13]), .A(inst_cellmath__62), .B(inst_cellmath__63[15]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1153 (.Y(x[14]), .A(inst_cellmath__62), .B(inst_cellmath__63[16]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1154 (.Y(x[15]), .A(inst_cellmath__62), .B(inst_cellmath__63[17]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1155 (.Y(x[16]), .A(inst_cellmath__62), .B(inst_cellmath__63[18]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1156 (.Y(x[17]), .A(inst_cellmath__62), .B(inst_cellmath__63[19]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1157 (.Y(x[18]), .A(inst_cellmath__62), .B(inst_cellmath__63[20]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1158 (.Y(x[19]), .A(inst_cellmath__62), .B(inst_cellmath__63[21]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1159 (.Y(x[20]), .A(inst_cellmath__62), .B(inst_cellmath__63[22]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1160 (.Y(x[21]), .A(inst_cellmath__62), .B(inst_cellmath__63[23]), .S0(inst_cellmath__72));
MX2XL inst_cellmath__61_0_I1161 (.Y(x[22]), .A(inst_cellmath__62), .B(inst_cellmath__63[24]), .S0(inst_cellmath__72));
assign inst_cellmath__44[3] = 1'B0;
assign inst_cellmath__47[2] = 1'B0;
assign inst_cellmath__47[3] = 1'B0;
assign inst_cellmath__47[4] = 1'B0;
assign inst_cellmath__47[5] = 1'B0;
assign inst_cellmath__47[6] = 1'B0;
assign inst_cellmath__47[7] = 1'B0;
assign inst_cellmath__48[0] = 1'B0;
assign inst_cellmath__48[24] = 1'B1;
assign inst_cellmath__49[1] = 1'B0;
assign inst_cellmath__49[9] = 1'B0;
assign inst_cellmath__49[10] = 1'B0;
assign inst_cellmath__49[11] = 1'B0;
assign inst_cellmath__49[12] = 1'B0;
assign inst_cellmath__49[13] = 1'B0;
assign inst_cellmath__49[14] = 1'B0;
assign inst_cellmath__49[15] = 1'B0;
assign inst_cellmath__49[16] = 1'B0;
assign inst_cellmath__49[17] = 1'B0;
assign inst_cellmath__49[18] = 1'B0;
assign inst_cellmath__49[19] = 1'B0;
assign inst_cellmath__49[20] = 1'B0;
assign inst_cellmath__49[21] = 1'B0;
assign inst_cellmath__49[22] = 1'B0;
assign inst_cellmath__49[23] = 1'B0;
assign inst_cellmath__49[24] = 1'B0;
assign inst_delta[1] = 1'B0;
assign inst_cellmath__56[0] = 1'B0;
assign inst_cellmath__56[1] = 1'B0;
assign inst_cellmath__56[2] = 1'B0;
assign inst_cellmath__56[3] = 1'B0;
assign inst_cellmath__56[4] = 1'B0;
assign inst_cellmath__56[5] = 1'B0;
assign inst_cellmath__56[6] = 1'B0;
assign inst_cellmath__56[7] = 1'B0;
assign inst_cellmath__56[8] = 1'B0;
assign inst_cellmath__56[9] = 1'B0;
assign inst_cellmath__56[10] = 1'B0;
assign inst_cellmath__56[11] = 1'B0;
assign inst_cellmath__56[12] = 1'B0;
assign inst_cellmath__56[13] = 1'B0;
assign inst_cellmath__56[14] = 1'B0;
assign inst_cellmath__56[15] = 1'B0;
assign inst_cellmath__56[16] = 1'B0;
assign inst_cellmath__56[17] = 1'B0;
assign inst_cellmath__56[18] = 1'B0;
assign inst_cellmath__56[19] = 1'B0;
assign inst_cellmath__56[20] = 1'B0;
assign inst_cellmath__56[21] = 1'B0;
assign inst_cellmath__56[22] = 1'B0;
assign inst_cellmath__56[23] = 1'B0;
assign inst_cellmath__56[24] = 1'B0;
assign inst_cellmath__63[0] = 1'B0;
assign inst_cellmath__63[1] = 1'B0;
endmodule

/* CADENCE  s7jzTwrYqw== : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



