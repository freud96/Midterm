/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:23:56 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42;
wire [22:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68;
wire [0:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195;
wire [20:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197;
wire [32:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N623,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5570,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5577,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5578,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5600,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5607,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5614,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5616,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5623,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5629,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5641,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5657,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5664,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5754,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5866,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5869,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6087,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6179,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6189,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6197,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6224,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6256,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6257,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6258,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6292,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6299,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6310,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6347,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6356,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6359,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6381,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6396,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7360,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7365,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7438,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7450,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7555,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7570,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7929,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8158,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8179,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8197,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8221,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8222,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8252,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8292,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8294,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8360,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8361,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8364,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8382,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8384,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8405,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8425,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8429,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8436,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8442,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8445,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8452,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8459,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8465,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8471,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8474,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8485,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8502,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8537,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8539,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8555,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8579,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8586,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8607,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8612,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8614,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8616,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8632,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8657,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8735,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8860,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8868,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8900,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9059,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9087,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9093,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10425,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10430,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10436,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10438,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10442,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10443,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10445,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10449,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10450,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10452,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10459,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10465,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10470,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10475,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10476,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10500,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10558,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10593,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10600,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10613,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10617,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10629,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10661,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10765,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10797,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10807,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10860,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10861,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10889,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11735,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11738,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11760,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11765,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11791,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11806,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11807,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11826,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11830,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11863,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11866,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11869,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11904,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11931,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12047,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12059,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12087,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12093,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12118,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12129,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12145,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12165,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12189,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12193,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12194,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12221,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12224,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12229,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12240,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12256,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12269,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12347,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12356,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12361,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12364,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12365,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12367,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12381,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12384,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12396,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12406,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12429,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12431,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12438,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12447,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12470,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12474,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12475,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12476,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12490,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12491,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12501,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12502,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12520,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12527,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12532,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12537,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12567,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12578,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12579,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12593,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12599,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12602,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12607,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12613,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12614,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12617,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12629,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12632,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12642,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12654,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12661,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12664,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12714,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12738,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12765,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12791,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12797,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12826,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12830,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12850,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12860,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12861,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12863,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12868,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12889,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12900,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13047,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13093,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13129,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13149,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13158,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13165,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13168,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13177,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13189,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13197,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13222,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13224,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13228,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13229,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13252,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13253,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13258,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13299,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13310,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15129,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15177,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15257,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15429,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15466,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15485,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15490,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15539,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16294,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16500,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16537,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16542,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16662,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16754,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17256,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23240,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23367,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45118,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45252,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45341,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45612,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45854;
wire N20585,N20596,N20746,N20748,N21279,N21282,N21470 
	,N21688,N22491,N22530,N22533,N22538,N22540,N22545,N22547 
	,N22552,N22554,N22559,N22561,N22566,N22575,N22580,N22583 
	,N22585,N22594,N22597,N22599,N22606,N22611,N22616,N22621 
	,N22624,N22626,N22636,N22641,N22648,N22651,N22672,N22682 
	,N22708,N22728,N22764,N22772,N22791,N22793,N22798,N22800 
	,N22812,N22814,N22816,N22826,N22828,N22830,N22833,N22835 
	,N22837,N22841,N22843,N22845,N22848,N22850,N22852,N22858 
	,N22860,N22864,N22866,N22868,N22871,N22873,N22875,N22881 
	,N22883,N22889,N22891,N22895,N22897,N22899,N22903,N22905 
	,N22907,N22910,N22919,N22973,N22978,N22985,N22992,N23039 
	,N23041,N23043,N23049,N23051,N23099,N23101,N23103,N23137 
	,N23601,N23606,N23608,N23613,N23615,N23620,N23628,N23630 
	,N23638,N23640,N23646,N23917,N23918,N23919,N23920,N23921 
	,N23922,N23923,N23924,N23925,N23926,N23927,N23928,N23929 
	;
reg x_reg_20__retimed_I14257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14257_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15184;
	end
assign N23646 = x_reg_20__retimed_I14257_QOUT;
reg x_reg_23__retimed_I14255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I14255_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547;
	end
assign N23640 = x_reg_23__retimed_I14255_QOUT;
reg x_reg_23__retimed_I14254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I14254_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15399;
	end
assign N23638 = x_reg_23__retimed_I14254_QOUT;
reg x_reg_20__retimed_I14251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14251_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999;
	end
assign N23630 = x_reg_20__retimed_I14251_QOUT;
reg x_reg_20__retimed_I14250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14250_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973;
	end
assign N23628 = x_reg_20__retimed_I14250_QOUT;
reg x_reg_20__retimed_I14247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14247_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15019;
	end
assign N23620 = x_reg_20__retimed_I14247_QOUT;
reg x_reg_20__retimed_I14245_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14245_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967;
	end
assign N23615 = x_reg_20__retimed_I14245_QOUT;
reg x_reg_20__retimed_I14244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14244_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15487;
	end
assign N23613 = x_reg_20__retimed_I14244_QOUT;
reg x_reg_20__retimed_I14242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14242_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253;
	end
assign N23608 = x_reg_20__retimed_I14242_QOUT;
reg x_reg_20__retimed_I14241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14241_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15113;
	end
assign N23606 = x_reg_20__retimed_I14241_QOUT;
reg x_reg_20__retimed_I14239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14239_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15386;
	end
assign N23601 = x_reg_20__retimed_I14239_QOUT;
reg x_reg_20__retimed_I14063_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14063_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15008;
	end
assign N23137 = x_reg_20__retimed_I14063_QOUT;
reg x_reg_20__retimed_I14046_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14046_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15490;
	end
assign N23103 = x_reg_20__retimed_I14046_QOUT;
reg x_reg_20__retimed_I14045_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14045_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464;
	end
assign N23101 = x_reg_20__retimed_I14045_QOUT;
reg x_reg_20__retimed_I14044_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14044_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320;
	end
assign N23099 = x_reg_20__retimed_I14044_QOUT;
reg x_reg_20__retimed_I14026_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14026_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15428;
	end
assign N23051 = x_reg_20__retimed_I14026_QOUT;
reg x_reg_20__retimed_I14025_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14025_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15283;
	end
assign N23049 = x_reg_20__retimed_I14025_QOUT;
reg x_reg_20__retimed_I14023_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14023_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232;
	end
assign N23043 = x_reg_20__retimed_I14023_QOUT;
reg x_reg_20__retimed_I14022_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14022_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208;
	end
assign N23041 = x_reg_20__retimed_I14022_QOUT;
reg x_reg_20__retimed_I14021_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14021_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069;
	end
assign N23039 = x_reg_20__retimed_I14021_QOUT;
reg x_reg_20__retimed_I14003_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14003_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597;
	end
assign N22992 = x_reg_20__retimed_I14003_QOUT;
reg x_reg_20__retimed_I14000_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I14000_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15105;
	end
assign N22985 = x_reg_20__retimed_I14000_QOUT;
reg x_reg_20__retimed_I13997_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13997_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219;
	end
assign N22978 = x_reg_20__retimed_I13997_QOUT;
reg x_reg_20__retimed_I13995_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13995_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15071;
	end
assign N22973 = x_reg_20__retimed_I13995_QOUT;
reg x_reg_20__retimed_I13973_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13973_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15448;
	end
assign N22919 = x_reg_20__retimed_I13973_QOUT;
reg x_reg_20__retimed_I13969_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13969_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15473;
	end
assign N22910 = x_reg_20__retimed_I13969_QOUT;
reg x_reg_20__retimed_I13968_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13968_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378;
	end
assign N22907 = x_reg_20__retimed_I13968_QOUT;
reg x_reg_20__retimed_I13967_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13967_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15524;
	end
assign N22905 = x_reg_20__retimed_I13967_QOUT;
reg x_reg_20__retimed_I13966_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13966_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15376;
	end
assign N22903 = x_reg_20__retimed_I13966_QOUT;
reg x_reg_20__retimed_I13965_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13965_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15352;
	end
assign N22899 = x_reg_20__retimed_I13965_QOUT;
reg x_reg_20__retimed_I13964_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13964_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15550;
	end
assign N22897 = x_reg_20__retimed_I13964_QOUT;
reg x_reg_20__retimed_I13963_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13963_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15207;
	end
assign N22895 = x_reg_20__retimed_I13963_QOUT;
reg x_reg_20__retimed_I13962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13962_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154;
	end
assign N22891 = x_reg_20__retimed_I13962_QOUT;
reg x_reg_20__retimed_I13961_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13961_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15064;
	end
assign N22889 = x_reg_20__retimed_I13961_QOUT;
reg x_reg_20__retimed_I13959_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13959_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15152;
	end
assign N22883 = x_reg_20__retimed_I13959_QOUT;
reg x_reg_20__retimed_I13958_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13958_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530;
	end
assign N22881 = x_reg_20__retimed_I13958_QOUT;
reg x_reg_20__retimed_I13956_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13956_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15044;
	end
assign N22875 = x_reg_20__retimed_I13956_QOUT;
reg x_reg_20__retimed_I13955_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13955_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513;
	end
assign N22873 = x_reg_20__retimed_I13955_QOUT;
reg x_reg_20__retimed_I13954_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13954_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361;
	end
assign N22871 = x_reg_20__retimed_I13954_QOUT;
reg x_reg_20__retimed_I13953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13953_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15463;
	end
assign N22868 = x_reg_20__retimed_I13953_QOUT;
reg x_reg_20__retimed_I13952_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13952_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15265;
	end
assign N22866 = x_reg_20__retimed_I13952_QOUT;
reg x_reg_20__retimed_I13951_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13951_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15127;
	end
assign N22864 = x_reg_20__retimed_I13951_QOUT;
reg x_reg_20__retimed_I13950_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13950_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15175;
	end
assign N22860 = x_reg_20__retimed_I13950_QOUT;
reg x_reg_20__retimed_I13949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13949_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14981;
	end
assign N22858 = x_reg_20__retimed_I13949_QOUT;
reg x_reg_20__retimed_I13947_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13947_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15539;
	end
assign N22852 = x_reg_20__retimed_I13947_QOUT;
reg x_reg_20__retimed_I13946_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13946_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15338;
	end
assign N22850 = x_reg_20__retimed_I13946_QOUT;
reg x_reg_20__retimed_I13945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13945_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15195;
	end
assign N22848 = x_reg_20__retimed_I13945_QOUT;
reg x_reg_20__retimed_I13944_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13944_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15435;
	end
assign N22845 = x_reg_20__retimed_I13944_QOUT;
reg x_reg_20__retimed_I13943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13943_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012;
	end
assign N22843 = x_reg_20__retimed_I13943_QOUT;
reg x_reg_20__retimed_I13942_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13942_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15290;
	end
assign N22841 = x_reg_20__retimed_I13942_QOUT;
reg x_reg_20__retimed_I13941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13941_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15241;
	end
assign N22837 = x_reg_20__retimed_I13941_QOUT;
reg x_reg_20__retimed_I13940_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13940_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15054;
	end
assign N22835 = x_reg_20__retimed_I13940_QOUT;
reg x_reg_20__retimed_I13939_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13939_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15573;
	end
assign N22833 = x_reg_20__retimed_I13939_QOUT;
reg x_reg_20__retimed_I13938_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13938_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15499;
	end
assign N22830 = x_reg_20__retimed_I13938_QOUT;
reg x_reg_20__retimed_I13937_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13937_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306;
	end
assign N22828 = x_reg_20__retimed_I13937_QOUT;
reg x_reg_20__retimed_I13936_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13936_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15161;
	end
assign N22826 = x_reg_20__retimed_I13936_QOUT;
reg x_reg_20__retimed_I13932_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13932_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14956;
	end
assign N22816 = x_reg_20__retimed_I13932_QOUT;
reg x_reg_20__retimed_I13931_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13931_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15420;
	end
assign N22814 = x_reg_20__retimed_I13931_QOUT;
reg x_reg_20__retimed_I13930_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13930_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15278;
	end
assign N22812 = x_reg_20__retimed_I13930_QOUT;
reg x_reg_20__retimed_I13925_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13925_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15135;
	end
assign N22800 = x_reg_20__retimed_I13925_QOUT;
reg x_reg_20__retimed_I13924_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13924_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14992;
	end
assign N22798 = x_reg_20__retimed_I13924_QOUT;
reg x_reg_20__retimed_I13922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13922_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15565;
	end
assign N22793 = x_reg_20__retimed_I13922_QOUT;
reg x_reg_20__retimed_I13921_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13921_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15409;
	end
assign N22791 = x_reg_20__retimed_I13921_QOUT;
reg x_reg_20__retimed_I13914_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13914_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15297;
	end
assign N22772 = x_reg_20__retimed_I13914_QOUT;
reg x_reg_20__retimed_I13911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13911_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15589;
	end
assign N22764 = x_reg_20__retimed_I13911_QOUT;
reg x_reg_20__retimed_I13906_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13906_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15123;
	end
assign N22728 = x_reg_20__retimed_I13906_QOUT;
reg x_reg_20__retimed_I13898_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13898_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15441;
	end
assign N22708 = x_reg_20__retimed_I13898_QOUT;
reg x_reg_20__retimed_I13887_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13887_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15518;
	end
assign N22682 = x_reg_20__retimed_I13887_QOUT;
reg x_reg_20__retimed_I13883_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13883_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15226;
	end
assign N22672 = x_reg_20__retimed_I13883_QOUT;
reg x_reg_20__retimed_I13874_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13874_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15372;
	end
assign N22651 = x_reg_20__retimed_I13874_QOUT;
reg x_reg_20__retimed_I13873_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13873_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14966;
	end
assign N22648 = x_reg_20__retimed_I13873_QOUT;
reg x_reg_20__retimed_I13870_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13870_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15559;
	end
assign N22641 = x_reg_20__retimed_I13870_QOUT;
reg x_reg_20__retimed_I13868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13868_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15100;
	end
assign N22636 = x_reg_20__retimed_I13868_QOUT;
reg x_reg_20__retimed_I13864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13864_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050;
	end
assign N22626 = x_reg_20__retimed_I13864_QOUT;
reg x_reg_20__retimed_I13863_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13863_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45835;
	end
assign N22624 = x_reg_20__retimed_I13863_QOUT;
reg x_reg_20__retimed_I13862_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13862_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15397;
	end
assign N22621 = x_reg_20__retimed_I13862_QOUT;
reg x_reg_20__retimed_I13860_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13860_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14991;
	end
assign N22616 = x_reg_20__retimed_I13860_QOUT;
reg x_reg_20__retimed_I13858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13858_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14944;
	end
assign N22611 = x_reg_20__retimed_I13858_QOUT;
reg x_reg_20__retimed_I13856_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13856_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15170;
	end
assign N22606 = x_reg_20__retimed_I13856_QOUT;
reg x_reg_20__retimed_I13853_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13853_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301;
	end
assign N22599 = x_reg_20__retimed_I13853_QOUT;
reg x_reg_20__retimed_I13852_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13852_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45811;
	end
assign N22597 = x_reg_20__retimed_I13852_QOUT;
reg x_reg_20__retimed_I13851_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13851_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15534;
	end
assign N22594 = x_reg_20__retimed_I13851_QOUT;
reg x_reg_20__retimed_I13847_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13847_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273;
	end
assign N22585 = x_reg_20__retimed_I13847_QOUT;
reg x_reg_20__retimed_I13846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13846_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45829;
	end
assign N22583 = x_reg_20__retimed_I13846_QOUT;
reg x_reg_20__retimed_I13845_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13845_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15192;
	end
assign N22580 = x_reg_20__retimed_I13845_QOUT;
reg x_reg_20__retimed_I13843_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13843_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15147;
	end
assign N22575 = x_reg_20__retimed_I13843_QOUT;
reg x_reg_20__retimed_I13839_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13839_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15325;
	end
assign N22566 = x_reg_20__retimed_I13839_QOUT;
reg x_reg_20__retimed_I13837_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13837_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247;
	end
assign N22561 = x_reg_20__retimed_I13837_QOUT;
reg x_reg_20__retimed_I13836_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13836_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45847;
	end
assign N22559 = x_reg_20__retimed_I13836_QOUT;
reg x_reg_20__retimed_I13834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13834_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481;
	end
assign N22554 = x_reg_20__retimed_I13834_QOUT;
reg x_reg_20__retimed_I13833_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13833_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45841;
	end
assign N22552 = x_reg_20__retimed_I13833_QOUT;
reg x_reg_20__retimed_I13831_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13831_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075;
	end
assign N22547 = x_reg_20__retimed_I13831_QOUT;
reg x_reg_20__retimed_I13830_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13830_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45817;
	end
assign N22545 = x_reg_20__retimed_I13830_QOUT;
reg x_reg_20__retimed_I13828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13828_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508;
	end
assign N22540 = x_reg_20__retimed_I13828_QOUT;
reg x_reg_20__retimed_I13827_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13827_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45823;
	end
assign N22538 = x_reg_20__retimed_I13827_QOUT;
reg x_reg_20__retimed_I13825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13825_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15583;
	end
assign N22533 = x_reg_20__retimed_I13825_QOUT;
reg x_reg_20__retimed_I13824_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13824_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15348;
	end
assign N22530 = x_reg_20__retimed_I13824_QOUT;
reg x_reg_20__retimed_I13812_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I13812_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15419;
	end
assign N22491 = x_reg_20__retimed_I13812_QOUT;
reg x_reg_23__retimed_I13554_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I13554_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15081;
	end
assign N21688 = x_reg_23__retimed_I13554_QOUT;
reg x_reg_23__retimed_I13476_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I13476_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15143;
	end
assign N21470 = x_reg_23__retimed_I13476_QOUT;
reg x_reg_23__retimed_I13410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I13410_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22];
	end
assign N21282 = x_reg_23__retimed_I13410_QOUT;
reg x_reg_23__retimed_I13409_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I13409_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455;
	end
assign N21279 = x_reg_23__retimed_I13409_QOUT;
reg x_reg_27__retimed_I13216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__retimed_I13216_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178;
	end
assign N20748 = x_reg_27__retimed_I13216_QOUT;
reg x_reg_27__retimed_I13215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__retimed_I13215_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594;
	end
assign N20746 = x_reg_27__retimed_I13215_QOUT;
reg x_reg_21__retimed_I13151_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I13151_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741;
	end
assign N20596 = x_reg_21__retimed_I13151_QOUT;
assign N23917 = !N20596;
assign N23922 = !N23917;
assign N23921 = !N23917;
assign N23920 = !N23917;
assign N23919 = !N23917;
assign N23918 = !N23917;
reg x_reg_22__retimed_I13146_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I13146_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163;
	end
assign N20585 = x_reg_22__retimed_I13146_QOUT;
assign N23923 = !N20585;
assign N23924 = !N23923;
assign bdw_enable = !astall;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45150 = !(a_exp[6] & a_exp[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16362 = !(a_exp[4] & a_exp[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328 = !(a_exp[2] & a_exp[1]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16357 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16362 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45152 = !((a_exp[7] & a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16357);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45150 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45152);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16464 = !(a_sign & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122 = !a_man[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16403 = !(a_man[0] | a_man[1]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16417 = !(a_man[12] | a_man[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16386 = !(a_man[18] | a_man[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16397 = !(a_man[16] | a_man[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16407 = !(a_man[14] | a_man[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16409 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16417 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16386) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16397) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16407;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23456 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16403) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16409);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213 = !(a_man[22] | a_man[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16411 = !(a_man[4] | a_man[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16380 = !(a_man[10] | a_man[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16390 = !(a_man[8] | a_man[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16401 = !(a_man[6] | a_man[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16393 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16411 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16380) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16390) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16401;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16376 = !(a_man[20] | a_man[19]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23456) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16393) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16376);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16464 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19) | a_sign) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268 = !a_exp[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289 = !a_exp[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264 = !a_exp[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7281 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287 = !a_exp[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280 = !a_exp[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293 = !a_exp[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7281 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267 = !a_exp[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[7] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7270 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7271 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7270);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[6] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7271 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[7] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45146 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16334 = !(a_exp[3] | a_exp[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16332 = !(a_exp[5] & a_exp[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16324 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16334 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16332);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16294 = ((a_exp[7] | a_exp[6]) | a_exp[0]) | a_exp[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16298 = ((a_exp[4] | a_exp[2]) | a_exp[3]) | a_exp[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16324 | a_exp[7]) & (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16294 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16298);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45132 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45119 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45118 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45119);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45146 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45132) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45118;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[29] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974 = !(a_exp[4] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45763 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45763;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406 = !(a_man[22] & a_man[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354 = !a_man[21];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341} = {1'B0, a_man[20]} + {1'B0, a_man[22]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965} = {1'B0, a_man[19]} + {1'B0, a_man[21]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6172 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5610 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6172;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6283 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6212, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6017} = {1'B0, a_man[17]} + {1'B0, a_man[19]} + {1'B0, a_man[22]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594} = {1'B0, a_man[18]} + {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6212};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201 = !a_man[16];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5833, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5644} = {1'B0, a_man[18]} + {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078} = {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5833} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6017};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6154 = a_man[15] | a_man[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870 = !a_man[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6261 = a_man[14] | a_man[16];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6317, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6131} = {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6261};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6154} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5644} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6317};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6377 = a_man[13] | a_man[15];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5940, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5749} = {1'B0, a_man[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6377};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5962 = (!a_man[15]) ^ a_man[17];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5962} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5940} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6131};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981 = !a_man[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5621 = a_man[12] | a_man[14];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5572, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6241} = {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5621};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6077 = (!a_man[14]) ^ a_man[16];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6077} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5572} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5749};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6108, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5915} = {1'B0, a_man[11]} + {1'B0, a_man[13]} + {1'B0, a_man[16]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605 = !a_man[19];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6051, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5866} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6108} + {1'B0, a_man[17]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6190 = (!a_man[13]) ^ a_man[15];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6051} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6241};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089 = !a_man[18];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6218, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6025} = {1'B0, a_man[10]} + {1'B0, a_man[12]} + {1'B0, a_man[15]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705 = !a_man[17];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5721, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6413} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5671, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6348} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6218} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5721};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6292 = (!a_man[12]) ^ a_man[14];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6292} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5671} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5866};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6326, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6141} = {1'B0, a_man[9]} + {1'B0, a_man[11]} + {1'B0, a_man[14]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6166, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5973} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6326} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6025} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6413};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5915} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6348} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6166};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6115 = a_man[22] | a_man[8];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5840, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5651} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6115} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821 = !a_man[15];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5581, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6248} = {1'B0, a_man[10]} + {1'B0, a_man[13]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5732, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6421} = {1'B0, a_man[21]} + {1'B0, a_man[7]} + {1'B0, a_man[9]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5922 = (!a_man[22]) ^ a_man[8];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5949, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5759} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5732} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5922};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5787, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5600} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5581} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6141} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5949};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5840} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5973} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5787};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308 = !a_man[14];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5680, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6357} = {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5849, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5656} = {1'B0, a_man[20]} + {1'B0, a_man[6]} + {1'B0, a_man[8]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929 = !a_man[13];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6223, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6034} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929} + {1'B0, a_man[11]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6060, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5876} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6223} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5849} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6421};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6274, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6085} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5680} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6248} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6060};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5651} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6274} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5600};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565 = !a_man[12];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6336, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6148} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5793, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5609} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6336};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5956, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5769} = {1'B0, a_man[19]} + {1'B0, a_man[5]} + {1'B0, a_man[7]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6174, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5983} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5956} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6034} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5656};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5895, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5700} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6357} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5793} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6174};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5759} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5895} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6085};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041 = !a_man[11];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5589, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6255} = {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5903, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5708} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5589};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6070, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5883} = {1'B0, a_man[18]} + {1'B0, a_man[4]} + {1'B0, a_man[6]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6281, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6092} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6148} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6070} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5769};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6388, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6197} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5609} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5903} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6281};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5876} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6388} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5700};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662 = !a_man[10];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5686, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6370} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662} + {1'B0, a_man[8]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6009, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5824} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5686} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6289, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6101} = {1'B0, a_man[16]} + {1'B0, a_man[2]} + {1'B0, a_man[4]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6123, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5933} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6289};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155 = !a_man[9];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5803, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5616} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308} + {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6182, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5988} = {1'B0, a_man[17]} + {1'B0, a_man[3]} + {1'B0, a_man[5]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5635, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6310} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6370} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5803} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5988};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5627, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6303} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6123} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5824} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5635};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6396, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6204} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6255} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6182} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5883};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6004, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5817} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6009} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5708} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6396};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6092} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5627} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5817};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5983} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6004} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6197};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6133, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5942} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6243, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6054} = {1'B0, a_man[21]} + {1'B0, a_man[14]} + {1'B0, a_man[0]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263 = !a_man[7];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5752, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5574} = {1'B0, a_man[2]} + {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6343, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6157} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6243} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6133} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5752};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5646 = a_man[22] | a_man[15];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6407, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6214} = {1'B0, a_man[1]} + {1'B0, a_man[3]} + {1'B0, a_man[6]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6233, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6045} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5646} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6407};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6318 = (!a_man[22]) ^ a_man[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778 = !a_man[8];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5910, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5717} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5857, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5664} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6214} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6318} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5717};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5734, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5560} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6045} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6343} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5857};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5742, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5566} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6101} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5910} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5616};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6117, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5923} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6233} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5933} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5742};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5734} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6310} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5923};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6204} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6117} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6303};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5601 = a_man[20] | a_man[13];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5867, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5674} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927 = !a_man[6];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6351, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6167} = {1'B0, a_man[1]} + {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5595, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6267} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5867} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5601} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6351};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5966, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5780} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5942} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6054} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5574};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6224, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6036} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6157} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5595} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5966};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5566} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6224} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5560};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6087, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5896} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5819 = a_man[19] | a_man[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378 = !a_man[5];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5702, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6391} = {1'B0, a_man[0]} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5695, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6381} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5819} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6087} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5702};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6276 = (!a_man[20]) ^ a_man[13];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6079, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5891} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5674} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6276} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6167};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5852, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5659} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5695} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6267} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6079};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5664} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5852} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6036};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5925, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5736} = {1'B0, a_man[18]} + {1'B0, a_man[11]} + {1'B0, a_man[2]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995 = !a_man[4];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6305, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6120} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5810, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5623} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5925} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6305};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6152 = a_man[17] | a_man[10];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5562, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6225} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5918, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5727} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6152} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5562};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716 = !a_man[3];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6038, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5854} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6297, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6110} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6120} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6038} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5736};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5958, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5774} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5918} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5623} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6297};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5629 = (!a_man[19]) ^ a_man[12];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6192, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5998} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5629} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5896} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6391};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6337, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6150} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6192} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5810} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6381};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5891} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5958} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6150};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5780} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6337} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5659};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6389 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723 = !a_man[1];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5894, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5699} = {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5786, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5598} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5754, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5575} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5598} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5894} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5669, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6347} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6272, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6084} = {1'B0, a_man[7]} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6163, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5971} = {1'B0, a_man[8]} + {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6134, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5945} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5786} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6272} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5971};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6347} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5754} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5945};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5980 = (!a_man[9]) ^ a_man[2];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5570, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6237} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5980};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740 = !a_man[0];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6050, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5862} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5648, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6320} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6163} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5669} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5862};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6134} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6237} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6320};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6171 = a_man[9] | a_man[2];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6056, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5872} = {1'B0, a_man[10]} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6314, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6127} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6171} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5872};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5937, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5748} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6021, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5837} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6050} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5748} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5570};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5837} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6127} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5648};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5848 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5578, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6246} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122} + {1'B0, a_man[4]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6207, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6013} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6056} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6246};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5828, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5640} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6409, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6215} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5937} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5640} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6314};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6013} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6021} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6215};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5947, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5755} = {1'B0, a_man[12]} + {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6096, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5906} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5578} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5755};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5713, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6399} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5911, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5718} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6399} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5828} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6207};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6409} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5906} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5718};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5577 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5577);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5848 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5869, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5675} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6002 = a_man[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6244, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6055} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6002} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5869} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5699} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6055};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6084} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6244} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5575};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6181 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5815 = (!a_man[5]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6352, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6169} = {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6352} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5815} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5675};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6279 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5976, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5789} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5604, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6278} = {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5604} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5789} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5976} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6169} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5703, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6392} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6088, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5899} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5899} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5703} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6088} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6278} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6315 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6200, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6007} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6392} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6200} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5820, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5631} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5820} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6007};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6173 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5563 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5634 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6309 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6339 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6188 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5634) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6309);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5823 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6203 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6227 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5823 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6203);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5898 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6339) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5563)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6227);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5739 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5739} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5901 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5706 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5944 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5901 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5898) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5706);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5631};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6020 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6091 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5607 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5835 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6091) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5607);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5771 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6020) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5944)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5835);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5982 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6356 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5856 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5982 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6356;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6239 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6173) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5771) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5856);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5875 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6247 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6130 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5875 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6247);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5758 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6138 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6015 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5758 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6138);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6137 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6130) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6015));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5704 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6315 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6239) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6090 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6100 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5704 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6279) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6090);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5606 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5979 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5989 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5606 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5979);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6100) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6181)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5989);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6355 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5871 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5658 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6355 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5871);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6245 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5757 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6420 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6245) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5757);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5658) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6420);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5776, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45273} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6374 = a_man[16] | a_man[9];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6259, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45245} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6030, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5843} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6374} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5776} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6259};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5960 = (!a_man[17]) ^ a_man[10];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6416, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6220} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6225} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5960} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5854};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5591, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6256} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6030} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5727} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6416};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5591} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5998} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5774};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6105 = a_man[15] | a_man[8];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45282, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45267} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6144, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45276} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6105} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45282};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45296 = (!a_man[16]) ^ a_man[9];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5653, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45239} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45273} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45296} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45245};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6072, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5885} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6144} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5843} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5653};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6110} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6072} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6256};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5839 = a_man[14] | a_man[7];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45300, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45286} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5839};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45242, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45293} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6322, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6136} = {1'B0, a_man[13]} + {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5650 = (!a_man[14]) ^ a_man[7];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45238, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45290} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45270, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5683} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5650} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6322} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45290};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45246, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45297} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45242} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45286} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45270};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45254 = (!a_man[15]) ^ a_man[8];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45262, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45249} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45238} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45254} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45267};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5687, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45259} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45276} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45300} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45262};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45239} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45246} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45259};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6220} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5687} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5885};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45252, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6285} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45279, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5799} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5947} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6136};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45283, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5618} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45252} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45293} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45279};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45249} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45283} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45297};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6290, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6103} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5713} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6285} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6096};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6290} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5683} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5618};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5799} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5911} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6103};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6135 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5649 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6135) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5649);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5970 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5970);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6401 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6401);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5952 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5952);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6380 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6380);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5932 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5932);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6359 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6359);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5914 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5691 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5914);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5641 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5691;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5773 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5641);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6196 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5773);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6389) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6196);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6283) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5610));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5681 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5619 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6358 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5619 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5681)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6358));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5657 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5657);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5890 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5890;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6003 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6258 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5816 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6258);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6003) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5816);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6415 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5934 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6415;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5744 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5744) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5934));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5770 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6189 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5770);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6189);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6230 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6230;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7528 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N706 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7528);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44981 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652 & a_exp[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071 = !a_exp[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45019 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45064 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45045 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45064) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45019));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45070 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45045);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45016 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45043 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45065 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45043) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45016));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45031 = !(a_exp[0] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45065);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45015 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45070) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45031);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45040 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45050 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45040 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45068 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45033 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45068 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45052 = !((a_exp[0] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45050) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45033);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45023 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45072 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45023 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45020 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45036 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45020 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45072) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45055 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45052) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45036);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45015 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45055);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44981 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N706 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7428 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45464 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45473 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45473) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45464));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45454 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45454));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6022 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6022 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5711 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5666 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5711;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6345 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6345) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5666));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6235 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5968 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6235;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5784 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5784) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5968));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6299 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6112 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5628 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6302 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5628) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6302);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6299));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6277 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6277) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5576 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5576 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6300 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45446 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6300;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45439 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45439) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5955 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45460 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5955;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45451 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45451) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45460));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7478 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7478));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6063 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6234 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6063;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6048 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6048) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6234));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7365 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7365) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7423 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7348 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7423) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7428));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N697 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7348);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N697 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7570 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5977 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5977 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6018 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5729 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6018;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6418 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6116 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6208 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5924 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6208 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6116) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5924);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6418) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5729));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7366 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7549 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N696 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7549);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N696 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12808 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7477 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7404 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7477);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N698 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7404);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N698;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12808 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11882 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11882 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7416 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N705 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7416);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N705 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7559 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N704 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7559);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N704 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7450 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N703 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7450);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N703 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7480 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N701 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7480);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N701 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7337 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N702 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7337);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N702 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8780 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8780;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8161 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8161;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9127 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9127;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8407 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8605 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8407);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9026 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9026;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8940 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7961 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9059 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8940 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7961);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8345 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9059);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8345 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8605;
assign N23925 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084;
assign N23926 = !N23925;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475 = !((a_exp[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543) | ((!a_exp[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7535 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7513 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7535);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N699 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7513);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N699 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12781 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7370 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N700 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7370);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[16] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N700 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12781 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11849 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11849 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8478 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8670 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8106 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8670);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8920 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8223 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8106 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8920);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8743 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8478 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8223);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8624 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8624 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8743;
assign N23927 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707;
assign N23928 = !N23927;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12225 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[41], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[40]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12225};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8405 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8210 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8405 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8040 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8192 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8252 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8192);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8909 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8252 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7934 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8909 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8024 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8151 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8465 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8151) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8728 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8024 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8465);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[22] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8210 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8040) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7934) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8728);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8652 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7968 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8774 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8652 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7968);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8898 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8774);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8349 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9067 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8080 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9067 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N761 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8080 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8349) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8898));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N761;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11854 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12363 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12261 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7460 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5672 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6032 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5672;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5846 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6032));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7566 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45504 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7566) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7460));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45494 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45504);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45494 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45771 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45771;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7349 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6333 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6146 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6146) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6333));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7510 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7438 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7510) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N694 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7438);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[10] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N694 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12835 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12835 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8678 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8749 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8678 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8597 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8749 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8058 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8635 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8484 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8635);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8325 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8058 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8484);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8597 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8325;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13146 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12916, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12581} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12261} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13146};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[40], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[39]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12363} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11854} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12916};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[22]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[40]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[40]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9111 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8919 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9053 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9111 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8936 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8584 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8992 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8584);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8821 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8759 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8936 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8992) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8821;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[21] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9053 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8759);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11913 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11913 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12658 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7492 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5737 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5737) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7456 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7379 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7456) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7492));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7379);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7833 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7833));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6394 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6394);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5733 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5766 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5733;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5587 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5587) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5766));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7400 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7324 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7400) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N692 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7324);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N692 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12863 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12863 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11894 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12422, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12066} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12658} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11894};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13186 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12298 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13297 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12127, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11750} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12298} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13186} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13297};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8186 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8657 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8186 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8783 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9010 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8950 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9010);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8444 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7977 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8444);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9076 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8950 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7977);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8905 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8783 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9076);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8085 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8248 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8353 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8085 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8248);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8905 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8353;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12785 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13130, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12772} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12785} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12127} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12066};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[39], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[38]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12422} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12581} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13130};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[39]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[39]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8502 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8074 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9142 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8502 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8074);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8138 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8767 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8844 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8138) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8767;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8158 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8844);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8454 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8411 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8454;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[20] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9142) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8158) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8411);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11947 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11947 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12692 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6257 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6068 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6257;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5881 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6068));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7387 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7343 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7387));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7524 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7343) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7524);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7809 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7809));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6368 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6179 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6179) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6368));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7331 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7544 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7331));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7469 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7544) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N690 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7469);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[6] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N690;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12892 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12892 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8579 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7984 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8857 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7984 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7895 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8000 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8857 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7895);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8638 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8579) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8000);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8519 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8169 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8519);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8425 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8123 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8169 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8425);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8618 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8273 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8618);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8537 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8273 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8377 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8123 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8537);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8377;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7918 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8448 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8026 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8448);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8338 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8711 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8338);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8562 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7918 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8026) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8711) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8562;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12078 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11813, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13105} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12692} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12078};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12439 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11905, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13196} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12439} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11813} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11750};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12816 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11931 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8798 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9089 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8471 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8798 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9089);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8259 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8522 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8739 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8259 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8522);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8317 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8471 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8739);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8173 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8317) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8846 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8101 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8846 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7989 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8218 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7989 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8586 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8101 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8218);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7937 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8432 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8586 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7937);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8432 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8173;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11703 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12331 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11688 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11721, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13010} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12331} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11703} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11688};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12551, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12186} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11931} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12816} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11721};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12477 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13222 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11978 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11978 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12721 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6075 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6075) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7531 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7487 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7531));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7412 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7487) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N689 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7412);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N689 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45756 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6393 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6393 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5801 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45756) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5614 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5614) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5801));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7473 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7434 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7473));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7355 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7434) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N688 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7355);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N688;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12926 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12926 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12115 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13304, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12923} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12721} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12115};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13168, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12800} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13222} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12477} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13304};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13265, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12888} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13105} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13168} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12186};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12635, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12275} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12551} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13196} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13265};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[38], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[37]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11905} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12772} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12635};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[38]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[38]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8625 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8671 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8528 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8571 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8921 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8528 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8571);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8744 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8921);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8867 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8671 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8744);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8053 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8107 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7903 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8053 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8107);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8590 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[19] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8625 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8867) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7903) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10403 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10442 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10576 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10442} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10403} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10576};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10425 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10457 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10493 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10855 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10920 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10666, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10529} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10855} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10493} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10920};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10457} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10425} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10666};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10778 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10992 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10592 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10737, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10610} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10992} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10592};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10809 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10809} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10737} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10529};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10838 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10892 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10936 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10554, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10401} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10892} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10838} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10936};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10710 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10653 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10433 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10573 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10988, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10842} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10410} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10433} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10573};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10819, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10684} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10653} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10710} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10988};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10554} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10610} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10819};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10939 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10939);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10690 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10568 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10774 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10568 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10828 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10774;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11029 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10786 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10917 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10515, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11011} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10786} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11029} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10917};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10513 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10981 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10763 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44729 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44729;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11008 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10782, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10656} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10763} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10981} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11008};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10629, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10492} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10513} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10515} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10782};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10401} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10629} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10684};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10649 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10640 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10497 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10675, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10543} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10640} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10649} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10497};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10702 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10862 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10870 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10655 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11005 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10566, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10417} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10655} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10870} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11005};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10946, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10808} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10862} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10702} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10566};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10427, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10923} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10675} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11011} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10946};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10842} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10427} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10492};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10424 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10848 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10724 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10832, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10694} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10848} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10424} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10724};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10996 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10583 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11026 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10715 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10443, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10935} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11026} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10583} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10715};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10480, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10974} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10443} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10996} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10417};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10601, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10455} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10832} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10543} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10480};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10656} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10601} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10923};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11010 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10776 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10598 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10717, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10591} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10776} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11010} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10598};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10726 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10512 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10739 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10960, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10824} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10512} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10726} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10739};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10928 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10439 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10686, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10557} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10928} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10439};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11000, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10853} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10686} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10960} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10935};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10748, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10621} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10717} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10694} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11000};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10808} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10748} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10455};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10483 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5978 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6099 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5978;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5909 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5909) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6099));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7318 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7419 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7318) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7375 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7419));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7555 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7375) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N687 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7555);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N687;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10452 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10454 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10469 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10792 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10925, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10784} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10469} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10454} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10792};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10613, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10470} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10452} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10483} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10925};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10860 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10926 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10833 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10581, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10432} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10926} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10860} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10833};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10881, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10740} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10557} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10581} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10824};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10644, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10505} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10591} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10613} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10881};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10974} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10644} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10621};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11019 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10807 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10528 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10893, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10750} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10807} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11019} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10528};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6403 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6210 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6210) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6403));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7516 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7362 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7516) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7320 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7362));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7498 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7320) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N686 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7498);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N686;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10944 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10822 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10597 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6412 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6412;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7418 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7462 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7418));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7562 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7462) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7518 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7562));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7446 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7518) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N685 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7446);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[1] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N685 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10805 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10544, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45592} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10597} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10822} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10805};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10845, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10709} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10944} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10893} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10544};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10660 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10593 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10569 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10811, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45621} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10593} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10660} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10569};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10495, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10991} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10784} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10811} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10432};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10530, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11028} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10845} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10470} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10495};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10530} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10853} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10505};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11007 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10556 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5928 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5928 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5643 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6040 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5832 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6040;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N623 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5643));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7360 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N623) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7407 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7360));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7506 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7407) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7464 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7506));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7390 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7464) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N684 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7390);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[0] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N684 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10673 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45631, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45618} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10556} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11007} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10673};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10476 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10458, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45584} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45631} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10476} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10750};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11016 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10913 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10890 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10609 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10558, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10408} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10890} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10609};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45595, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45581} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10913} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11016} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10558};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10827 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45774 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10445 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45774) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10630 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10671 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10902 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10825, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10688} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10671} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10630} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10902};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45624, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45608} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10445} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10827} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10825};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10729, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45612} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45595} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45592} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45624};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10759, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10635} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10458} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10709} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10729};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10759} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10740} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11028};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10731 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10722 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10645 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45583, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45569} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10722} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10731} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10645};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10987 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10620 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10787, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10661} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10987} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10620};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10560 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45611, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45598} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10560} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10787} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10408};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45587, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45572} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45583} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45618} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45611};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11013, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45576} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45584} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45621} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45587};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10991} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11013} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10635};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10451 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10633 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10461 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10434, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10927} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10633} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10451} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10461};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11001 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10907 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10972 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10706 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10398, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10895} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10972} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10706};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10711, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10582} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10907} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11001} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10398};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45575, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10883} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10688} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10434} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10711};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45615, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45601} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45608} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45581} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45575};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45612} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45615} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45576};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10990 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10683 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10804 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10679, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10548} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10683} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10990} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10804};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10718 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10814 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10428 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10538 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10918, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10775} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10428} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10538};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10951, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10815} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10814} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10718} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10918};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45620, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10847} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10661} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10679} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10951};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45604, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10534} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45569} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45598} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45620};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45572} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45604} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45601};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10519 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10712 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10533 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10625 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10865 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10970 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10500, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10995} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10865} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10970};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10617, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10477} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10625} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10533} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10500};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10889 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10430 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10894 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10449, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10940} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10430} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10889} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10894};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11006, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10858} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10617} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10712} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10940};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10994 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10444 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10839, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10700} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10444} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10994} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10775};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10516 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10619 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10967, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10829} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10516} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10619};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10797 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10781 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10416 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10801, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10670} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10781} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10416};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10720, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10596} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10797} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10967} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10670};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10547 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10708 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10574, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10423} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10708} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10547} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10801};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10487, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10980} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10449} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10720} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10423};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10700} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11006} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10980};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10637 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10604, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10462} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10637} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10895} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10574};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10872, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10732} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10548} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10839} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10815};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10462} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10487} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10732};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10636, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10496} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10927} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10582} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10604};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10872} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10847} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10496};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10883} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10636} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10534};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10436 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10517 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10979 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10882 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10764, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10639} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10979} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10517} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10882};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10885, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10743} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10829} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10436} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10764};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10885} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10596} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10858};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10540 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10788 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10693 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10600 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10930, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10789} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10693} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10600};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10412, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10909} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10788} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10995} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10930};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10477} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10412} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10743};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10450 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10962 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10422 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10676 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10765 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10817, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10681} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10676} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10765};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11020, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10422} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10962} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10817};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10523 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10699 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10947 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10415 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10734, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10606} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10947} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10415};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10585, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10438} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10699} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10523} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10734};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10789} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11020} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10438};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10585} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10639} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10909};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11015 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10874 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10504 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11037 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10898, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10504} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11037};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10605 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10465, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10605} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10898} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10681};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10874} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10606} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10465};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10888 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10618 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10953 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10510 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10749 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10852 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10627, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10749} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10852};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10510} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10953} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10627};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10692 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10481 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10587 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10840} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10481} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10587};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10840;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10861 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10790 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10982 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10861 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10790) & (!(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10414 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10816 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10982 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10414) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10584 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10692) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10816)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10969 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10966 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10584 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10969) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10479 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10650 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10966) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10618)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10479);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10745 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10950 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10650 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10888) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10745);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11035 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10672 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10871 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11035) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10672);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10472 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10950) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11015)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10871);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10942 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10975 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10472 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10450) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10942);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10747 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10975;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11036 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10747 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10540) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11036);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10674 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10945 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10674 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10575 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10575));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10697 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11014 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10697);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10519)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11014);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10828) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10690));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10723 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10785 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10873 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10545 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10873));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10978 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10545);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10659 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10978);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10961 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10785)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[32] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10723) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10961;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13228, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12514} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[32]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13228;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12514;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23314 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23314;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13204 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11971 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7963 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8238 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7963 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9061 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8076 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7922 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8076) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8941 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8868 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8504 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8868 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8607 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8941 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8504);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8200 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8607);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8238 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9061) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8200;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12992 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12850 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12373, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12008} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12992} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11971} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12850};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12246, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11873} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12373} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13010} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12800};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13262 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8264 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8722 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8415 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8722);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8108 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8264 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8415);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9070 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8203 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8849 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9070 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8203);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7885 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8803 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8849 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7885);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9055 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8673 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9055 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8972 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8673);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9096 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8803 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8972);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8108 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9096;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12651 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12510 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13207, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12834} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12651} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13262} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12510};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11738 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12369 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11751 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11759, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13046} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12369} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11738} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11751};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13076, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12726} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11759} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13207} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12923};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13028 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8751 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9005 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8751) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8981 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7946 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8440 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8981 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7946);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8014 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9005 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8440);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8551 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8877 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219)) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8809 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8060 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8809 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8327 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8382 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8060 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8327);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8287 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8877 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8382);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N753 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8287 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8551) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8014));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N753;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12290 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12006 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12620, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12254} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12290} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13028} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12006};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12009 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12009 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12751 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12953 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12145 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11885, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13177} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12751} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12145};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12283, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11911} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11885} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12620} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13046};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12159, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11784} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12008} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12283} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12726};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12950, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12611} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13076} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11873} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12159};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12337, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11974} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12246} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12888} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12950};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[37], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[36]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12275} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13204} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12337};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[37]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[37]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8508 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8013 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9068 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8013 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8612 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9124 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8393 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9124);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7993 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8393);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8243 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7993);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[18] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8508 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9068) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8612) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8243);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9042 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8052 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8695 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23415 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9042 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8052) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8695);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9095 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8477 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9095 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8589 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8477);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23415 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8589);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12710 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8775 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8034 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8775);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8081 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8720 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8081);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7926 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8034) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7926) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8720);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11994 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10638 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10499 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10638);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10908 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10800 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10411 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10800;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10411) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10908);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12038, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13331} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11994} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12611} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[36], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[35]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12710} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11974} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12038};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[18]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[36]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[36]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11775 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12399 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11814 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12224, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11853} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12399} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11775} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11814};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12880 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13298 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12684 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12547 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12015, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13313} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12684} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13298} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12547};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11667, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12959} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12880} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12224} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12015};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12181 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12042 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12042 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12780 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12567, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12200} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12780} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12181} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8402 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9135 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8660 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9135);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9079 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8402 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8660);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8208 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9079);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8515 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9013 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8293 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8906 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9013) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8293) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7932 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8515 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8906);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8208 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7932;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11921 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13062 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12324 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12041 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13283, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12902} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12324} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13062} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12041};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12730, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12378} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11921} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12567} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13283};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12406, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12047} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13177} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12254} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12730};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12982, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12645} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12834} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11667} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12406};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8485 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8307 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8808 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8307 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8326 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8596 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8326) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23407 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8808) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8596);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8485 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23407);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12906 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12859, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12524} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12982} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11784} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12906};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13067 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8214 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7897 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8214 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8796 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8987 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8796 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8994 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8170 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8994);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7951 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7897 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8987) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8170;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8428 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8044 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8686 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8275 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8126 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8686 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8275);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8932 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8428 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8126);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7951 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8932;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13213 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12920 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & N23928) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & N23926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12434 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11874 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | N23926);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | N23928);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12775 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12470 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12392} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12775} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12470};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12909 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13095, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12737} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11874} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12434} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12909};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12349, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11986} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12920} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13213} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13095};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11791, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13084} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12349} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11853} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13313};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13113, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12756} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11791} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12959} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12047};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12072, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11694} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11911} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13113} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12645};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11943, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13235} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12072} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13067} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12524};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[35], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[34]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12859} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13331} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11943};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9102 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8679 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7996 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8268 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8114 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7996 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8268);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8372 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8679) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8114);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[17] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9102 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8372);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[17]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[35]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[35]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9133 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8148 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9133 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8292 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9051 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8555 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8292 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9051);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8639 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8881 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8639);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8401 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8232 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8658 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8881) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8401) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8232);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[16] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8148) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8658);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12711 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11807 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13335 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12873, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12540} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11807} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12711} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13335};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12583 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8342 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8300 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9141 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8300);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8135 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8196 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8135);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8891 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8564 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8891);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8155 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8196 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8564);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8963 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9141 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8155);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8236 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9017 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8236);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8030 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8842 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9017 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8030);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8665 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125)) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8842);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8963 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8665;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12843 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11963 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11962, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13253} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12843} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12583} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11963};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13054, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12706} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12873} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12200} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11962};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13100 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12358 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12074 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11774, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13061} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12358} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13100} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12074};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12216 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12572 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8435 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9093 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8865 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9093) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8694 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8435 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8865);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8220 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8474 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7902 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8220) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8474);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8175 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7902 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8175 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8694;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12503 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12714, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12357} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12572} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12216} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12503};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12683, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12323} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12714} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11774} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12737};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12139, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11765} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11986} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12902} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12683};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12532, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12165} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13054} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12378} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12139};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8538 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8124 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8538));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8858 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8815 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8858 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8986 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7950 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23399 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8815 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8986) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7950);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8124 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23399);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8784 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8400 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8514 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8400 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8952 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8656 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8086 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8952 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8656);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[16] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8784) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8514) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8086);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13125 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12193, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11821} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12532} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12756} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13125};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10971 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10971) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10475 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10475);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10713 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10854 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10498 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10854 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10849 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10498;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45208 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45200 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45208)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45200);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10849) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10713);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12798 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12798 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28] ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45526 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45206 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45530 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45206;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45530) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45526);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11779 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11779 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13244, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12867} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13084} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12165} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12365 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12894, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12561} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13244} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12188} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12365};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11844, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13140} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11694} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12193} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12894};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12205 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12718 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12778, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12431} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12205} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12718};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[34], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[33]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11844} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13235};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[16]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[34]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[34]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9033 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8580 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8794 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8254 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7896 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8794) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8254);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8212 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8305 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8212);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8426 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8305);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[15] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9033 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8580) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7896) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8426);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9138 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9085 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9138);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8887 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8960 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8644 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7957 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8153 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8644 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7957) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7983 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8960 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8153);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8352 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7983);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9085) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8887) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8352);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12415 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13254 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12951 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11842 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12745 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11809, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13099} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12392} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11842} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12745};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12509, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12147} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12951} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13254} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11809};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11740, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13027} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12540} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13253} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12509};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12842, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12502} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12706} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11740} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11765};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11812 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12316, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11953} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12842} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12415} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11812};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23307 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23307;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12004 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12874 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11697 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8321 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8648 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8321);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8439 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8944 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8439);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9063 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8648 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8944);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8202 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9063);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8873 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7965 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8873);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8179 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8241 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8179 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8896 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7965 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8241);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8056 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8507 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8056);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8771 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8507 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7924 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8896 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8771);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8202 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7924;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12136 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12546, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12180} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11697} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12874} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12136};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13224, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12849} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12546} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12357} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13061};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12476, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12114} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12323} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13224} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13027};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8360 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8864 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8360) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8316 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8655 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8316 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8413 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8472 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8413) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8174 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8472);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8864 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8655) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8174);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11682 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11920, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13215} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11682} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12476} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12502};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13018, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12677} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12004} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12867} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11920};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11980, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13275} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11821} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12316} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13018};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[33], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[32]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12431} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11980} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13140};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[15]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[33]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[33]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13103 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12716 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12716 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23303 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25] ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23303;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12925 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8630 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8110 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8973 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8851 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8574 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7994 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8851 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9099 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8973 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7994);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8368 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8110 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9099);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8630 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8368;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11766 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12986 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13290 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12368, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12005} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12986} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11766} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13290};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13133 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12391 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & N23928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12110 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13300, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12919} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12391} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13133} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12110};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12333, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11970} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13300} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12368} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13099};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11996 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12614 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12250 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12426 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12537 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12582, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12217} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12426} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12250} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12537};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13261, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12882} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12614} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11996} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12582};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12297, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11930} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13261} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12333} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12147};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10588 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10588) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10875 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10733 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10949 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10603 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10459 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10603) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10949)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10459);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[23] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10733) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10875);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[23];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11683 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23226 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11683 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23226;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13185, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12818} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12297} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12114};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12653, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12289} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12925} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13103} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13185};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8346 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9062 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8827 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8075 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8827);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8895 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9062 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8075);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8388 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8455 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8388) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8346 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8895) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8455) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12630 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8398 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8781 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8398);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8247 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8315 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9128 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8315);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7973 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9128);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8512 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8247 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7973);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8512;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13055 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12774 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12648 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12613, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12249} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12774} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13055} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12648};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11875 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12589 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12803, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12464} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11875} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12589};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12910 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11732 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12171 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13334, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12952} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11732} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12910} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12171};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13068, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12722} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12803} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12613} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13334};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13034, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12691} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12180} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13068} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12882};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12999, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12661} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12849} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13034} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11930};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12588 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12263, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11893} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12999} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12630} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12588};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13295 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11702, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12991} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13295} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12263} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13215};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12106, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11728} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12653} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11953} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11702};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[32], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[31]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12106} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12561} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13275};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8938 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8071 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8384 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8496 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8384);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8473 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9113 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8473 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8133 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7901 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8823 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7901);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8610 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9113 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8133) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8823);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[14] = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8938 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8071) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8496) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8610;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[14]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[32]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[32]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8046 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8046);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8404 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8839 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8956 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8839);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8067 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8786 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8956) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8067);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[29] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8404) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8786);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8582 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8913 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8687 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8913);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8640 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8582) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8687;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8215 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8378 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8215) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[28] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8378);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313 = 1'B0 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8565 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8031 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7920 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8409 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8031) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7920) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8892 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[27] = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8565) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8409) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8892);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[27]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8437 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8222 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8050 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8176 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8222) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8050) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[26] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8437 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8176);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[26]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8588 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8079 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8588);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8348 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7966 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8459 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8348 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7966);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9065 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8650 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7925 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9065) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8650);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8897 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[25] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8079 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8459) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7925) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8897);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[25]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810 = !(N23926 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[42] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8975 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8369 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8975) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8632 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8369) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8924 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8531 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8747 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8924 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8531);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8267 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[24] = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8632) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8747) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8267);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[42]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[24]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9007 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8018 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9007 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8121 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8755 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8121);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8880 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8755);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8834 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8880));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8183 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8489 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8704 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8489;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8553 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8183) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8704) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9131 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8834 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8553);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[23] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8018 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9131);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[41] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[42];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[41]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[23]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[41]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15428 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12918 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12749 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12965, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12626} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12749} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12918} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12818};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45799 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45799 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12826 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[23] ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12826;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12046 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12397 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12791, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12447} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12046} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12661} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12397};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9097 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8479 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9097);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8204 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8675 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8204);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9025 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8627 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9025 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8922 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8971 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7941 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8922 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8971);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8319 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7941) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23391 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8675 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8627) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8319);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8479 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23391);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11898 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12155, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11782} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12217} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12919} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12005};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13170 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12284 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12646 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12837, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12497} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12284} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13170} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12646};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12033 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12573 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12427 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8423 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8464 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8272 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8423 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8464);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8120 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8272 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8251 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8856 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8251 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8355 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7892 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8355 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8811 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8856 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7892);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8682 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8983 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8682);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9106 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8811 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8983);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8120 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9106;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12704 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12647, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12285} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12427} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12573} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12704};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12400, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12040} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12033} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12837} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12647};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11800 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13020 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13328 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11696, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12985} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13020} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11800} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13328};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13107, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12750} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11696} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12464} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12952};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12857, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12516} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13107} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12400} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12722};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12123, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11747} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12155} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11970} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12857};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12220 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12088, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11711} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12123} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11898} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12220};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12053, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11676} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12088} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12791} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11893};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12438, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12081} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12965} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12289} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12053};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[31], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[30]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12677} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12438} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11728};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8160 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8524 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8160) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8568 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9023 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8946 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8524 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8568) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9023);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8361 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8946);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7883 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9090 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8103 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7883 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9090);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[13] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8361 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8103);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[13]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[31]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[31]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45780 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45780) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10954 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10464 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21] = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10464) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10954);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13252 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13252 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9126 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8395 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8065 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7970 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8065);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9009 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7970);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8779 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8395 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9009);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23383 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9126 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8779);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8702 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8244 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8702);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23383 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8244);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12821 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12823, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12481} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12691} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12821};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12579 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13093 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9015 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8191 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8445 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8295 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8191 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8445);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8884 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7915 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8916 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8884 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7915);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8560 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8295 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8916);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9015 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8560;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12350 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12804 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11957, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13247} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12350} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13093} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12804};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12352 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11916 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12870, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12534} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12352} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11916};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12207 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12942 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12069 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12679, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12318} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12942} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12207} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12069};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12433, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12073} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12870} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11957} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12679};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12189, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11815} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12249} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12433} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12040};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11938, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13231} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11782} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12189} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12516};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11846 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11901, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13192} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11747} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11938} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11846};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11863, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13157} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12579} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12823} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11901};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12037 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11668 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12213 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12632, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12269} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12037} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11668} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12213};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12601, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12232} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11711} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12632} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12447};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12761, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12411} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11863} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12626} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12601};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[30], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[29]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12991} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12761} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12081};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8480 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8696 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8480) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9045 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8009 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9045);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8674 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9098 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8999 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8674 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9098;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8282 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8009 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8999);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[12] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8696 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8282);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[12]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[30]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[30]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13142, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12779} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12285} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12497} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12985};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12738 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13208 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11836 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12707, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12351} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13208} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12738} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11836};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12472, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12109} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12707} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12534} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13247};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8914 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8199 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8469 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8199);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8862 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8914 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8469);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8666 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7986 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8735 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8666 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7986);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8099 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9037 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8099 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8845 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8735 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9037);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8172 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8862 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8845);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8312 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8420 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8429 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8420);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8429 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8172;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11987 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12463 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12606 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11990, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13286} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12463} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11987} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12606};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12680 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12319 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13285 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12202, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11829} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13285} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12319} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11731, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13022} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12680} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11990} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12202};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12221, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11848} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11731} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12472} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12073};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12889, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12554} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13142} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12750} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12221};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8726 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8576 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8726);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8271 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8576);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8907 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8422 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8907);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8535 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8422);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8855 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7998 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8855);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8271) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8535) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7998);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12121 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13138 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12666, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12306} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12121} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12889} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13138};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12958 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23421 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23421 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21] ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12784 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13333 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11717, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13003} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12784} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12958} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13333};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11685, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12970} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12481} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12666} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11717};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10549 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10680 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10680) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10549));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10820 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10820) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13149 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13149);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8334 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7913 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8022 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7913);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8838 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8334) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8707 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8838) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8707) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13031 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11976, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13267} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11815} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13031};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11841 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12456, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12095} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11841} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11976} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13231};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12417, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12061} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13192} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12456} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12269};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13323, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12938} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11685} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13157} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12417};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[29], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[28]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11676} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13323} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12411};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8350 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8144 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8614 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8350 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8144);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8900 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8552 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8082 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8552);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8778 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8245 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7927 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8778 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8245);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[11] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8614 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8900) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8082) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7927);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[29]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[11]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[29]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12619 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12440 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12948 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11753, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13039} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12440} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12619} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12948};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12384 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13127 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12836 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12940, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12603} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13127} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12384} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12836};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11689 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11954 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8766 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8280 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9060 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8280 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8197 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9060);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8033 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8766) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8197);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8715 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9117 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8073 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9117 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8136 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8344 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8136 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8452 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8073 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8344);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9019 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8715 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8452);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9019 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8033;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13281 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13158, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12793} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11954} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13281};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11768, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13058} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11689} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12940} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13158};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13180, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12811} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12318} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11768} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13022};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12927, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12592} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12779} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13180} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11848};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12777 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12696, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12339} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12554} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12927} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12777};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13162, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12796} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12696} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11753} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12306};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13132 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8733 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9087 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8619 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8045 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9087 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8619);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7985 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8213 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7985 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8376 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8213);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8733) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8045) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8376);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12329 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12240 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12978 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12101 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12027, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13326} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12978} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12240} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12101};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12505, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12141} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12027} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13286} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11829};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12023 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12498 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12640 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12271, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11903} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12498} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12023} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12640};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11830 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12903 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13195, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12825} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11830} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12903};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12765 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13248 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11867 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12973, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12633} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13248} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12765} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11867};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12740, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12386} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13195} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12271} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12973};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13217, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12844} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12351} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12740} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13058};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12256, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11888} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12505} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12109} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13217};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45525 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12152 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45525) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26]) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12152;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12432 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12010, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13306} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12256} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12329} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12432};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12490, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12129} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13267} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13132} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12010};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12239, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11869} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13003} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12490} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12095};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13126, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12768} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13162} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12970} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12239};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[28], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[27]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12232} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13126} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12938};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8373 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9048 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8061 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8373) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9048) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9105 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8752 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9105);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8328 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8752) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[10] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8061 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8328);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[10]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[28]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[28]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12255 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12610 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11786, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13078} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12255} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12592} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12610};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12079 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20]) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20] ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11892 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10631 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[18] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10631) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[18] & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11803, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13097} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12603} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12793} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13326};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12134 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13011 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12056 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12939 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13043, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12698} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12056} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12939};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12098, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11720} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13011} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12134} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13043};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13163 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12871 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12277 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13006, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12667} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12871} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13163} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12277};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12770, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12420} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13006} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12098} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11903};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13324 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12762 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12418 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12308, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11940} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12762} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13324} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12418};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11723 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12064, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11686} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12308} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12825};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12541, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12174} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12064} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12770} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12386};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12291, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11924} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11803} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12141} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12541};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12961, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12622} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12811} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12291};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12727, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12375} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11892} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12079} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12961};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13199, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12830} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12727} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11786} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12339};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12771 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9115 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7960 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8436 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8763 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8436 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8684 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8499 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8684);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[6] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9115 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7960) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8763) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8499);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13260 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12071 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12049, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11670} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11888} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13260} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12071};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11701 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13187 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11883 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12758, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12407} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13187} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11701} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11883};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12527, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12161} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12049} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12771} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12758};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12279, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11907} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13039} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12527} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12129};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12945, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12605} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13199} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12796} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12279};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[27], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[26]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12061} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12945} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12768};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8294 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8955 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7980 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8955 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7914 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8708 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8403 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8250 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7914) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8708) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8403;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[9] = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8294 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7980) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8250;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[9]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[27]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[27]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13237, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12861} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13306} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12375} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13078};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12424 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12248 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45786 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10755 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45786) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45792 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10897 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45792) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10897) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10755);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11908 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12797 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11760 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12832, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12493} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12797} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11908} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11760};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12062 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12533 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12673 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12131, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11756} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12533} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12062} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12673};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12799, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12458} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12131} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12832} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11940};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11839, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13129} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12633} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12799} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11686};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13258, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12876} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13097} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11839};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12659 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12995, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12654} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12844} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13258} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12659};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11824, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13115} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12248} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12424} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12995};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8968 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8526 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8800 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8526);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8848 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8262 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8848 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8414 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8719 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8669 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8414 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8719);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[5] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8968 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8262) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8669);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12543 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11692 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12083, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11705} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12543} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11924} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11692};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12817 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12993 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13176 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12786, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12441} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12993} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12817} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13176};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12563, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12194} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12083} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12622} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12786};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12312, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45350} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12563} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11824} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12161};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12977, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12639} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13237} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12830} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12312};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[26], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[25]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12977} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11869} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12605};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8012 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8127 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8012);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8734 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8621 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8098 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8860 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8098);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8171 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8539 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8734 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8621) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8860) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8171;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9110 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8539);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[8] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8127 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9110);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[8]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[26]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[26]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9116 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8498 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9116 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8343 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8498);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8604 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8237 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8005 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8893 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8005;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8451 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8237 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8893);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8324 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8451);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[7] = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8343 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8604) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8324;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11872 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12068 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12265 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12703, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12347} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12265};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12966 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11684 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12864, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12529} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12966} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12703} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11684};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13200 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12453 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12313 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11948, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13241} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12453} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13200} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12313};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11909, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13202} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12864} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12698} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11948};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11870, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13165} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12667} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11720} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11909};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13033 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12575, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12211} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13033} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11870} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12420};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12296 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12326, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11966} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12575} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12174} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12296};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11856, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13150} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12068} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11872} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12326};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13276, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12897} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11670} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12407} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11856};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9122 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8872 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8594 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8700 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8390 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8700) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23375 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8872 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8594) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8390);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9122 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23375);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11806 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12983 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13029, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12687} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11806} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12876} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12983};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12652 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12475 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12809 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12118, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11742} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12475} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12652} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12809};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12596, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12226} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13029} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12654} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12118};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45345, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45394} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13115} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12596} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12194};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13012, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45377} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13276} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12861} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45345};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[25], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[24]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11907} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13012} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12639};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[25]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[7]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[25]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13166 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12332 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12167 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13050 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12971 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12096 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11762, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13052} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12971} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12347} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12096};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12675, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12314} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13050} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12167} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11762};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12642, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12281} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11756} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12675} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12493};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12607, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12243} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12332} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12458} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12642};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13293, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12913} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12607} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13129} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12211};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11687 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12819, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12479} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13293} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13166} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11687};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13315, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12933} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12819} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12441};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12829 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12702 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11944 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12501, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12135} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12702} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12829} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11944};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11725, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13015} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12501} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12529} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13241};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13263 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11691, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12981} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11725} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13202} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13263};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13329, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12946} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13165} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11691} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12243};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12116 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12469 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13064, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12717} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12116} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13329} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12469};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11932 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8397 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7930 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8397 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8016 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8903 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8016);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8948 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9073 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8948);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7974 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8461 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7974);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[3] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7930 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8903) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9073) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8461);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12742 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12644 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12361, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12000} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12742} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11932} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12644};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11896, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13189} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11966} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13064} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12361};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45389, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45721} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13150} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11896} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12226};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45371, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45358} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13315} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12897} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45389};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[24], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45342} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45350} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45371} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45377};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9024 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7938 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9024) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9041 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7938);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8221 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8364 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8051 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8364);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8318 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8221) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8051) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[6] = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9041 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8318);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[6]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[24]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[24]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15184 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12461 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12105 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12637 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12183, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11810} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12105} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12461} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12637};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11934, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13227} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12000} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12183} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12717};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12099 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11729 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11718 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13190 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12491 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12321, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11959} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13190} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11718} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12491};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11794 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13086 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13238 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12344 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13025, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12682} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13238} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13086} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12344};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13210, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12840} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11794} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12321} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13025};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12545 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12467, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12103} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13210} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12314} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12545};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12429, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12070} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12281} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12467} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12981};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12922, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12585} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11729} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12099} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12070};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8374 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8813 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8167 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8636 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8167 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8488 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8813 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8636);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9032 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8488);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8374) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9032);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12029 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13223 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12282 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12394, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12035} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13223} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12029} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12282};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11739 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11922 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13102, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12747} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11739} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12429} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11922};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11973, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13264} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12035} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12922} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12747};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12511 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11808 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11752 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11743 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12526 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12969, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12629} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11743} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11752} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12526};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11983 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12478 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13004 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11927, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13220} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12478} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13004};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11708, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12997} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11983} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12969} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13220};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12732 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12130 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12862 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12656, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12295} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12130} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12732} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12862};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12112, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11735} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11927} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12656} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11959};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12814, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12474} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12682} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11708} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11735};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12989, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12649} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12840} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11808} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12814};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8540 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8990 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8820 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8736 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8380 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8736 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8094 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8380);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8933 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8820 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8094);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9036 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8003 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9036 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23367 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8990 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8933) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8003);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8540 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23367);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8446 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8957 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8446);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8023 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8516 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8023);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8790 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8709 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7981 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9081 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7981);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8089 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8709 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9081);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[1] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8957 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8516) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8790) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8089);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12237 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12251, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11880} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12989} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12511} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12237};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12274 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12685 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12841 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13205 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12955, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12617} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12841} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12685} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13205};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12007, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13302} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12274} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12251} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12955};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12287, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11918} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13052} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12135} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12112};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13173, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12805} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13015} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12287} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12103};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13026 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13214 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12219, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11843} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13026} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13173} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13214};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12941 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12848 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11912 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13135, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12776} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12848} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12941} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11912};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12884, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12549} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12219} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12946} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13135};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12693, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12335} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11810} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12007} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12549};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45718, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45705} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11973} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13227} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12693};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12853, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12512} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12394} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12913} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13102};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45711, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45698} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12853} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12479} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13189};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12975 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12288 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12802 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12150, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11778} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12288} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12975} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12802};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12628, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12264} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12687} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12150} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11742};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45692, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45679} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12884} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12512};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45708, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45695} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11934} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12264} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45692};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45677, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45724} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45698} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45718} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45695};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8879 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8017 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8879);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8331 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8442 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8290 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8331) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8442) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8063 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8184 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8063);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8978 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8184);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45700 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8017 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8290) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8978) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45353, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45687} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12628} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12933} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45711};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45380, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45713} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45721} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45708} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45687};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45700} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45677} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45713};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7929 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8418 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8976 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8418);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9074 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8163 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9074);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8266 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8163);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8852 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8634 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8852);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45391 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8976 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8266) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8634;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45400, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45386} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45394} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45353} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45358};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45391} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45380} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45386};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8150 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8663 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8150);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8091 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8663);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9030 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8297 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8789 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8297);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8616 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8789);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8727 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8616 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8038 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45720 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8091 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9030) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8038;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13017 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11722 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12044, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13337} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13017} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12805} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11722};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12723, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12371} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12044} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12776} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11843};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13159 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12146 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12075, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11699} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11918} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13159} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12146};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11904 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12380 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13277 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12688 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13040 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12389, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12030} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12688} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13040};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12059, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11681} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13277} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12380} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12389};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12444, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12087} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12295} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12059} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12997};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12746 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11890, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13183} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12746} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12444} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12474};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12833 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12783, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12437} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11890} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12649} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12833};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12752, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12404} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11904} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12075} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12783};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11783, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13071} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12752} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12585} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13302};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45668, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13036} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13264} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11783};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45684, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[19]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45679} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45668} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45705};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45684} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45720} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45724};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8874 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45383 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8874 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45368 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8180 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45341 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8180 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8699 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8322 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9121 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8699) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8322;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45355 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9121 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45397 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45383 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45368) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45341) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45355);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45397} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45400} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45342};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8157 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8843 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8453 = ((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8303 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8453);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8303 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8566 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[0] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8157 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8843) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8410) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8566);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12504 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12325 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12676 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11851, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13143} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12325} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12504} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12676};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11818, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13109} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11851} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11880} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12617};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12137 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11961 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12317 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11673, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12964} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11961} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12137} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12317};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13310, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12930} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11699} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11673} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12437};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12669 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12828 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12409, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12051} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13183} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12669} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12828};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12896 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12162 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12016 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13098, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12741} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12162} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12896} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12016};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12764, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12416} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13098} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12629} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11681};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12032 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13154, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12789} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12764} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12087};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12133 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13255 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12935, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12599} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12133} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12789} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13255};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12943 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11787 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11965 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12564 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13229, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12854} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11965} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11787} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12564};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12178, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11805} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13229} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12030} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12741};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11833, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13124} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12178} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12943} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12416};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13063 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12229, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11859} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11833} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13063};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11951 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11764 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12311 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12021, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13319} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11764} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11951} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12311};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13119, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12759} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12229} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12935} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12021};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12377, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12011} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12409} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13143} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13119};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13270, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12891} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13310} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13109} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12377};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13198 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13008 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11773 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12496 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12625, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12259} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11773} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13154} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12496};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12593, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12223} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13008} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13198} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12625};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12557, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12190} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13337} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12593} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12404};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12520, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12157} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11818} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12371} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12557};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[18], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[17]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13071} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13270} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12157};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[18]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[19], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[18]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12335} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12520} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13036};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12712 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12241 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12877 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13077 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12423, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12067} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12877} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13077};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13316 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12304, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11937} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13316} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12423} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12854};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12879, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12544} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12241} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11805};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12571, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12204} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12879} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12712} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13124};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12487 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12734, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12381} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12487} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12571} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11859};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12196, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11826} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12259} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12964} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12734};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13080, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12729} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12223} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12930} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12196};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[17], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[16]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12190} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13080} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12891};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[17] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8991 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8379 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8991);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7899 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8492 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7899 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8935 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8313 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7953 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8935 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8277 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8689 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8819 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8689);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8234 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8277 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8819);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[1] = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8379 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8492) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7953) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8234);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[1]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[19]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15524 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444 = !(N22905 | N23646);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15035 = !(N23051 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13047 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12356 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12538 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12689, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12328} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12356} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13047} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12538};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12868 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12705 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13233 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11746, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13032} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12705} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12868} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13233};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13060, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12709} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12689} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12204} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11746};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12536, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12169} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13319} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13060} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12381};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12934 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12195 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11822 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12175 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12595 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13038, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12694} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12175} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11822} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12595};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13131, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12773} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12195} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12934} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13038};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13161 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13002, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12664} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13131} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11937} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13161};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11968, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13259} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13002} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12544};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13243 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11942 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12355, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11993} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13243} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11968} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11942};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12875 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11757 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13056 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13289, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12907} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11757} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12875} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13056};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11796, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13092} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13289} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12355} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12599};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12900, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12566} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12051} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11796} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12759};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[15], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[14]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11826} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12536} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12566};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[16], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[15]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12900} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12011} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12729};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[16] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15141 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[15] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12454 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12214, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11840} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12067} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12773} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12454};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11997 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12093, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11716} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12214} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12664} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11997};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13096 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13116 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12039, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13332} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13096} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13116};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12227 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11857 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12387 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13148 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13327 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12860, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12523} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13327} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13148} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12460, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12100} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12387} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11857} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12860};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12748, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12396} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12227} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13332} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12460};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12128, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11749} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12039} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12694} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12748};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12917, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12578} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12128} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11840};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12700 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12172 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12794, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12451} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12700} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12917} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12172};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12480, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12120} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12093} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13259} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12794};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12143, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11771} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12907} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11993} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12480};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[14], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[13]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12143} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13092} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12169};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[14] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12531 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12348 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11866, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13160} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12348} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12531} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11716};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13191, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12820} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12328} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11866};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[13], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[12]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12709} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13191} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11771};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15155 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[13] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15456 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15155;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12164 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11988 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12720, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12364} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11988} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12164} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12578};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12343 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13291 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11801 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12003, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13296} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13291} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12343} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11801};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12604, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12236} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12003} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12720} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12451};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[12], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[11]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12120} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12604} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12820};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15531 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[12] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13094 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12665 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11811, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13106} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12665} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12396} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13282 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11906, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13197} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11811} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13094} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13282};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11719 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12908 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12827, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12488} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11719} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11749} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12908};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11781, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13066} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12827} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11906} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13296};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[11], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[10]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13160} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11781} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12236};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[11] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11792 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12736 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12574 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12901 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12552, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12187} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12574} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12736} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12901};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12636, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12273} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11792} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12488} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12552};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[10], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[9]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12364} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12636} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13066};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14950 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[10] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[10]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13083 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11939 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12208 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13169, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12801} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12100} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12208};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13266, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12886} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13083} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13106} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13169};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[9], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[8]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13266} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13197} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12273};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15322 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[9] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12856 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11941, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13236} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12523} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12856} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12385 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12247, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11871} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11941} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12568} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12385};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[8], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[7]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12247} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12187} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12886};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15038 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[8] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12024 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11835 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12198 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12670, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[5]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11835} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12024} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12198};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[7], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[6]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12801} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12670} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11871};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15403 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[7] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12154 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12602 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13128 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13074, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[4]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12602} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12154} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13128};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13322 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13069 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13305, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12924} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13069};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12766 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12367 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13299 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11845, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[1]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13299};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12587, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[2]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12367} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11845};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12374, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[3]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12766} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12924} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12587};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12160, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[4]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13305} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13322} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12374};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[6], DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[5]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13236} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13074} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12160};
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[6] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15492 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[5] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15201 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[4] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[3] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15580 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[3] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[2] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[2] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[1] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15519 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[1] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[1]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15144 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[2] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15129 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15519 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15144);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15270 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[1] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[1]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14960 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15129 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15270);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15429 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[3] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15453 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14960 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15580) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15429);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15199 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15201) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15453)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[4]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[4]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15345 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[5] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14974 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[6] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14994 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15345) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14974;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15068 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15492) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15199) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14994);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15257 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[7] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15023 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15068) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15403)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15257);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15556 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[8] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14970 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15023 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15038) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15556);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15177 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[9] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15498 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14970) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15322)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15177);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15466 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[10] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[10]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15097 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[11] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15327 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15466) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15097;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15485 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14950) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15498) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15327);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15379 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[12] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15560 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15485) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15531)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15379);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15011 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[13] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15298 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[14] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15311 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15011) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15298;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15084 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15560 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15456) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15311);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15590 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[15] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15210 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[16] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15000 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15590 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15210);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15084) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15141)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15000);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15297 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15412 = !N22772;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[17] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15376 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15044 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303 = ((!N22903) & (!N23646)) | (!N22875);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15424 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108) & (!(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15032 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15424);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15283 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15032);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15553 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303 & N23051) | N23049);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[49] = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15412) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15035)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15553);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[49];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45117 = !(N21282 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15143 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15565 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15490 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091 = !((N23630 & N23628) | N23103);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15409 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091) & (!N22793)) | (!N22791);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15081 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15391 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15137 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15391);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15399 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15001 = ((!N21688) & (!N23640)) | (!N23638);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15366 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015 & N21470) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15001;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45155 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15366 ^ N21279;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45117 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45155);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15064 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587 = !((N23103 & N23101) | N23099);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181 = ((!N22891) & (!N22889)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14966 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[28] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181 ^ N22648;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[28] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15550 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15352 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15207 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469 = ((!N22899) & (!N22897)) | (!N22895);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15397 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[29] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469 ^ N22621;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[29] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45835 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15338 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15019 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14940 = !(N22850 | N23620);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15539 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15195 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15457 = ((!N22852) & (!N22850)) | (!N22848);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14940) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15457);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[45] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056 & N22624) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056) & N22626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[45] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45829 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15054 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15386 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15312 = !(N22835 | N23601);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15241 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15573 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15166 = ((!N22837) & (!N22835)) | (!N22833);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15312) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15166);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[44] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426 & N22583) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426) & N22585));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[44] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45847 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15518 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15265 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15463 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15127 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383 = ((!N22868) & (!N22866)) | (!N22864);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15448 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15515 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15113 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15515);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15369 = ((!N22919) & (!N23608)) | (!N23606);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383 & N22682) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[47] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972 & N22559) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972) & N22561));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[47];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45841 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15226 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14981 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15175 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15499 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102 = ((!N22860) & (!N22858)) | (!N22830);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15161 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15223 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15487 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15223);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15086 = ((!N22826) & (!N23615)) | (!N23613);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102 & N22672) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15086);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[46] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342 & N22552) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342) & N22554));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[46] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45811 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15110 = !(N22873 | N23646);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978 = ((!N22907) & (!N22905)) | (!N22903);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14963 = ((!N22875) & (!N22873)) | (!N22871);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15110) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14963);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[41] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225 & N22597) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225) & N22599));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[41] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15483 = !(N22978 | N22793);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14985 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15334 = ((!N22791) & (!N22978)) | (!N21688);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14985 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15483) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15334);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45805 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15534 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[40] = !((N22594 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45805) | ((!N22594) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[40] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45817 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15135 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15473 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15393 = !(N22800 | N22910);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15152 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15008 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261 = ((!N22883) & (!N22881)) | (!N23137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330 = !((N23043 & N23041) | N23039);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14992 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15249 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330) & (!N22800)) | (!N22798);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15393) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15249);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[42] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516 & N22545) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516) & N22547));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[42] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45823 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15420 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15105 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15028 = !(N22814 | N22985);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15435 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15290 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562 = ((!N22845) & (!N22843)) | (!N22841);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14956 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15278 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15543 = ((!N22816) & (!N22814)) | (!N22812);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15028) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15543);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[43] = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140 & N22538) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140) & N22540));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[43] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15100 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15190 = !(N22992 | N22866);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15505 = !N22868;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15052 = ((!N22864) & (!N22992)) | (!N22919);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15308 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15505 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15190) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15052);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[39] = (!N22636) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15308;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23358 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[39] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23358;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15325 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15571 = !(N22828 | N22858);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15354 = !N22860;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15416 = ((!N22830) & (!N22828)) | (!N22826);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15026 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15354 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15571) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15416);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[38] = (!N22566) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15026;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[38] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15123 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14988 = !(N23601 | N22889);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15071 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15510 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587) & (!N23601)) | (!N22837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15107 = !((N22973 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14988) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15510);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[36] = (!N22728) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15107;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23255 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[36] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23255;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15559 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15275 = !(N23620 | N22899);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15211 = !N22897;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15132 = ((!N22895) & (!N23620)) | (!N22852);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15390 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15211 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15275) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15132);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[37] = (!N22641) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15390;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23324 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[37] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23324;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15372 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[32] = N22651 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[32] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567 = !((N22772 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23433 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15147 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[33] = !((N22575 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23433) | ((!N22575) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[33] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15583 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15078 = !(N22910 | N22883);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15441 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15594 = ((!N23137) & (!N22910)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15187 = !((N22708 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15078) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15594);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[34] = (!N22533) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15187;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[34] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15358 = !(N22985 | N22845);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15589 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15215 = ((!N22841) & (!N22985)) | (!N22816);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479 = !((N22764 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15358) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15215);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23439 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15348 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[35] = !((N22530 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23439) | ((!N22530) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[35];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14944 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[31] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383 ^ N22611;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[31] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15170 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[30] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102 ^ N22606;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[30] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15419 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173));
assign N23929 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[26] = !((N22491 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261) | ((!N22491) & N23929));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[26] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14991 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[25] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978 ^ N22616;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[25] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16497 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15192 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[27] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562 ^ N22580;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[27] & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16534 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16552 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16497)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16534);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16522 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16542 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16522);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16562 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16493 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16542) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16562);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16537 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16552)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16493);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16548 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16569 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16548);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16500 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16519 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16569) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16500);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16489 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16509 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16526 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16546 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16509) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16526);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16488 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16519) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16546);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16516 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16537 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16488);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16535 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16] | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16554 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16486 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16535) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16554);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16564 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20] | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16557 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16514 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16564) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16557);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16553 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16486) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16514));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16516) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16553);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0] = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16556 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16506 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16525 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16556 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16506);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16515 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16533 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16551 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16515 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16533);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45547 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16525) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16551);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16541 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16561 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16492 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16541 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16561);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45552 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16492;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45547) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45552);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45549 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45549;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45000 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16508 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16545 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16566 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16508) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16545);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16504 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16566)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16504);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16643 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16643 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45000) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23240 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23239 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23240 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23239));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16663 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16719 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16663) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16662 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16719));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45854 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16646 = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45854) | (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[4] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16646;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16754 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16754;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16727 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16662) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16742 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16684 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16742));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16684) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[2] = (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636) ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N683 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16727));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17223 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N683 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[22] = !((N23918 & N23924) | ((!N23918) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17223));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16790 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16685 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16790) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16789 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16685));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16693 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16789) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755 | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16704 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16809 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16809) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N682 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16693));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17207 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N682 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[21] = !((N23922 & N23924) | ((!N23922) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17207));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16810 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16756 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16810));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16817 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16756) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[3] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16668 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16775 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16668));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16775) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N681 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16817));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17267 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N681 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[20] = !((N23919 & N23924) | ((!N23919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17267));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16776 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16718 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16776));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16783 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16795 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16741 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16795));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16741 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N680 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16783));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17251 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N680 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[19] = !((N23921 & N23924) | ((!N23921) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17251));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16703 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16703 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N679 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17234 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N679 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[18] = !((N23920 & N23924) | ((!N23920) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17234));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16667 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16667 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N678 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17217 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N678 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[17] = !((N23921 & N23924) | ((!N23921) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17217));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16794 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16794 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N677 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17202 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N677 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[16] = !((N23919 & N23924) | ((!N23919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17202));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319 = !DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16724 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16724 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N675 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17244 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N675 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[14] = !((N23921 & N23924) | ((!N23921) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17244));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16691 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16691 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N674 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17227 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N674 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[13] = !((N23918 & N23924) | ((!N23918) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17227));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16814 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16814 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N673 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17211 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N673 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[12] = !((N23920 & N23924) | ((!N23920) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17211));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16762 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16762);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16746 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16746 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N672 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17270 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N672 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[11] = !((N23918 & N23924) | ((!N23918) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17270));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N671 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17254 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N671 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[10] = !((N23920 & N23924) | ((!N23920) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17254));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N670 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17237 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N670 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[9] = !((N23922 & N23924) | ((!N23922) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17237));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N669 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17220 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N669 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[8] = !((N23919 & N23924) | ((!N23919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17220));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N668 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17205 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N668 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[7] = !((N23920 & N23924) | ((!N23920) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17205));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N667 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17263 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N667 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[6] = !((N23922 & N23924) | ((!N23922) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17263));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N666 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17247 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N666 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[5] = !((N23919 & N23924) | ((!N23919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17247));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N665 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17230 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N665 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[4] = !((N23920 & N23924) | ((!N23920) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17230));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17213 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731;
assign x[3] = !((N23918 & N23924) | ((!N23918) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17198 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820;
assign x[2] = !((N23921 & N23924) | ((!N23921) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17198));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17256 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752;
assign x[1] = !((N23921 & N23924) | ((!N23921) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17256));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17239 = (DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680;
assign x[0] = !((N23919 & N23924) | ((!N23919) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17239));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16343 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128) & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N585 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16343;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N595 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N585 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[30] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N595 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N713 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[4];
assign x[27] = (N20596 & N20746) | (N20748 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N713);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N712 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[3];
assign x[26] = (N20596 & N20746) | (N20748 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N712);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N711 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[2];
assign x[25] = (N20596 & N20746) | (N20748 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N711);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N710 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759;
assign x[24] = (N20596 & N20746) | (N20748 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N710);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N709 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722;
assign x[23] = (N20596 & N20746) | (N20748 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N709);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17141 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[6] | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7494 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N708 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7494 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44986 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N707 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44986 | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N493 = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N708 ^ DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N707;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[31] = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17141) | (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N493)) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8]) | DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45115 = !((DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725 & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45148 = !(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45115 & (!DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991));
assign x[15] = !((N23918 & N23924) | ((!N23918) & DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45148));
reg x_reg_28__I4378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I4378_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[29];
	end
assign x[28] = x_reg_28__I4378_QOUT;
reg x_reg_30__I4380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I4380_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[30];
	end
assign x[30] = x_reg_30__I4380_QOUT;
reg x_reg_31__I4381_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I4381_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[31];
	end
assign x[31] = x_reg_31__I4381_QOUT;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[0] = x[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[1] = x[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[2] = x[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[3] = x[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[4] = x[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[5] = x[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[6] = x[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[7] = x[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[8] = x[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[9] = x[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[10] = x[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[11] = x[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[12] = x[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[13] = x[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[14] = x[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[15] = x[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[16] = x[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[17] = x[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[18] = x[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[19] = x[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[20] = x[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[21] = x[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[22] = x[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[23] = x[23];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[24] = x[24];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[25] = x[25];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[26] = x[26];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[27] = x[27];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[28] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[18] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[48] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[30] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[1] = 1'B0;
assign x[29] = x[28];
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urT3TA7ZrhpN : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



