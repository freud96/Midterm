/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:23:42 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42;
wire [22:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82;
wire [0:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195;
wire [32:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N682,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N684,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N688,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N696,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N698,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N734,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N735,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N739,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N740,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N743,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N746,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N747,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N751,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N753,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N754,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4079,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4113,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4134,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4141,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4162,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4166,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4168,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4176,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4190,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4204,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4205,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4210,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4224,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4233,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4238,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4262,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4283,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4289,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4303,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4312,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4314,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4319,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4320,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4326,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4330,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4331,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4338,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4342,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4350,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4363,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4366,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4369,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4396,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4403,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4412,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4422,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4425,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4438,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4461,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4469,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4471,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4482,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4483,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4489,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4559,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4585,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4590,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4607,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4632,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5388,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5433,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5462,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5489,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5500,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5837,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5839,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5852,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5854,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5857,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5867,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5871,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5879,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5892,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5893,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5900,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5908,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5913,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5964,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5979,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5980,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6063,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6079,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6141,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6166,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6168,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6186,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6199,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6223,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6242,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6248,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6260,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6289,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6304,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6309,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6311,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6315,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6319,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6323,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6325,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6327,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6331,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6340,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6342,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6350,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6353,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6357,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6358,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6361,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6396,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6419,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6433,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6438,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6444,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6452,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6458,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6471,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6474,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6482,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6483,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6500,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6514,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6535,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6572,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6585,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6599,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6603,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6625,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6646,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6647,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6671,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7561,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7599,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7642,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7644,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7652,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7674,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7675,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7684,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7698,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7702,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7703,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7705,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7706,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7709,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7710,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7713,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7714,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7715,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7718,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7721,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7723,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7724,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7725,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7727,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7728,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7729,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7730,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7731,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7732,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7743,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7747,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7751,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7754,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7760,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7761,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7762,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7764,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7765,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7766,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7767,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7768,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7769,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7770,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7771,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7772,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7773,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7774,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7779,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7780,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7782,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7783,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7785,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7788,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7791,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7792,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7793,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7794,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7795,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7796,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7797,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7798,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7801,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7803,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7804,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7806,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7807,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7809,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7811,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7813,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7815,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7816,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7817,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7819,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7821,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7822,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7824,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7826,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7828,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7829,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7830,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7833,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7834,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7836,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7855,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7864,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7867,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7871,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7885,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7889,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7891,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7892,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7896,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7900,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7949,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8652,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8656,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8671,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8675,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8688,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8696,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8702,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8705,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8708,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8709,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8710,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8711,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8713,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8714,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8715,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8717,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8718,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8719,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8720,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8721,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8723,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8725,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8726,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8727,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8728,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8729,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8731,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8732,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8735,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8740,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8743,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8746,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8756,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8758,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8760,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8761,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8762,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8763,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8764,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8765,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8767,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8768,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8769,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8771,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8773,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8774,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8776,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8777,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8780,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8783,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8784,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8785,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8787,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8789,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8791,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8792,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8793,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8795,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8796,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8797,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8798,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8801,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8802,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8803,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8804,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8806,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8810,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8813,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8814,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8815,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8816,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8819,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8820,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8821,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8823,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8826,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8827,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8828,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8830,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8833,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8835,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8836,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8839,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8841,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8844,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8852,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8855,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8857,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8867,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8879,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8880,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8892,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8893,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8896,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8904,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8980,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9105,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9113,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9134,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9136,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9147,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9162,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9163,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9176,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9179,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9186,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9195,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9205,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9210,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9223,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9224,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9238,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9260,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9309,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9311,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9312,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9315,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9319,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9326,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9330,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9333,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9337,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9338,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9340,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9363,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9366,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9396,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9403,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9419,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9431,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9433,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9438,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9444,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9458,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9462,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9469,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9482,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9489,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9514,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9572,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9581,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9585,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9593,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9603,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9607,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9625,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9642,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9644,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9647,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9653,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9671,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9674,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9702,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9703,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9705,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9709,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9710,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9711,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9714,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9716,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9718,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9719,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9722,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9725,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9726,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9727,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9729,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9730,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9731,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9732,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9734,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9735,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9739,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9740,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9746,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9753,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9758,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9760,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9761,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9762,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9763,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9764,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9765,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9766,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9767,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9769,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9771,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9773,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9774,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9776,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9779,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9781,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9784,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9787,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9789,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9791,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9792,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9793,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9794,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9796,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9797,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9798,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9799,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9802,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9805,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9807,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9811,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9814,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9815,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9816,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9820,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9821,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9823,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9824,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9826,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9827,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9828,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9829,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9831,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9833,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9835,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9836,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9844,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9852,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9856,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9864,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9879,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9885,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9889,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9891,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9893,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9896,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9904,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9913,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9949,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9964,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9979,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9980,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10079,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10091,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10100,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10105,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10122,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10134,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10159,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10163,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10179,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10186,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10190,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10195,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10199,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10223,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10224,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10256,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10262,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10264,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10286,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10290,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10303,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10304,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12100,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12163,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12179,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12210,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12260,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12264,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12320,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12350,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12384,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12444,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12466,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13332,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13337,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13340,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13358,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13384,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13388,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13398,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13475,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37720;
wire N9100,N18660,N18664,N18667,N18678,N18835,N18839 
	,N18879,N18881,N18886,N18971,N18990,N19000,N19010,N19020 
	,N19030,N19040,N19050,N19060,N19070,N19080,N19099,N19109 
	,N19119,N19129,N19139,N19149,N19159,N19223,N19233,N19275 
	,N19410,N19633,N19768,N19891,N19900,N19909,N20144,N20175 
	,N20182,N20492,N20538,N20660,N21070,N21075,N21080,N21085 
	,N21090,N21100,N21105,N21765,N21769,N21782,N21795,N21988 
	,N21993,N21999,N22003,N22305,N22309,N22618,N22929,N22939 
	,N22949,N22959,N22969,N22979,N22989,N23008,N23018,N23035 
	,N23050,N23060,N23070,N23080,N23090,N23100,N23110,N23120 
	,N23130,N23140,N23142,N23333,N23335,N23378,N23556,N23579 
	,N23859,N23861,N23943,N23945,N24239,N24241,N24248,N24250 
	,N24268,N24432,N24633,N24635,N24642,N24644,N24653,N24662 
	,N25288,N25295,N25297,N25313,N25457,N25627,N25766,N25768 
	,N25852,N25854,N26198,N26206,N26208,N26228,N26230,N26236 
	,N26238,N26244,N26246,N26248,N26252,N26254,N26256,N26646 
	,N26654,N26704,N26726,N26734,N26736,N26742,N26744,N26750 
	,N26752,N26758,N26760,N26766,N26768,N27092,N27094,N27100 
	,N27102,N27231,N27448,N27456,N27640,N27844,N27939,N28088 
	,N28113,N28287,N28313,N29392,N29396,N29398,N29426,N29430 
	,N29442,N29446,N29448,N29450,N29452,N29454,N29456,N29458 
	,N29460,N29462,N29464,N29466,N29468,N29470,N29472,N29474 
	,N29476,N29478,N29480,N29482,N29484,N29486,N29488,N29490 
	,N29492,N29494,N29496,N29498,N29502,N29506,N29510,N29556 
	,N29560,N29566,N29570,N29580,N29592,N29598,N29610,N29612 
	,N29614,N29616,N29618,N29620,N29622,N29624,N29626,N29653 
	,N29655,N29667,N29669,N29673,N29679,N29681,N30223,N30224 
	,N30225,N30226,N30227,N30228,N30229,N30230,N30231,N30232 
	,N30233,N30234,N30235,N30236,N30237,N30238,N30239,N30240 
	,N30241,N30242,N30243,N30244,N30245,N30246,N30247,N30248 
	,N30249,N30250,N30251,N30252,N30253,N30254,N30255,N30256 
	,N30257,N30258,N30259,N30260,N30261,N30262,N30263,N30264 
	,N30265,N30266,N30267,N30268,N30269,N30270,N30271,N30272 
	,N30273,N30274,N30275,N30276,N30277,N30278,N30279,N30280 
	,N30281,N30282,N30283,N30284,N30285,N30286,N30287,N30288 
	,N30289,N30290,N30291,N30292,N30293,N30294,N30295,N30296 
	,N30297,N30298,N30299,N30300,N30301,N30302,N30303,N30304 
	,N30305,N30306,N30307,N30308,N30309,N30310,N30311,N30312 
	,N30313,N30315,N30316,N30323,N30329,N30336,N30343,N30352 
	,N30360,N30368,N30373;
reg x_reg_L0_31__retimed_I15390_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15390_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002;
	end
assign N29681 = x_reg_L0_31__retimed_I15390_QOUT;
reg x_reg_L0_31__retimed_I15389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15389_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921;
	end
assign N29679 = x_reg_L0_31__retimed_I15389_QOUT;
reg x_reg_L0_31__retimed_I15387_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15387_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330;
	end
assign N29673 = x_reg_L0_31__retimed_I15387_QOUT;
reg x_reg_L0_31__retimed_I15386_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15386_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355;
	end
assign N29669 = x_reg_L0_31__retimed_I15386_QOUT;
reg x_reg_L0_31__retimed_I15385_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15385_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276;
	end
assign N29667 = x_reg_L0_31__retimed_I15385_QOUT;
reg x_reg_L0_31__retimed_I15380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15380_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10109;
	end
assign N29655 = x_reg_L0_31__retimed_I15380_QOUT;
reg x_reg_L0_31__retimed_I15379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15379_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9746;
	end
assign N29653 = x_reg_L0_31__retimed_I15379_QOUT;
reg x_reg_L0_31__retimed_I15368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15368_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9486;
	end
assign N29626 = x_reg_L0_31__retimed_I15368_QOUT;
reg x_reg_L0_31__retimed_I15367_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15367_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9098;
	end
assign N29624 = x_reg_L0_31__retimed_I15367_QOUT;
reg x_reg_L0_31__retimed_I15366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15366_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8668;
	end
assign N29622 = x_reg_L0_31__retimed_I15366_QOUT;
reg x_reg_L0_31__retimed_I15365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15365_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9982;
	end
assign N29620 = x_reg_L0_31__retimed_I15365_QOUT;
reg x_reg_L0_31__retimed_I15364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15364_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9147;
	end
assign N29618 = x_reg_L0_31__retimed_I15364_QOUT;
reg x_reg_L0_31__retimed_I15363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15363_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8791;
	end
assign N29616 = x_reg_L0_31__retimed_I15363_QOUT;
reg x_reg_L0_31__retimed_I15362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15362_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[32];
	end
assign N29614 = x_reg_L0_31__retimed_I15362_QOUT;
reg x_reg_L0_31__retimed_I15361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15361_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9601;
	end
assign N29612 = x_reg_L0_31__retimed_I15361_QOUT;
reg x_reg_L0_31__retimed_I15360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15360_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9212;
	end
assign N29610 = x_reg_L0_31__retimed_I15360_QOUT;
reg x_reg_L0_31__retimed_I15354_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15354_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[31];
	end
assign N29598 = x_reg_L0_31__retimed_I15354_QOUT;
reg x_reg_L0_31__retimed_I15351_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15351_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[30];
	end
assign N29592 = x_reg_L0_31__retimed_I15351_QOUT;
reg x_reg_L0_31__retimed_I15345_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15345_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[29];
	end
assign N29580 = x_reg_L0_31__retimed_I15345_QOUT;
reg x_reg_L0_31__retimed_I15340_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15340_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[27];
	end
assign N29570 = x_reg_L0_31__retimed_I15340_QOUT;
reg x_reg_L0_31__retimed_I15338_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15338_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11918;
	end
assign N29566 = x_reg_L0_31__retimed_I15338_QOUT;
reg x_reg_L0_31__retimed_I15335_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15335_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[26];
	end
assign N29560 = x_reg_L0_31__retimed_I15335_QOUT;
reg x_reg_L0_31__retimed_I15333_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15333_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9153;
	end
assign N29556 = x_reg_L0_31__retimed_I15333_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15636 (.Y(N30223), .A(N29556));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15637 (.Y(N30224), .A(N30223));
reg x_reg_L0_31__retimed_I15310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15310_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12415;
	end
assign N29510 = x_reg_L0_31__retimed_I15310_QOUT;
reg x_reg_L0_31__retimed_I15308_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15308_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12222;
	end
assign N29506 = x_reg_L0_31__retimed_I15308_QOUT;
reg x_reg_L0_31__retimed_I15306_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15306_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12080;
	end
assign N29502 = x_reg_L0_31__retimed_I15306_QOUT;
reg x_reg_L0_31__retimed_I15304_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15304_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9890;
	end
assign N29498 = x_reg_L0_31__retimed_I15304_QOUT;
reg x_reg_L0_31__retimed_I15303_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15303_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9089;
	end
assign N29496 = x_reg_L0_31__retimed_I15303_QOUT;
reg x_reg_L0_31__retimed_I15302_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15302_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8744;
	end
assign N29494 = x_reg_L0_31__retimed_I15302_QOUT;
reg x_reg_L0_31__retimed_I15301_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15301_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9983;
	end
assign N29492 = x_reg_L0_31__retimed_I15301_QOUT;
reg x_reg_L0_31__retimed_I15300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15300_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9611;
	end
assign N29490 = x_reg_L0_31__retimed_I15300_QOUT;
reg x_reg_L0_31__retimed_I15299_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15299_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9072;
	end
assign N29488 = x_reg_L0_31__retimed_I15299_QOUT;
reg x_reg_L0_31__retimed_I15298_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15298_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8731;
	end
assign N29486 = x_reg_L0_31__retimed_I15298_QOUT;
reg x_reg_L0_31__retimed_I15297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15297_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9860;
	end
assign N29484 = x_reg_L0_31__retimed_I15297_QOUT;
reg x_reg_L0_31__retimed_I15296_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15296_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9469;
	end
assign N29482 = x_reg_L0_31__retimed_I15296_QOUT;
reg x_reg_L0_31__retimed_I15295_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15295_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9237;
	end
assign N29480 = x_reg_L0_31__retimed_I15295_QOUT;
reg x_reg_L0_31__retimed_I15294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15294_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8866;
	end
assign N29478 = x_reg_L0_31__retimed_I15294_QOUT;
reg x_reg_L0_31__retimed_I15293_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15293_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9120;
	end
assign N29476 = x_reg_L0_31__retimed_I15293_QOUT;
reg x_reg_L0_31__retimed_I15292_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15292_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8771;
	end
assign N29474 = x_reg_L0_31__retimed_I15292_QOUT;
reg x_reg_L0_31__retimed_I15291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15291_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9417;
	end
assign N29472 = x_reg_L0_31__retimed_I15291_QOUT;
reg x_reg_L0_31__retimed_I15290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15290_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9035;
	end
assign N29470 = x_reg_L0_31__retimed_I15290_QOUT;
reg x_reg_L0_31__retimed_I15289_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15289_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10167;
	end
assign N29468 = x_reg_L0_31__retimed_I15289_QOUT;
reg x_reg_L0_31__retimed_I15288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15288_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9807;
	end
assign N29466 = x_reg_L0_31__retimed_I15288_QOUT;
reg x_reg_L0_31__retimed_I15287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15287_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10202;
	end
assign N29464 = x_reg_L0_31__retimed_I15287_QOUT;
reg x_reg_L0_31__retimed_I15286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15286_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9846;
	end
assign N29462 = x_reg_L0_31__retimed_I15286_QOUT;
reg x_reg_L0_31__retimed_I15285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15285_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9497;
	end
assign N29460 = x_reg_L0_31__retimed_I15285_QOUT;
reg x_reg_L0_31__retimed_I15284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15284_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9105;
	end
assign N29458 = x_reg_L0_31__retimed_I15284_QOUT;
reg x_reg_L0_31__retimed_I15283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15283_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9156;
	end
assign N29456 = x_reg_L0_31__retimed_I15283_QOUT;
reg x_reg_L0_31__retimed_I15282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15282_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8798;
	end
assign N29454 = x_reg_L0_31__retimed_I15282_QOUT;
reg x_reg_L0_31__retimed_I15281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15281_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8789;
	end
assign N29452 = x_reg_L0_31__retimed_I15281_QOUT;
reg x_reg_L0_31__retimed_I15280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15280_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10124;
	end
assign N29450 = x_reg_L0_31__retimed_I15280_QOUT;
reg x_reg_L0_31__retimed_I15279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15279_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9811;
	end
assign N29448 = x_reg_L0_31__retimed_I15279_QOUT;
reg x_reg_L0_31__retimed_I15278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15278_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9426;
	end
assign N29446 = x_reg_L0_31__retimed_I15278_QOUT;
reg x_reg_L0_31__retimed_I15276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15276_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[24];
	end
assign N29442 = x_reg_L0_31__retimed_I15276_QOUT;
reg x_reg_L0_31__retimed_I15270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15270_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[25];
	end
assign N29430 = x_reg_L0_31__retimed_I15270_QOUT;
reg x_reg_L0_31__retimed_I15268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15268_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[28];
	end
assign N29426 = x_reg_L0_31__retimed_I15268_QOUT;
reg x_reg_L0_31__retimed_I15255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15255_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9397;
	end
assign N29398 = x_reg_L0_31__retimed_I15255_QOUT;
reg x_reg_L0_31__retimed_I15254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15254_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9015;
	end
assign N29396 = x_reg_L0_31__retimed_I15254_QOUT;
reg x_reg_L0_31__retimed_I15252_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15252_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[22];
	end
assign N29392 = x_reg_L0_31__retimed_I15252_QOUT;
reg x_reg_L0_31__retimed_I14964_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14964_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[18];
	end
assign N28313 = x_reg_L0_31__retimed_I14964_QOUT;
reg x_reg_L0_31__retimed_I14962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14962_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[20];
	end
assign N28287 = x_reg_L0_31__retimed_I14962_QOUT;
reg x_reg_L0_31__retimed_I14921_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14921_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[19];
	end
assign N28113 = x_reg_L0_31__retimed_I14921_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15638 (.Y(N30225), .A(N28113));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15639 (.Y(N30226), .A(N30225));
reg x_reg_L0_31__retimed_I14912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14912_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[21];
	end
assign N28088 = x_reg_L0_31__retimed_I14912_QOUT;
reg x_reg_L0_31__retimed_I14868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14868_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[23];
	end
assign N27939 = x_reg_L0_31__retimed_I14868_QOUT;
reg x_reg_L0_31__retimed_I14846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14846_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9564;
	end
assign N27844 = x_reg_L0_31__retimed_I14846_QOUT;
reg x_reg_L0_31__retimed_I14791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14791_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9476;
	end
assign N27640 = x_reg_L0_31__retimed_I14791_QOUT;
reg x_reg_L0_31__retimed_I14734_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14734_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9344;
	end
assign N27456 = x_reg_L0_31__retimed_I14734_QOUT;
reg x_reg_L0_31__retimed_I14731_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14731_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9030;
	end
assign N27448 = x_reg_L0_31__retimed_I14731_QOUT;
reg x_reg_L0_31__retimed_I14653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14653_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8717;
	end
assign N27231 = x_reg_L0_31__retimed_I14653_QOUT;
reg x_reg_L0_31__retimed_I14604_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14604_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8857;
	end
assign N27102 = x_reg_L0_31__retimed_I14604_QOUT;
reg x_reg_L0_31__retimed_I14603_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14603_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9840;
	end
assign N27100 = x_reg_L0_31__retimed_I14603_QOUT;
reg x_reg_L0_31__retimed_I14601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14601_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8872;
	end
assign N27094 = x_reg_L0_31__retimed_I14601_QOUT;
reg x_reg_L0_31__retimed_I14600_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14600_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10127;
	end
assign N27092 = x_reg_L0_31__retimed_I14600_QOUT;
reg x_reg_L0_31__retimed_I14504_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14504_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9039;
	end
assign N26768 = x_reg_L0_31__retimed_I14504_QOUT;
reg x_reg_L0_31__retimed_I14503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14503_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10021;
	end
assign N26766 = x_reg_L0_31__retimed_I14503_QOUT;
reg x_reg_L0_31__retimed_I14501_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14501_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9739;
	end
assign N26760 = x_reg_L0_31__retimed_I14501_QOUT;
reg x_reg_L0_31__retimed_I14500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14500_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10134;
	end
assign N26758 = x_reg_L0_31__retimed_I14500_QOUT;
reg x_reg_L0_31__retimed_I14498_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14498_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9073;
	end
assign N26752 = x_reg_L0_31__retimed_I14498_QOUT;
reg x_reg_L0_31__retimed_I14497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14497_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8758;
	end
assign N26750 = x_reg_L0_31__retimed_I14497_QOUT;
reg x_reg_L0_31__retimed_I14495_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14495_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9364;
	end
assign N26744 = x_reg_L0_31__retimed_I14495_QOUT;
reg x_reg_L0_31__retimed_I14494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14494_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9108;
	end
assign N26742 = x_reg_L0_31__retimed_I14494_QOUT;
reg x_reg_L0_31__retimed_I14492_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14492_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8760;
	end
assign N26736 = x_reg_L0_31__retimed_I14492_QOUT;
reg x_reg_L0_31__retimed_I14491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14491_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9243;
	end
assign N26734 = x_reg_L0_31__retimed_I14491_QOUT;
reg x_reg_L0_31__retimed_I14488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14488_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9757;
	end
assign N26726 = x_reg_L0_31__retimed_I14488_QOUT;
reg x_reg_L0_31__retimed_I14479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14479_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10092;
	end
assign N26704 = x_reg_L0_31__retimed_I14479_QOUT;
reg x_reg_L0_31__retimed_I14458_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14458_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9773;
	end
assign N26654 = x_reg_L0_31__retimed_I14458_QOUT;
reg x_reg_L0_31__retimed_I14455_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14455_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9227;
	end
assign N26646 = x_reg_L0_31__retimed_I14455_QOUT;
reg x_reg_L0_31__retimed_I14320_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14320_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10156;
	end
assign N26256 = x_reg_L0_31__retimed_I14320_QOUT;
reg x_reg_L0_31__retimed_I14319_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14319_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9408;
	end
assign N26254 = x_reg_L0_31__retimed_I14319_QOUT;
reg x_reg_L0_31__retimed_I14318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14318_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9607;
	end
assign N26252 = x_reg_L0_31__retimed_I14318_QOUT;
reg x_reg_L0_31__retimed_I14317_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14317_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10026;
	end
assign N26248 = x_reg_L0_31__retimed_I14317_QOUT;
reg x_reg_L0_31__retimed_I14316_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14316_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9265;
	end
assign N26246 = x_reg_L0_31__retimed_I14316_QOUT;
reg x_reg_L0_31__retimed_I14315_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14315_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10208;
	end
assign N26244 = x_reg_L0_31__retimed_I14315_QOUT;
reg x_reg_L0_31__retimed_I14313_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14313_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8903;
	end
assign N26238 = x_reg_L0_31__retimed_I14313_QOUT;
reg x_reg_L0_31__retimed_I14312_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14312_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9085;
	end
assign N26236 = x_reg_L0_31__retimed_I14312_QOUT;
reg x_reg_L0_31__retimed_I14310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14310_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8816;
	end
assign N26230 = x_reg_L0_31__retimed_I14310_QOUT;
reg x_reg_L0_31__retimed_I14309_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14309_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9370;
	end
assign N26228 = x_reg_L0_31__retimed_I14309_QOUT;
reg x_reg_L0_31__retimed_I14301_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14301_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10035;
	end
assign N26208 = x_reg_L0_31__retimed_I14301_QOUT;
reg x_reg_L0_31__retimed_I14300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14300_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9852;
	end
assign N26206 = x_reg_L0_31__retimed_I14300_QOUT;
reg x_reg_L0_31__retimed_I14297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14297_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8742;
	end
assign N26198 = x_reg_L0_31__retimed_I14297_QOUT;
reg x_reg_L0_31__retimed_I14154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14154_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10310;
	end
assign N25854 = x_reg_L0_31__retimed_I14154_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15640 (.Y(N30227), .A(N25854));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15641 (.Y(N30228), .A(N30227));
reg x_reg_L0_31__retimed_I14153_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14153_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8975;
	end
assign N25852 = x_reg_L0_31__retimed_I14153_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15642 (.Y(N30229), .A(N25852));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15643 (.Y(N30230), .A(N30229));
reg x_reg_L0_31__retimed_I14121_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14121_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8710;
	end
assign N25768 = x_reg_L0_31__retimed_I14121_QOUT;
reg x_reg_L0_31__retimed_I14120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14120_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9687;
	end
assign N25766 = x_reg_L0_31__retimed_I14120_QOUT;
reg x_reg_L0_31__retimed_I14062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14062_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9666;
	end
assign N25627 = x_reg_L0_31__retimed_I14062_QOUT;
reg x_reg_L0_31__retimed_I13990_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13990_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9219;
	end
assign N25457 = x_reg_L0_31__retimed_I13990_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15644 (.Y(N30231), .A(N25457));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15645 (.Y(N30232), .A(N30231));
reg x_reg_L0_31__retimed_I13930_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13930_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10108;
	end
assign N25313 = x_reg_L0_31__retimed_I13930_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15646 (.Y(N30233), .A(N25313));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15647 (.Y(N30234), .A(N30233));
reg x_reg_L0_31__retimed_I13923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13923_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9352;
	end
assign N25297 = x_reg_L0_31__retimed_I13923_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15648 (.Y(N30235), .A(N25297));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15649 (.Y(N30236), .A(N30235));
reg x_reg_L0_31__retimed_I13922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13922_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9745;
	end
assign N25295 = x_reg_L0_31__retimed_I13922_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15650 (.Y(N30237), .A(N25295));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15651 (.Y(N30238), .A(N30237));
reg x_reg_L0_31__retimed_I13919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13919_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8774;
	end
assign N25288 = x_reg_L0_31__retimed_I13919_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15652 (.Y(N30239), .A(N25288));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15653 (.Y(N30240), .A(N30239));
reg x_reg_L0_31__retimed_I13661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13661_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9894;
	end
assign N24662 = x_reg_L0_31__retimed_I13661_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15654 (.Y(N30241), .A(N24662));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15655 (.Y(N30242), .A(N30241));
reg x_reg_L0_31__retimed_I13657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13657_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9284;
	end
assign N24653 = x_reg_L0_31__retimed_I13657_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15656 (.Y(N30243), .A(N24653));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15657 (.Y(N30244), .A(N30243));
reg x_reg_L0_31__retimed_I13653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13653_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9125;
	end
assign N24644 = x_reg_L0_31__retimed_I13653_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15658 (.Y(N30245), .A(N24644));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15659 (.Y(N30246), .A(N30245));
reg x_reg_L0_31__retimed_I13652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13652_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9517;
	end
assign N24642 = x_reg_L0_31__retimed_I13652_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15660 (.Y(N30247), .A(N24642));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15661 (.Y(N30248), .A(N30247));
reg x_reg_L0_31__retimed_I13649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13649_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10255;
	end
assign N24635 = x_reg_L0_31__retimed_I13649_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15662 (.Y(N30249), .A(N24635));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15663 (.Y(N30250), .A(N30249));
reg x_reg_L0_31__retimed_I13648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13648_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8914;
	end
assign N24633 = x_reg_L0_31__retimed_I13648_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15664 (.Y(N30251), .A(N24633));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15665 (.Y(N30252), .A(N30251));
reg x_reg_L0_31__retimed_I13572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13572_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8852;
	end
assign N24432 = x_reg_L0_31__retimed_I13572_QOUT;
reg x_reg_L0_31__retimed_I13503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13503_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9677;
	end
assign N24268 = x_reg_L0_31__retimed_I13503_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15666 (.Y(N30253), .A(N24268));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15667 (.Y(N30254), .A(N30253));
reg x_reg_L0_31__retimed_I13495_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13495_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10044;
	end
assign N24250 = x_reg_L0_31__retimed_I13495_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15668 (.Y(N30255), .A(N24250));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15669 (.Y(N30256), .A(N30255));
reg x_reg_L0_31__retimed_I13494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13494_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6236;
	end
assign N24248 = x_reg_L0_31__retimed_I13494_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15670 (.Y(N30257), .A(N24248));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15671 (.Y(N30258), .A(N30257));
reg x_reg_L0_31__retimed_I13491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13491_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9064;
	end
assign N24241 = x_reg_L0_31__retimed_I13491_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15672 (.Y(N30259), .A(N24241));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15673 (.Y(N30260), .A(N30259));
reg x_reg_L0_31__retimed_I13490_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13490_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9447;
	end
assign N24239 = x_reg_L0_31__retimed_I13490_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15674 (.Y(N30261), .A(N24239));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15675 (.Y(N30262), .A(N30261));
reg x_reg_L0_31__retimed_I13379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13379_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8821;
	end
assign N23945 = x_reg_L0_31__retimed_I13379_QOUT;
reg x_reg_L0_31__retimed_I13378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13378_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10073;
	end
assign N23943 = x_reg_L0_31__retimed_I13378_QOUT;
reg x_reg_L0_31__retimed_I13344_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13344_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9832;
	end
assign N23861 = x_reg_L0_31__retimed_I13344_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15676 (.Y(N30263), .A(N23861));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15677 (.Y(N30264), .A(N30263));
reg x_reg_L0_31__retimed_I13343_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13343_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10191;
	end
assign N23859 = x_reg_L0_31__retimed_I13343_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15678 (.Y(N30265), .A(N23859));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15679 (.Y(N30266), .A(N30265));
reg x_reg_L0_31__retimed_I13240_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13240_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9181;
	end
assign N23579 = x_reg_L0_31__retimed_I13240_QOUT;
reg x_reg_L0_31__retimed_I13231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13231_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8851;
	end
assign N23556 = x_reg_L0_31__retimed_I13231_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15680 (.Y(N30267), .A(N23556));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15681 (.Y(N30268), .A(N30267));
reg x_reg_L0_31__retimed_I13163_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13163_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[0];
	end
assign N23378 = x_reg_L0_31__retimed_I13163_QOUT;
reg x_reg_L0_31__retimed_I13148_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13148_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9763;
	end
assign N23335 = x_reg_L0_31__retimed_I13148_QOUT;
reg x_reg_L0_31__retimed_I13147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13147_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8844;
	end
assign N23333 = x_reg_L0_31__retimed_I13147_QOUT;
reg x_reg_L0_31__retimed_I13074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13074_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[38];
	end
assign N23142 = x_reg_L0_31__retimed_I13074_QOUT;
reg x_reg_L0_31__retimed_I13073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13073_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[20];
	end
assign N23140 = x_reg_L0_31__retimed_I13073_QOUT;
reg x_reg_L0_31__retimed_I13070_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13070_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[19];
	end
assign N23130 = x_reg_L0_31__retimed_I13070_QOUT;
reg x_reg_L0_31__retimed_I13067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13067_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[18];
	end
assign N23120 = x_reg_L0_31__retimed_I13067_QOUT;
reg x_reg_L0_31__retimed_I13064_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13064_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[17];
	end
assign N23110 = x_reg_L0_31__retimed_I13064_QOUT;
reg x_reg_L0_31__retimed_I13061_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13061_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[16];
	end
assign N23100 = x_reg_L0_31__retimed_I13061_QOUT;
reg x_reg_L0_31__retimed_I13058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13058_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[15];
	end
assign N23090 = x_reg_L0_31__retimed_I13058_QOUT;
reg x_reg_L0_31__retimed_I13055_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13055_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[14];
	end
assign N23080 = x_reg_L0_31__retimed_I13055_QOUT;
reg x_reg_L0_31__retimed_I13052_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13052_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[13];
	end
assign N23070 = x_reg_L0_31__retimed_I13052_QOUT;
reg x_reg_L0_31__retimed_I13049_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13049_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[12];
	end
assign N23060 = x_reg_L0_31__retimed_I13049_QOUT;
reg x_reg_L0_31__retimed_I13046_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13046_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[11];
	end
assign N23050 = x_reg_L0_31__retimed_I13046_QOUT;
reg x_reg_L0_31__retimed_I13041_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13041_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[8];
	end
assign N23035 = x_reg_L0_31__retimed_I13041_QOUT;
reg x_reg_L0_31__retimed_I13035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13035_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[5];
	end
assign N23018 = x_reg_L0_31__retimed_I13035_QOUT;
reg x_reg_L0_31__retimed_I13032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13032_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[10];
	end
assign N23008 = x_reg_L0_31__retimed_I13032_QOUT;
reg x_reg_L0_31__retimed_I13025_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13025_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[4];
	end
assign N22989 = x_reg_L0_31__retimed_I13025_QOUT;
reg x_reg_L0_31__retimed_I13022_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13022_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[1];
	end
assign N22979 = x_reg_L0_31__retimed_I13022_QOUT;
reg x_reg_L0_31__retimed_I13019_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13019_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[2];
	end
assign N22969 = x_reg_L0_31__retimed_I13019_QOUT;
reg x_reg_L0_31__retimed_I13016_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13016_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[3];
	end
assign N22959 = x_reg_L0_31__retimed_I13016_QOUT;
reg x_reg_L0_31__retimed_I13013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13013_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[9];
	end
assign N22949 = x_reg_L0_31__retimed_I13013_QOUT;
reg x_reg_L0_31__retimed_I13010_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13010_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[7];
	end
assign N22939 = x_reg_L0_31__retimed_I13010_QOUT;
reg x_reg_L0_31__retimed_I13007_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13007_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[6];
	end
assign N22929 = x_reg_L0_31__retimed_I13007_QOUT;
reg x_reg_L0_31__retimed_I12919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12919_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12365;
	end
assign N22618 = x_reg_L0_31__retimed_I12919_QOUT;
reg x_reg_L0_31__retimed_I12818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12818_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102;
	end
assign N22309 = x_reg_L0_31__retimed_I12818_QOUT;
reg x_reg_L0_31__retimed_I12816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12816_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240;
	end
assign N22305 = x_reg_L0_31__retimed_I12816_QOUT;
reg x_reg_L0_31__retimed_I12715_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12715_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944;
	end
assign N22003 = x_reg_L0_31__retimed_I12715_QOUT;
reg x_reg_L0_31__retimed_I12713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12713_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075;
	end
assign N21999 = x_reg_L0_31__retimed_I12713_QOUT;
reg x_reg_L0_31__retimed_I12711_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12711_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437;
	end
assign N21993 = x_reg_L0_31__retimed_I12711_QOUT;
reg x_reg_L0_31__retimed_I12710_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12710_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298;
	end
assign N21988 = x_reg_L0_31__retimed_I12710_QOUT;
reg x_reg_L0_31__retimed_I12644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12644_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12246;
	end
assign N21795 = x_reg_L0_31__retimed_I12644_QOUT;
reg x_reg_L0_31__retimed_I12639_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12639_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12328;
	end
assign N21782 = x_reg_L0_31__retimed_I12639_QOUT;
reg x_reg_L0_31__retimed_I12634_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12634_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12055;
	end
assign N21769 = x_reg_L0_31__retimed_I12634_QOUT;
reg x_reg_L0_31__retimed_I12632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12632_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12188;
	end
assign N21765 = x_reg_L0_31__retimed_I12632_QOUT;
reg x_reg_L0_31__retimed_I12380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12380_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11950;
	end
assign N21105 = x_reg_L0_31__retimed_I12380_QOUT;
reg x_reg_L0_31__retimed_I12378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12378_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12362;
	end
assign N21100 = x_reg_L0_31__retimed_I12378_QOUT;
reg x_reg_L0_31__retimed_I12374_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12374_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12115;
	end
assign N21090 = x_reg_L0_31__retimed_I12374_QOUT;
reg x_reg_L0_31__retimed_I12372_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12372_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11927;
	end
assign N21085 = x_reg_L0_31__retimed_I12372_QOUT;
reg x_reg_L0_31__retimed_I12370_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12370_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12335;
	end
assign N21080 = x_reg_L0_31__retimed_I12370_QOUT;
reg x_reg_L0_31__retimed_I12368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12368_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11901;
	end
assign N21075 = x_reg_L0_31__retimed_I12368_QOUT;
reg x_reg_L0_31__retimed_I12366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12366_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12138;
	end
assign N21070 = x_reg_L0_31__retimed_I12366_QOUT;
reg x_reg_L0_31__retimed_I12237_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12237_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11976;
	end
assign N20660 = x_reg_L0_31__retimed_I12237_QOUT;
reg x_reg_L0_31__retimed_I12190_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12190_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400;
	end
assign N20538 = x_reg_L0_31__retimed_I12190_QOUT;
reg x_reg_L0_31__retimed_I12181_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12181_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22];
	end
assign N20492 = x_reg_L0_31__retimed_I12181_QOUT;
reg x_reg_L0_31__retimed_I12116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12116_QOUT <= a_exp[5];
	end
assign N20182 = x_reg_L0_31__retimed_I12116_QOUT;
reg x_reg_L0_31__retimed_I12113_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12113_QOUT <= a_exp[6];
	end
assign N20175 = x_reg_L0_31__retimed_I12113_QOUT;
reg x_reg_L0_31__retimed_I12103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12103_QOUT <= a_exp[0];
	end
assign N20144 = x_reg_L0_31__retimed_I12103_QOUT;
reg x_reg_L0_31__retimed_I12021_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12021_QOUT <= a_exp[1];
	end
assign N19909 = x_reg_L0_31__retimed_I12021_QOUT;
reg x_reg_L0_31__retimed_I12017_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12017_QOUT <= a_exp[2];
	end
assign N19900 = x_reg_L0_31__retimed_I12017_QOUT;
reg x_reg_L0_31__retimed_I12013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12013_QOUT <= a_exp[4];
	end
assign N19891 = x_reg_L0_31__retimed_I12013_QOUT;
reg x_reg_L0_31__retimed_I11972_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11972_QOUT <= a_exp[3];
	end
assign N19768 = x_reg_L0_31__retimed_I11972_QOUT;
reg x_reg_L0_31__retimed_I11920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11920_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647;
	end
assign N19633 = x_reg_L0_31__retimed_I11920_QOUT;
reg x_reg_L0_31__retimed_I11828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11828_QOUT <= a_man[0];
	end
assign N19410 = x_reg_L0_31__retimed_I11828_QOUT;
reg x_reg_L0_31__retimed_I11770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11770_QOUT <= a_man[1];
	end
assign N19275 = x_reg_L0_31__retimed_I11770_QOUT;
reg x_reg_L0_31__retimed_I11753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11753_QOUT <= a_man[3];
	end
assign N19233 = x_reg_L0_31__retimed_I11753_QOUT;
reg x_reg_L0_31__retimed_I11749_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11749_QOUT <= a_man[2];
	end
assign N19223 = x_reg_L0_31__retimed_I11749_QOUT;
reg x_reg_L0_31__retimed_I11721_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11721_QOUT <= a_man[7];
	end
assign N19159 = x_reg_L0_31__retimed_I11721_QOUT;
reg x_reg_L0_31__retimed_I11717_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11717_QOUT <= a_man[10];
	end
assign N19149 = x_reg_L0_31__retimed_I11717_QOUT;
reg x_reg_L0_31__retimed_I11713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11713_QOUT <= a_man[6];
	end
assign N19139 = x_reg_L0_31__retimed_I11713_QOUT;
reg x_reg_L0_31__retimed_I11709_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11709_QOUT <= a_man[8];
	end
assign N19129 = x_reg_L0_31__retimed_I11709_QOUT;
reg x_reg_L0_31__retimed_I11705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11705_QOUT <= a_man[11];
	end
assign N19119 = x_reg_L0_31__retimed_I11705_QOUT;
reg x_reg_L0_31__retimed_I11701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11701_QOUT <= a_man[12];
	end
assign N19109 = x_reg_L0_31__retimed_I11701_QOUT;
reg x_reg_L0_31__retimed_I11697_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11697_QOUT <= a_man[13];
	end
assign N19099 = x_reg_L0_31__retimed_I11697_QOUT;
reg x_reg_L0_31__retimed_I11689_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11689_QOUT <= N30313;
	end
assign N19080 = x_reg_L0_31__retimed_I11689_QOUT;
reg x_reg_L0_31__retimed_I11685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11685_QOUT <= a_man[5];
	end
assign N19070 = x_reg_L0_31__retimed_I11685_QOUT;
reg x_reg_L0_31__retimed_I11681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11681_QOUT <= a_man[9];
	end
assign N19060 = x_reg_L0_31__retimed_I11681_QOUT;
reg x_reg_L0_31__retimed_I11677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11677_QOUT <= a_man[14];
	end
assign N19050 = x_reg_L0_31__retimed_I11677_QOUT;
reg x_reg_L0_31__retimed_I11673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11673_QOUT <= a_man[15];
	end
assign N19040 = x_reg_L0_31__retimed_I11673_QOUT;
reg x_reg_L0_31__retimed_I11669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11669_QOUT <= a_man[18];
	end
assign N19030 = x_reg_L0_31__retimed_I11669_QOUT;
reg x_reg_L0_31__retimed_I11665_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11665_QOUT <= a_man[20];
	end
assign N19020 = x_reg_L0_31__retimed_I11665_QOUT;
reg x_reg_L0_31__retimed_I11661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11661_QOUT <= a_man[17];
	end
assign N19010 = x_reg_L0_31__retimed_I11661_QOUT;
reg x_reg_L0_31__retimed_I11657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11657_QOUT <= a_man[19];
	end
assign N19000 = x_reg_L0_31__retimed_I11657_QOUT;
reg x_reg_L0_31__retimed_I11653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11653_QOUT <= a_man[16];
	end
assign N18990 = x_reg_L0_31__retimed_I11653_QOUT;
reg x_reg_L0_31__retimed_I11645_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11645_QOUT <= a_man[21];
	end
assign N18971 = x_reg_L0_31__retimed_I11645_QOUT;
reg x_reg_L0_22__retimed_I11608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I11608_QOUT <= a_man[22];
	end
assign N18886 = x_reg_L0_22__retimed_I11608_QOUT;
reg x_reg_L0_31__retimed_I11606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11606_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N577;
	end
assign N18881 = x_reg_L0_31__retimed_I11606_QOUT;
reg x_reg_L0_31__retimed_I11605_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11605_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487;
	end
assign N18879 = x_reg_L0_31__retimed_I11605_QOUT;
reg x_reg_L0_23__retimed_I11588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I11588_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580;
	end
assign N18839 = x_reg_L0_23__retimed_I11588_QOUT;
reg x_reg_L0_23__retimed_I11586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I11586_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026;
	end
assign N18835 = x_reg_L0_23__retimed_I11586_QOUT;
reg x_reg_L0_16__retimed_I11519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I11519_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82;
	end
assign N18678 = x_reg_L0_16__retimed_I11519_QOUT;
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15682 (.Y(N30269), .A(N18678));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15683 (.Y(N30270), .A(N30269));
reg x_reg_L0_21__retimed_I11514_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I11514_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759;
	end
assign N18667 = x_reg_L0_21__retimed_I11514_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15684 (.Y(N30271), .A(N18667));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15689 (.Y(N30276), .A(N30271));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15688 (.Y(N30275), .A(N30271));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15687 (.Y(N30274), .A(N30271));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15686 (.Y(N30273), .A(N30271));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15685 (.Y(N30272), .A(N30271));
reg x_reg_L0_31__retimed_I11513_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11513_QOUT <= a_sign;
	end
assign N18664 = x_reg_L0_31__retimed_I11513_QOUT;
reg x_reg_L0_31__retimed_I11511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11511_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639;
	end
assign N18660 = x_reg_L0_31__retimed_I11511_QOUT;
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15690 (.Y(N30277), .A(N18660));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15697 (.Y(N30284), .A(N30277));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15696 (.Y(N30283), .A(N30277));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15695 (.Y(N30282), .A(N30277));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15694 (.Y(N30281), .A(N30277));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15693 (.Y(N30280), .A(N30277));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15692 (.Y(N30279), .A(N30277));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15691 (.Y(N30278), .A(N30277));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13316), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[5]), .D(a_exp[6]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639), .A(a_exp[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13316));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360), .A(a_exp[3]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I4 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345), .A(a_exp[1]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I5 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345), .B(a_exp[2]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I6 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I7 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5347), .A(a_exp[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I8 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5347), .B(a_exp[5]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I9 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I10 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I11 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[1]), .B(a_exp[2]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I12 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I13 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[1]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I14 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A(a_exp[0]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .A(a_man[21]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I16 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .B(a_man[19]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I17 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4212), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4168), .A(a_man[15]), .B(a_man[17]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4489));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I18 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181), .A(a_man[22]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I19 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4153), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181), .B(a_man[20]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I20 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4528), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4374), .A(a_man[16]), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I21 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4212), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4153), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4374));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I22 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181), .B(a_man[20]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I23 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .A(a_man[20]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I24 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4113), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .B(a_man[18]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I25 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4554), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4064), .A(a_man[14]), .B(a_man[16]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4113));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I26 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3994), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4554), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4168));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I27 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I28 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I29 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .B(a_man[19]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I30 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958), .A(a_man[19]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I31 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958), .B(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I32 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4176), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3959), .A(a_man[13]), .B(a_man[15]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4449));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I33 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4331), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4176), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4064));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I34 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I35 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .B(a_man[18]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I36 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368), .A(a_man[18]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I37 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4387), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368), .B(a_man[16]), .CI(a_man[13]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I38 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4516), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4577), .A(a_man[12]), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4387));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I39 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3953), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4516), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3959));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I40 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I41 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I42 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958), .B(a_man[17]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I43 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052), .A(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I44 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4319), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4166), .A(a_man[10]), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I45 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4012), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4571), .A(a_man[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I46 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4141), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4471), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4319), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4012));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I47 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4294), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4141), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4577));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I48 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I49 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454), .A(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I50 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3943), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4109), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I51 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4075), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4600), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4571), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4166));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I52 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4229), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4075), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4471));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I53 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I54 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I55 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I56 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I57 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548), .A(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I58 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4560), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4403), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958), .B(a_man[21]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I59 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145), .A(a_man[15]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I60 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4215), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I61 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4438), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4342), .A(a_man[13]), .B(a_man[22]), .CI(a_man[10]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I62 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4283), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4130), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4560), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4215), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4342));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I63 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4411), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3989), .A(a_man[9]), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4283));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I64 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4378), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I65 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4504), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4348), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4378), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4438), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4109));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I66 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4504), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4600));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I67 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I68 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4307), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4360), .A(a_man[9]), .B(a_man[12]), .CI(a_man[7]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I69 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4297), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4144), .A(a_man[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I70 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4493), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4608), .A(a_man[6]), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4297));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I71 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4156), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4001), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4403), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4493), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4360));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I72 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4190), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4307), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4156));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I73 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4348), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4190), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3989));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I74 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I75 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I76 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236), .A(a_man[13]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I77 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4026), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4592), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I78 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4427), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4271), .A(a_man[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I79 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4169), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4014), .A(a_man[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I80 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4366), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4118), .A(a_man[5]), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4169));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I81 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4334), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4180), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4592), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4366), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4608));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I82 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4061), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4026), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4427), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4334));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I83 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4061), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4224));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I84 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I85 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922), .A(a_man[12]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I86 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4623), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4453), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I87 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4041), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4613), .A(a_man[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15725 (.Y(N30312), .A(a_man[4]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15726 (.Y(N30313), .A(N30312));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I88 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4235), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4351), .A(N30313), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4041));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I89 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4204), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4050), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4453), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4235), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4118));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I90 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4247), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4478), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4271), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4204));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I91 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4001), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4247), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4243));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I92 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I93 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I94 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I95 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322), .A(a_man[11]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I96 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4483), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454), .B(a_man[9]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I97 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4103), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4596), .A(a_man[3]), .B(a_man[5]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4613));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I98 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4076), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4103), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4351));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I99 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4120), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3999), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4483), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4144), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4076));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I100 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4180), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4120), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4478));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I102 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015), .A(a_man[10]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I103 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4352), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4193), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I104 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4219), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368), .B(a_man[16]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I105 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3946), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4507), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4193), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4596));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I106 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3985), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4232), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4352), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4014), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I107 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3985), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3999));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I109 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I110 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4006), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4457), .A(a_man[3]), .B(a_man[6]), .CI(a_man[1]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104), .A(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I112 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4249), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4584), .A(a_man[15]), .B(a_man[22]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I113 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4065), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4006), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4249), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4220));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415), .A(a_man[9]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I115 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3970), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415), .B(a_man[7]), .CI(N30313));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I116 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I117 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4532), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4380), .A(a_man[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4183), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4106));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I118 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4574), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4468), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4065), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3970), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4532));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I119 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3919), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4574), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4232));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508), .A(a_man[7]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I122 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4369), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4029), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I124 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4090), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4369), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4029), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4584));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I125 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4624), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4456), .A(a_man[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I126 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4121), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4604), .A(a_man[2]), .B(a_man[5]), .CI(a_man[0]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I127 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4564), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4404), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4624), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4121), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4457));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I128 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4440), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3987), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4090), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4564), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4636));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I129 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4440), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4507), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4468));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I132 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I133 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080), .A(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I134 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4079), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3923), .A(N30313), .B(a_man[13]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I135 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4170), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4016), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I136 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4207), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4053), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4079), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4170), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3995));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I137 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3960), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4524), .A(a_man[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4456), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4604));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I138 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4469), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4207), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3960), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4404));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I139 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4380), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4469), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3987));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I140 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614), .A(a_man[5]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I142 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4355), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4194), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I143 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4549), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4230), .A(a_man[19]), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4355));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I144 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4597), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4476), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4549), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4053));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I145 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3935), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4597), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4338));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I148 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4638), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I149 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4107), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4494), .A(a_man[0]), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4638));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I150 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4392), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4016), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4107), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4230));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I151 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4441), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4289), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I152 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3948), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4510), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4194), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4289), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4494));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I153 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4300), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4115), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3923), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4441), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3948));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I154 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4300), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4476));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428), .A(a_man[3]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15698 (.Y(N30285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15699 (.Y(N30286), .A(N30285));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I157 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3938), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4499), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104), .B(a_man[10]), .CI(N30286));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I158 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4032), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I159 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4472), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4314), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4032), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4158));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287), .A(a_man[4]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15700 (.Y(N30287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15701 (.Y(N30288), .A(N30287));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I161 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4383), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4039), .A(N30288), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I162 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4221), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4069), .A(a_man[17]), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4039));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I163 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4580), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4377), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4383), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4221));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I164 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4238), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4115));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I165 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I166 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I168 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4210), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4056), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958), .B(a_man[9]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I169 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4406), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4393), .A(a_man[16]), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4210));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I170 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4134), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4314), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4406), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4069));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I171 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4134), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4510), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4377));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381), .A(a_man[2]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4488), .A(a_man[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I175 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3963), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4488));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I176 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4251), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4601), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3963), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4393));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I177 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4303), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I178 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4526), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4056), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4149), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3936));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I179 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4162), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4499), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4303), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4526));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I180 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4251), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4162), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3920));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I183 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4267), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I184 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4197), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4047), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I185 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4316), .A(a_man[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I186 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4329), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4174), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4267), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4197), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4316));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I187 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4241), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .A(a_man[1]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I189 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4083), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4198));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I190 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4432), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4533), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4241), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4083));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I191 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4093), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4276));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I193 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4386), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104), .B(a_man[13]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I194 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4139), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I195 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4112), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4139), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4557));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I196 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3992), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4112), .B(a_man[14]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4174));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I197 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3992), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4533));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I198 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I200 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I201 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I202 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949), .A(a_man[0]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I203 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4318), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145), .B(a_man[5]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I204 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3976), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4099), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4227));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I205 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4020), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4047), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3976));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I206 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4020), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4084));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I207 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I208 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4569), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4410), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I209 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4502), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052), .B(N30313), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I210 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4165), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4410), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4336));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I211 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4619), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4569), .B(N30288), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4165));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I212 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4619), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3952), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4437));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I213 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I215 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4035), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4607), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I216 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3967), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I217 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4347), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4189), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4607), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4575));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I218 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4073), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4035), .B(N30286), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4347));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I219 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4539), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4073), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3983));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I221 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4213), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I222 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4155), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4326), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I223 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4529), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4155), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4059), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4092));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I224 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4254), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4455), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4529));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I225 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4010), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4254), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4218));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I226 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I227 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4621));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4087), .A(a_man[9]), .B(N30288));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3931), .A(a_man[9]), .B(N30288));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I231 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4632), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3931));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I232 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4436), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4087), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4632));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I233 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4436), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4189), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4455));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I234 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I235 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4490), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I236 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4024), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4343), .A(N30286), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I237 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3997), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4024), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4326));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I238 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3997), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4376), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3971));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I239 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I240 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3984));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I241 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4202), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4049), .A(a_man[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I242 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4519), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I243 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4591), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4425), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4519), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4343));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I244 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4463), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4556), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4591), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4208));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4463));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4128));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I248 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4481), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I249 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4622), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4481));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I250 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4143), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I251 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4270), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4461), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4049), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4143));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I252 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4622), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4461));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I253 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4270), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4225));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I255 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4512), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I256 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4543), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I257 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4543), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3982), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4587));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I259 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4167), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236), .B(N30313), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I260 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4320), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I261 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4167), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4320), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3978));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I262 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I263 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3945), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I264 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4412), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3998), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I265 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3998));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I266 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4412), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4609));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I269 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4439), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4350), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I270 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4191), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I271 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611), .A(N30288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4439), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4233));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I272 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4191), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4119));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4559), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I275 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4379), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I276 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131), .A(N30286), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4379), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4350));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I277 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I278 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4467), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I279 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4467), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4217));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I280 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I281 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .B(N30288), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4308));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I282 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I283 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949), .B(N30286), .CI(a_man[6]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I285 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I287 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287), .B(N30286));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I289 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I290 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I291 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3961), .A(a_man[1]), .B(a_man[0]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4071), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I296 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4030), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4071), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4226));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I297 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4312), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4184), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3961), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4030));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I298 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4537), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I299 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4137), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I300 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4497), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4537), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4137));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I301 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4578), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3975), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4312), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4497));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I302 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4205), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4617), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4578), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4563), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4196), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4205), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4045));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I305 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4101), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4513), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4563), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I306 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4546), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3951), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4265));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4491), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4110), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4101), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4546));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I310 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4266), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4559), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4491));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I311 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I312 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4173), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4401), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4582), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4173));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I314 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4486), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I315 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4081), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I316 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4306), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4486), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4081));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4583), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4401), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4306));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4330), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4266), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4583));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I319 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I320 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I321 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3944), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4396), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3990));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I322 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4443), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4550), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4330), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3944));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I323 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4301), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I325 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4356), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4301), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4626));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I326 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3918), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4512), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4443), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4356));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I327 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4111), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19007), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3918), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I328 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I329 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4422), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4542), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I330 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4585), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4111), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4422));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4451), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4328), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I335 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4008), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4328));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15727 (.Y(N30315), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4008));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15728 (.Y(N30316), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4161), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405), .B0(N30315));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042), .A(N30316));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I338 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4240), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4240));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I344 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4150), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4637), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4150));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4354), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4637));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4509), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4354));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I349 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I350 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4055), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4055));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I354 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I355 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I357 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3962), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I358 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4534), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3962));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I359 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4324), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4534));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4324));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I361 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I362 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I363 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I364 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4602), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I365 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4602));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4206), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4370));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4363), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4515), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4200), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4363));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I372 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4187), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4025), .A(a_man[19]), .B(a_man[22]), .CI(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I373 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605), .A(a_man[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4528), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4025));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4515), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I378 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I379 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344), .A(a_man[18]), .B(a_man[20]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4187));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I381 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4423), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I384 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I385 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I386 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4102), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4258));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I387 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I388 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I389 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4021), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4423), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4590));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I390 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940), .A(a_man[21]), .B(a_man[19]));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I392 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4021), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I395 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4480), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3916), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4074), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4480), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3916));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I404 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I405 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3981), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I406 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I407 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4040), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4612), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4040));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4140), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4293), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3981), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4140));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4293), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152), .A(a_man[22]), .B(a_man[21]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I417 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253), .A(a_man[22]), .B(a_man[20]));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I419 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4418), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288));
AOI2BB2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I423 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4498), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I424 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4442), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4498));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I425 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4262), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4442));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I426 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4418), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4262));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I427 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253));
OAI2BB2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4482), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4482));
OA22X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921), .B0(a_man[22]), .B1(a_man[21]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I432 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4085), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I436 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4244), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3929), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4085));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I438 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I439 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I442 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I443 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I444 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I445 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I446 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I447 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348), .B(a_exp[4]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I448 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5489));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15730 (.Y(N30323), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5524));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778), .A(N30323));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15702 (.Y(N30289), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15706 (.Y(N30293), .A(N30289));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15705 (.Y(N30292), .A(N30289));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15704 (.Y(N30291), .A(N30289));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15703 (.Y(N30290), .A(N30289));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N750), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17]));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I460 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I464 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I466 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I467 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I471 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I472 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N751), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5389));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I473 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N751), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I474 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18]));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I479 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5500), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I480 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5500));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I481 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N752), .B(N30293));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I483 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I484 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I485 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I486 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I489 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I490 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5400));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I495 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N754), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5513));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N754), .B(N30293));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I498 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I500 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I501 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I502 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I503 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5413));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I504 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N755), .B(N30293));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I505 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I506 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I510 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I511 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I512 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I516 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I521 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I523 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I533 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I540 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I541 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I542 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I543 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I550 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5869), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6057), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6248), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6633), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6171), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5869), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6057));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I576 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I578 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I586 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I594 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I595 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I596 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I599 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I600 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6355), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6521));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I604 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I605 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6483), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6552), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6667));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I619 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6127), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I621 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15732 (.Y(N30329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .A(N30329));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6018), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6197), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6127), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6018), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[28]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6483), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6552), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6197));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255), .A(1'B0), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6074), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6440), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6440));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6538), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I645 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5890), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6156), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6538), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6618), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5890));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[27]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6509), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6156));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I651 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476), .A(1'B1), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[27]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I656 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6033), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6141), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I665 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I666 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6391), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6141), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5959), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6391));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[26]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6033), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5927));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I673 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197), .A(1'B1), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[26]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391), .A(N29673), .B(N29667));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5907), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6174), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5907));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I684 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6635));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I685 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I686 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6458));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I687 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6095), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6557), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6285), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6095));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I701 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6174), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6357), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6525), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5994));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I702 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929), .A(1'B1), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[25]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I704 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4570), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4570), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5548), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5548), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N748), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5477));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N748), .B(N30293));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3942), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3942), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I723 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5501), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I724 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5580), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5580));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N747), .B(N30293));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5378), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5378));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N749), .B(N30292));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8982), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8982));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9472), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I740 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5861), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6237), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6407), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6131), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6237), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6407), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5945));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15744 (.Y(N30373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .A(N30373));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6591), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6591));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[42]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6513));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5980), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I764 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I765 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I766 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6318), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5980), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37720));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I767 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6408), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I768 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6408));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I769 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I770 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6160), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I774 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6347), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I777 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I778 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I779 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5862), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6160), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6347), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5862));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6132), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6318), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6485), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I782 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[24]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[41]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[42]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I786 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I787 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6473), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I788 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I789 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I790 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6301), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I791 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I793 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I794 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6654), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I795 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I796 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6009), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6077), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6473), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6301), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6654), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6009));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I798 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I799 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6189), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I800 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I801 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I802 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[23]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6077), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6189), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6543), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6368));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I805 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I806 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I807 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I808 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5455), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I809 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5454), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5571), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5455), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I810 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5454));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I811 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N746), .B(N30292));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I812 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4037), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I818 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5408), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5407), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5433), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5408), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5407));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I823 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N745), .B(N30292));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I824 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9016), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I825 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9016));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I827 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9506), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I828 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I832 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I833 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6443), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I834 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6078), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I835 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6270), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I836 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6542), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6443), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6078), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6270));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I837 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I838 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9163), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I839 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[41]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[40]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9163));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I840 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[41]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[23]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[41]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I841 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I842 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6334), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6221), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6334));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I844 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5846), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I845 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6395), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5846));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I846 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6499), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I847 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6499));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I848 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5965), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6145), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5965), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6609), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6145));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6221), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6395), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6577), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6036));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I857 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I858 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I860 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I861 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6576), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I862 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6396), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5931), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6576));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I865 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I867 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5505), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I869 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I870 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5575), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5574), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5505), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5575), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5574));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I876 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N744), .B(N30292));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I877 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I878 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I879 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4129), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I880 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4129), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I881 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I882 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I884 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5529), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I885 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5528), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5579), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5529), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5528));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I887 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N743), .B(N30292));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I888 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9052), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I889 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9052));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I890 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I891 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6610), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I893 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I894 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5878), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I895 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5964), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6610), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6066), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5878));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6257), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5964), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6257));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10137), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I900 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9919), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9538), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10137));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I901 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[40]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[39]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9307), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9919));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I902 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[40]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[22]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[40]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I903 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I904 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I905 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I906 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391), .B(N29566));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I907 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6288), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6361), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6099));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I911 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I912 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6677), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I913 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I914 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5912), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I915 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5997), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6677), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6639), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5912));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I916 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[21]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6361), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5997));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9539), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I919 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I920 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I921 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I922 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I923 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I924 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5481), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5480), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5442), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5481), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5480));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N742), .B(N30291));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I931 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I932 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I933 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I934 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4078), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I935 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4237), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15734 (.Y(N30336), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4078), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4237));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394), .A(N30336));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I937 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4005), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I938 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4565), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4005));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I939 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I940 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4214), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4633), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4062));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I941 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I942 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I943 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5437), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I946 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5436), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5437), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I947 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5436));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I948 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N741), .B(N30291));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9083), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9083));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8836), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I954 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9373), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8836));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I955 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9235), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I960 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9056), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8718), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9238), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9235));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6414), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I963 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6322), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6595), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I965 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6678), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6414), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6322), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6595));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I966 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I967 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6135), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I968 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6678), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5951), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6135));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I969 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I970 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9779), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I971 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10126), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9763), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9056), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9779), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8994));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I972 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[39]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[38]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9538), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9373), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10126));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I973 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12222), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12080), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[39]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[21]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[39]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970), .A(N22618), .B(N29506));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5986), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I976 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6051), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5986));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6350), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I978 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6242), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6350));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I979 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6166), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6166));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I981 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6083), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I984 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6277), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I985 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5865), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6083), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6447), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6277));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6051), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6242), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6413), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5865));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9569), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9569), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I990 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I992 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I993 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I994 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5427), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5390), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5427), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I997 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5388), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5390), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5388));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I999 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N740), .B(N30291));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1002 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4000), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4402), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4562));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1004 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1005 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1006 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1007 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5381), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1008 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5556), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5381), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1009 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5555), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5556), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1010 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5555));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N739), .B(N30291));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1012 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9121), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1013 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9121));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1016 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1017 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8769), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8867));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1018 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6117), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5898), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6117));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6305), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1025 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1026 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1027 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6659), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1028 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6305), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6477), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6659));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1029 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5898), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6448), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6012), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6084));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1032 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1033 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9392), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1034 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8844), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8769), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9392), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8718));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1035 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1036 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6339), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1038 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5970), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6149), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6339));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1039 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1040 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1041 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6502), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5851), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6502), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1043 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6227), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5851));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1044 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1046 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1047 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1048 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1049 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9271), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9299), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1053 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8694), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10206), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9271), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9299));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1054 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9509), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9010), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9814), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8694));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1055 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1056 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6492), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1057 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6387), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6492));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1058 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6387), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5838), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5838));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1061 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5918), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1062 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1063 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1064 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1065 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6028), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6212), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142));
NOR3X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1066 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6102), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6000));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1067 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1068 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1069 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1070 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9600), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1073 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1074 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1075 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9702), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1076 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1077 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1078 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1079 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5547), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5509), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5547), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5508), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5509), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5508));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1083 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N738), .B(N30291));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15736 (.Y(N30343), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934), .A(N30343));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1085 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4492), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1086 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4492), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5499), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1090 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5463), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5499), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1091 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5462), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5463), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5462));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1093 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N737), .B(N30290));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1094 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9157), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1095 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9157));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1097 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8904), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1099 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10280), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9926), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9702), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8904));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1100 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10159), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9796), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8679), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9429), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10280));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1101 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10249), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9890), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10159), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10103), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9116));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1102 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9601), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10185), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9509), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10249));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1103 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[38]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[37]), .A(N23335), .B(N23333), .CI(N29612));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1104 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446), .A(N23142), .B(N23140), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[38]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1105 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323), .A(N29502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1109 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6340), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1113 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6306), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6340));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6584), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1115 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6478), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6584));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1116 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6228), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1117 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6306), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6478), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6228));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6400), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5936), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6116), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6658));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1119 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9044), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9853), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6016), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1124 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6247), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6016));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1125 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1126 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1127 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6373));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1128 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6169), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1129 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5901), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6548), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6418), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5901), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6548), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1132 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6247), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5990), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6353), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6418));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1133 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1134 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1135 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9318), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9853), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9991));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1136 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9181), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8821), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9318), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9796));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1137 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1138 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8708), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1139 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1140 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9463), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6153), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1142 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6505), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6342), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6153), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6505), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6342));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5853), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6043), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5853), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6232), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1148 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6587), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6043), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6232));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1149 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1150 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1151 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10194), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9835), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8708), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9463), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9618));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1152 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1157 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8726), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9313), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9365));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1158 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10073), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9709), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10194), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8726), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9926));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1159 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9885), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1161 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1165 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9582), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9885), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8936), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9075));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1166 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1168 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1169 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1171 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5373), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5453), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5373), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5418), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5453), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5417), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5418), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N736), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5417));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N736), .B(N30290));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1180 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4594), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4594), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1183 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5541), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1184 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5406), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5541), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1185 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5584), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5406), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1186 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5583), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5584), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N735), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5583));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N735), .B(N30290));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9196), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9196));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5922), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6107), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6468), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5922), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6107), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6468));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1196 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6293), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1197 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6647), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1198 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6003), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1200 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5887), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6293), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6647), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6184), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6003));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1201 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5887));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1202 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1203 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1204 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8828), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10165), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9740), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9230));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1205 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9221), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8852), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9582), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8828), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10045));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1206 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9089), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9221), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8940), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9709));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1207 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9954), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9574), .A(N23945), .B(N23943), .CI(N29496));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1208 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9279), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8909), .A(N29498), .B(N23579), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9954));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1210 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1211 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1212 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1213 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1215 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1217 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7522), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7554), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7670));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1218 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1219 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7595), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1224 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1225 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7986), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1226 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7754), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7595), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7986));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1227 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7568), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7754));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7685), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8043), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1232 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7861), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1233 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7821), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7685), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8043), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7861));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1234 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7888), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1235 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7821), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7888), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7626));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1236 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1237 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1238 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1239 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1240 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1241 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7648), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7957), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7744));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1242 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1243 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7794), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7546), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1247 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8039), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7915), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7527), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7546), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7667));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1248 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7894), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7910), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7794), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8039));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1249 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7703), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7648), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7894));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1251 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1252 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8077), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1255 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7615), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7867), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8077), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8060));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1256 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1257 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8035), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7847), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1260 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7981), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1261 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7864), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8035), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7847), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7981));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1262 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7723), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7594), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7613), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7864));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1263 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7723), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7521), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7771));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1264 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1265 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1266 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7599), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1269 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7765), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7732), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7599), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7741));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1270 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7541), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7987), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8062), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7765), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7747));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1271 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7915), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7594));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8049), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1276 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1277 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7905), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7782), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7745), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8049), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7539));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1278 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7801), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1279 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7677), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1280 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1281 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1282 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7556), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8001), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7801), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7677), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8073));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1283 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8057), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1287 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1288 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7803), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7684), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8061), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7859), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7693));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1289 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7586), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8030), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7556), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8057), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7803));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1290 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7695), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7905), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7586));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1291 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7788), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7938), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7811), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1296 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7662), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7533), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7938), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7811));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1297 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8009), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7887), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7788), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7662));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1298 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7695), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8009), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7987));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1299 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1300 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1301 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1302 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7822), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7551), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1305 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8019), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7896), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7822), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7551), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7588));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1306 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7560), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1310 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7772), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7650), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7994), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7560), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7565));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1311 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8052), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7926), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8019), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7772), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8001));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1312 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7832), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7715), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7782), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7533), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8052));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1313 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7832), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7887), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7567));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1314 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1315 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7813), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1316 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7873), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1319 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1320 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7989), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7865), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7577), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7873), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7992));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1321 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7705), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7813), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7611), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7989));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1322 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1323 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7932), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1325 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7674), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7544), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7932), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7906));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1326 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7947), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7824), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7674), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7896));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1327 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7736), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7605), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7684), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7947));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1328 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8030), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7715));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1329 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1330 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7624), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8068), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5456), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1335 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5494), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5456), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1336 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5573), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5494), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5537), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5573), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1338 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5536), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5537), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5536));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N734), .B(N30290));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[1]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15707 (.Y(N30294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15715 (.Y(N30302), .A(N30294));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15714 (.Y(N30301), .A(N30294));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15713 (.Y(N30300), .A(N30294));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15712 (.Y(N30299), .A(N30294));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15711 (.Y(N30298), .A(N30294));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15710 (.Y(N30297), .A(N30294));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15709 (.Y(N30296), .A(N30294));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15708 (.Y(N30295), .A(N30294));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7885), .A(N30302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1343 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7959), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7834), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7624), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8068), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7885));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1344 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15716 (.Y(N30303), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15724 (.Y(N30311), .A(N30303));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15723 (.Y(N30310), .A(N30303));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I15722 (.Y(N30309), .A(N30303));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15721 (.Y(N30308), .A(N30303));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15720 (.Y(N30307), .A(N30303));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15719 (.Y(N30306), .A(N30303));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15718 (.Y(N30305), .A(N30303));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15717 (.Y(N30304), .A(N30303));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8007), .A(N30311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7886), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7664), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1349 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7889), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7767), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7886), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7690), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7664));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1350 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7916), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7793), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7959), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8007), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7889));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7895), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7582), .A(N30311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1354 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7642), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8088), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7895), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7582));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1355 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7596), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8041), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7865), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7642), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7544));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1356 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7628), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7916), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7596));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1357 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7628), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7605));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1358 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1359 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7815), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8088), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7834), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7767));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1361 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1362 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1363 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7606), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7649), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7943), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7639));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1364 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059), .A(N30302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1365 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4028), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4429), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4598));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1372 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3956), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4367), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4028), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4520));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3956), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5410), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N608), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5447), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5410), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5527), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5447), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5490), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5527), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1378 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5488), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5490), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1379 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5488));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N733), .B(N30290));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1381 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7764), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7900), .A(N30311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1384 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7855), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7764), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7977), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7900));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1385 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7569), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7687), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7855));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1386 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7843), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7727), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7815), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7569), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7793));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1387 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7843), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7824), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8075));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1388 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1389 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1390 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7797), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1392 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7558), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7724), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7702), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1395 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7652), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7724), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7702));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7816), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7967), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1399 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7580), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8021), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7816), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7967), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7737));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1400 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7534), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7558), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7652), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7580));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7809), .A(N30302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7762), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7655), .A(N30311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1404 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7898), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7762), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7655));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1405 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7783), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8054), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7898), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7738));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1406 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8064), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7534), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7783));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1407 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8064), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8041), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7727));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7564), .A(N30301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7570), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1411 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7868), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7564), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7570));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1413 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7826), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7706), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7868), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7955), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7524));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8053), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7714), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7770), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1417 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7791), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1418 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7515), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7962), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7770), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7791));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1419 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7796), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8053), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7714), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8038), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7725), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7971), .A(N30311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1423 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7548), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7993), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7725), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7971));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1424 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8078), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7949), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7796), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7548), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8021));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1425 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8031), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7907), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7826), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8078));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1426 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8031), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7697), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7936));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1427 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7890), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8040), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7730), .A(N30310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1432 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7768), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7644), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7890), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8040), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7730));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8029), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7884), .A(N30301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7804), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1436 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8013), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7891), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7884), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7804));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1437 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8044), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7768), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7750), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8013));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1438 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7757), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7774), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7706));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1439 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7757), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7665), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7907));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7637), .A(N30301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1442 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1443 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7983), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7858), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7637), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7643));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1444 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1445 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7792), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1446 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1447 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7668), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7537), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7542), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7792), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7557));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1448 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7698), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7962), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7983), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7668));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1449 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7729), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7993), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7698));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1450 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7729), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7631));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7862), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1456 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7881), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7862), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7543));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8046), .A(N30310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1458 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7912), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7786), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7881), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8046), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7858));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1459 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7939), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7817), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7912), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7644), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7891));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1460 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7939), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7918), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7598));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7877), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1464 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7713), .A(N30301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7718), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1466 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8024), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7901), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7713), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7718));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1467 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7806), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7689), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7877), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7532), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8024));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7954), .A(N30301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7961), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7798), .A(N30310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1471 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7561), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8005), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7961), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7798));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1472 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7591), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8034), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7806), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7561), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7537));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1473 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7591), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7571), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7817));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1474 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7575));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7549), .A(N30310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1479 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7710), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7630), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7616), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7549));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1480 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8058), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7930), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7710), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7760), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8005));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1481 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8058), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7786), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8034));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19018), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1483 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1484 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1485 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7601), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8047), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7935), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7617));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1486 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8027), .A(N30300), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8033), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1489 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7848), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7731), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8027), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8033), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7948));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1490 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7951), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7828), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7901), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7601), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7848));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1491 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7951), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7689), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7930));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7785), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1495 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7996), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7871), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7780), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7785));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7870), .A(N30310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1497 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7528), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7972), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7996), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7870), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8047));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1498 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7528), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7828));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1500 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7621), .A(N30309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1501 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1502 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1503 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1504 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7819), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8010), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7536));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1505 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7678), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7621), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7694), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7819));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1506 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7731), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7678), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7972));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7883), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8020), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7531), .A(N30300), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1510 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7941), .A(N30309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1511 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8069), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7942), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8020), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7531), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7941));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1512 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8069), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7871), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7550));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7851), .A(N30300), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7766), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1516 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7892), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7851), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7766));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1517 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7892), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7942));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1521 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7965), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7840), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8084), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7608));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7699), .A(N30309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1523 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7965), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7699), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7769));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8014), .A(N30309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7604), .A(N30300), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1527 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7604), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7840));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7925), .A(N30300), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7833), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1531 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7833));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7779), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1533 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7681), .A(N30299), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1535 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7587), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7681));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517), .A(N30309));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7850), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(N30299), .C(N30308));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1540 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7721), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7850), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7612), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1541 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7974), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1542 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7573), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7530), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7721), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7974));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1543 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7921), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7779), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7573), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7903), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7709), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8026), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7921), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7903));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7982), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7712), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7709), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7830), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8083), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7911), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7830), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8083));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1550 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7911));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7795), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7953), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7982), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7520));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7686), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7883), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7795), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7660), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8006), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7692));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7673), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7563), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7686), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7660));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7931), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19018), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7673), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8016), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7610), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8016), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7701));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7743), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7931), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7610));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7623));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7552), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7538), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7552));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7818), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7538));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7940), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7818));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8048), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8048));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8036), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7973));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1576 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8036));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1578 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7902), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7902));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7829), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7963), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7829));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7751), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7963));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7676), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7751));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7797), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7676));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1586 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7761), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7645), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7761));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7645));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7929));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8076), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7807), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[32]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7807));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1594 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1595 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10214), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9468), .A(N29614), .B(N29598));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1596 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10214));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9468));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1599 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[37]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[36]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9279), .B(N29610), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10192));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1600 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[37]), .B(N23130), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[37]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1604 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37712));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1605 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6133), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6133));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6182), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6182));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5917), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5917), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6292), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6103));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5882), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6261), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6534));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5942), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6125), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6664), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6017), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5942), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6125), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6313), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6664));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1619 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6482), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8851), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6017), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6482));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1621 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9692), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .A1(N30268), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1622 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9347), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1627 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9162), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8801), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10276), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9347), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9433));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10027), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5870), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6140), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6522), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5870), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6058));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6250), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6603), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6420), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6140), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6250), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6603), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6420));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1645 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8945), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10286), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8859), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9503), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8738));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1646 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8648), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10027), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8945));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9668), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9266), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1654 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9526), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9134), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9774), .B(N30308), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9266));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1656 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9923), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1663 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10263), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9904), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9923), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8971), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9111));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1664 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9716), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9326), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9526), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9660), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10263));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1665 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9354), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9191), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10165), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9716));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1666 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9983), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8648), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9835), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9354));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6315), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6484), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6668), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1673 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6315), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6484), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6668));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6020), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6378), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6199), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6554), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6020), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6378), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6199));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10199), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9386), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1684 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10089), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9726), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9386), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1685 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9294), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10199), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10089));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1686 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8748), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10286), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8801), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9294));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1687 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10109), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8748), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9960), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8977));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1688 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9004), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8671), .A(N29490), .B(N24432), .CI(N29655));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1689 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9862), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9478), .A(N29494), .B(N29492), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9004));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6438), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6537), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6155), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6073), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6267), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6438), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6537));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10191), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6155), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6617), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5975));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8925), .A0(N30266), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30268));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1699 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8967), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10303), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9862), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9574), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8925));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1700 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[36]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[35]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8909), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8967));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1701 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[36]), .B(N23120), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[36]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1702 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1704 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7897), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7651), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7773));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[30]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9596), .A(N29592), .B(N29580));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9596), .B(N29598));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6570), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6109), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6032), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6570), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6497));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5924), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9832), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6109), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5924), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6390));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9909), .A0(N30264), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30266));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1723 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1724 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5858), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6075), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6269), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6619));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6441), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6157), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5978), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5858), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6441), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6345), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6157));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9844), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390));
NAND2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[1]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962), .AN(N30299), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808), .A(N30308), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1740 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9913), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1741 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8895), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9844), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9693), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9913));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8896), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9541), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8762), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1748 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9877), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9496), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8896), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9541), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8762));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1749 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10050), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8895), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9877), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9134));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1750 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9486), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10050), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10079));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10235), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9766), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .S0(N30299));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9421), .A(N30308), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1758 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9732), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9340), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9421));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1761 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8737), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10235), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9732), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10098));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1764 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1765 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1766 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1767 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1768 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9695), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9301), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9955), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9007), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9148));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1769 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9659), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9695), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9726));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1770 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9072), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8731), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9904), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8919));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6034), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5843), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1774 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5928), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6034), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5843), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5928));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1777 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6392), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6219), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1778 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6573), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1779 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6392), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6573));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9457), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1782 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9576), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8673), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1786 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8764), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10097), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8673), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9340));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1787 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9462), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9078), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9530), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9457), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8764));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1788 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8710), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9496), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9462));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1789 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9843), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9456), .A(N25768), .B(N25766), .CI(N29486));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1790 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10229), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9869), .A(N29624), .B(N29488), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9843));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1791 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9127), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8776), .A(N29653), .B(N29626), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10229));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1793 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6423), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1794 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1795 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6251), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1796 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5872), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6423), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6251));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9137), .A0(N30262), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30264));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1798 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9771), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9382), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9127), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8671), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9137));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1799 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8880), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10221), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9478), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9771));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1800 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[35]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[34]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10303), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8880));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1801 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6137), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1802 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6417), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6599), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1805 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1806 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6493), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6417), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6599), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6325), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5953));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1807 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[17]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6137), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6493));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1808 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[35]), .B(N23110), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[35]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1809 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1810 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6374), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1811 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6549), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1812 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5900), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6088), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6374), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6549), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5900), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6088));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6452), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5991), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6452), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10251), .A0N(N29592), .A1N(N29580), .B0(N29598));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1818 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10251));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908), .A(N29592), .B(N29580));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1823 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8042), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1824 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1825 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1827 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7919), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8045));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1828 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7633), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7759));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7597), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7728), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8042), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7597));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1832 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7728), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1833 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[27]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1834 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9495), .A(N29426), .B(N29570));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1835 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9495), .B(N29580));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1836 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1837 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1838 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6671), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1839 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6094), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1840 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1841 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6457), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6671), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6094), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5906));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1842 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9064), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6556), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6457));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10118), .A0(N30260), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30262));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1844 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1845 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1846 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1847 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6359), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1848 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5908), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5908));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5995));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6254), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5874), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6062), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6636));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6175), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6359), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6527), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6254));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1857 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1858 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8793), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1860 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9502), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9070), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8793));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1861 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10208), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9852), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9502), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10058));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1862 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9428), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9043), .A(N26246), .B(N26244), .CI(N26248));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1865 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1867 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9493), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1869 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9312), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10129), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10267), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9493));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1870 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9986), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .S0(N30299));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9040), .A(N30308), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9186), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1876 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10278), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9922), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9986), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9040), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9186));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1877 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9274), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8903), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10278), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10097));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1878 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1879 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9878), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1880 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1881 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1882 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1884 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1885 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5947), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1887 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6409), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1888 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6592), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6409), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1889 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6486), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6239), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5947), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6592));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1890 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6486));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1891 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1893 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9540), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9338), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9376), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8732));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1894 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10243), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9886), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9878), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9733), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9540));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1895 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9237), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8866), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9274), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10243), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9078));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1900 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6544), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1901 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5893), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1902 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1903 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6272), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6079), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1904 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6544), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5893), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6272));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1905 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1906 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10051), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1907 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9575), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9102), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9613), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10051));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .S0(N30298));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8702), .A(N30307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1911 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1912 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9799), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9414), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8702), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10216));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1913 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1914 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8823), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1915 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1916 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8961), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9914), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1919 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10306), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8961), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9914));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1920 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10068), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9575), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9799), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10306));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1921 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10035), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10068), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9110), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9886));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1922 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9999), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9629), .A(N26208), .B(N26206), .CI(N29478));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1923 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10170), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9816), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9043), .B(N29480), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9999));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1924 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8858), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9456), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9428), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10170));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7866), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7545), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7866), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7991));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1931 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9396), .A(N29560), .B(N29430));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1932 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9396), .B(N29570));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1933 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9257), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8887), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8858), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9869), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1934 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9896), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10118), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8776), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9257));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1935 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8796), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9382), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9896));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1936 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[34]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[33]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10221), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10067), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8796));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1937 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[34]), .B(N23100), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[34]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1938 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1939 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1940 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1941 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1942 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6615));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1943 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6044), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6044));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1946 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6436), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1947 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1948 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6265), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6436), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5973));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5886), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5854), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5886));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6311), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5941), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6123), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6588), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5854));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1954 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6231), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6311));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1955 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9309), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9319), .A0N(N29426), .A1N(N29570), .B0(N29580));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1960 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9319));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707), .A(N29426), .B(N29570));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1963 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9118), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1965 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8915), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9118), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9518));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1966 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[33]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[32]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10132), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9699), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8915));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1967 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[33]), .B(N23090), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[33]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1968 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1969 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1970 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1971 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1972 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6569), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1973 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6216), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6108), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6569), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6294));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15738 (.Y(N30352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6648), .A(N30352));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5921), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6183), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6467), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6648));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1978 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1979 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6541), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1981 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6512), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6188), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6541));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5892), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5979), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1984 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1985 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5860), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6007));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6236), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6512), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5892), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5979), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5860));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9363), .A0(N30258), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30260));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8768), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1990 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10017), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9650), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8887), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9363), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8768));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1992 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1993 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6428), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1994 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I1996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6428), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6608), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6144));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1997 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I1998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6498), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15740 (.Y(N30360), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5845), .A(N30360));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10044), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6220), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5963), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6498), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5845));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8659), .A0(N30256), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30258));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2002 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9085), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9922), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9149), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8935));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2004 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2005 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2006 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10300), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2007 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2008 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2009 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8672), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10161), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10300), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9531));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2010 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10105), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9414), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8672), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9185));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .S0(N30298));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2012 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10018), .A(N30307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2013 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9377), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2016 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9838), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9450), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10018), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9377), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10275));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2017 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2018 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9765), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9223), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6335), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2025 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5847), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2026 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6500), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2027 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6222), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6611), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6335), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5847), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6500));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2028 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6146), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2029 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6038), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6222), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6146), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6038));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2032 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9685), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2033 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9612), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8756), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9685));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2034 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9348), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9838), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9765), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9612));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2035 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9860), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9469), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10105), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9348), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9703));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2036 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9051), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8714), .A(N26238), .B(N26236), .CI(N29484));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2038 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8998), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2039 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2040 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2041 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2043 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8890), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8998), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9138), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2044 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9297), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2046 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .S0(N30298));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2047 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9654), .A(N30307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2048 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9872), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9297), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9654));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2049 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8855), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5913), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2053 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6460), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2054 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6562), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5913), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6460));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2055 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6289), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2056 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6178), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6289), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2057 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2058 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2061 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9653), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9260), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8855), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9295), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9948));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2062 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9385), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8890), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9872), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9653));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2063 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9120), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9385), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9956), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8970));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2064 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8873), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10218), .A(N29476), .B(N26198), .CI(N29482));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2065 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9823), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9434), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8873), .B(N25627), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8714));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2066 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9019), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9629), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9051), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9823));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2067 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2068 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7937), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2069 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2070 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[23]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9291), .A(N29442), .B(N27939));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9291), .B(N29430));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2073 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9201), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8835), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9019), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9816), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2074 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9620), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8659), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9201));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2075 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9037), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9620), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9650));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2076 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[32]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10256), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10017), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9037));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2077 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[32]), .B(N23080), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[32]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2078 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2079 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6356), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2083 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5871), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2084 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2085 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6356), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5871), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6059), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2086 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6249), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6421), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6604), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6331), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6249), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6421), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6604));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2090 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2091 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6382), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6560), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2093 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6638), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6206), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6382), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6560));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2094 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5911), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2095 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5911), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2097 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9677), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6098), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6287));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9595), .A0(N30254), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30256));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2099 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10110), .A0N(N29560), .A1N(N29430), .B0(N29570));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2100 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10110));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2102 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775), .A(N29560), .B(N29430));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9547), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2105 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9967), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9591), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8835), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9595), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9547));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6082), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6165), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37704), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6165), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2109 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5950), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6082), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37704));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6274), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6446), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6241), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6274), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6446));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2113 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2115 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9284), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5950), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6241), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6625), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5984));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2116 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8839), .A0(N30244), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30254));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2117 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10134), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9224), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9450), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9985));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5987), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2119 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6167), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6053), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6449), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2124 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6628), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6243));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2125 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6053), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5952));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2126 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6167), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19032));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2127 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2128 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2129 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2132 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2133 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9689), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9296), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8667), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9568));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2134 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9423), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9039), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9689), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10231));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2136 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2137 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2138 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2139 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9135), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8783), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8666));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2140 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9800), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2142 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .S0(N30298));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9261), .A(N30307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8787), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9727), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2148 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8922), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10264), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9261), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8787), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9727));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2149 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8701), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10021), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9135), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9800), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8922));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2150 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9156), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8798), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8701), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9006));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2151 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9891), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9511), .A(N26760), .B(N26758), .CI(N29456));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2152 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8719), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2157 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10146), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9789), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9032), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9176), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8719));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2158 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2159 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2161 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9333), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2165 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9981), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2166 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9944), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10121), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9333), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9981));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2167 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8733), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10195), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9944));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2168 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6041), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2169 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2171 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6041), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6229), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5937));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6401), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6401), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6479), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6585), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6119));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .S0(N30298));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8888), .A(N30307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2180 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9836), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2182 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8955), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10261), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8888), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9836));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2183 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9460), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8783), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8955), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10264));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2184 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10167), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9807), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8733), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9260), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9460));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2185 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9928), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9551), .A(N29468), .B(N26654), .CI(N29454));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2186 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8911), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9511), .B(N29474), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9928));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2187 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9636), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10218), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9891), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8911));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6040), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6399), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6226), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6399), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6582));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6114), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8914), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6114), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5935));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2196 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9821), .A0(N30252), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30244));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2197 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8840), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10179), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9636), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9434), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9821));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2198 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9787), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8839), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8840));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2200 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2201 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2202 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2203 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8981), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8656), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9787), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9738), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9921));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2204 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9391), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9229), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8981));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2205 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2206 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2207 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2208 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2210 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10273), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2211 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8678), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10102), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9927), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10273));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2212 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[31]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[30]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9391), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8678), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8699));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2213 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[31]), .B(N23070), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[31]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2215 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9161), .A0N(N29442), .A1N(N27939), .B0(N29430));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9161));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2217 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2218 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555), .A(N29442), .B(N27939));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2219 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2224 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2225 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8810), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8976), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9154), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9345));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2226 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9753), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9360), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9591), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8810), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8656));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2227 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[30]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9990), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9012));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6021), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6669), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6316), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2232 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6129), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6669), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6316), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2233 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6379), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2234 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2235 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6021), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6092), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6379), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6198));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2236 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[30]), .B(N23060), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[30]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2237 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2238 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2239 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2240 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2241 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2242 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6364), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2243 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6069), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5881), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6181), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6364), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6069), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5881));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6260), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2248 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10255), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6532), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6260));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2249 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9049), .A0(N30250), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30252));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2251 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2252 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2255 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9758), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2256 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9207), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8841), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8696), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8814), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9758));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2257 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8784), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2260 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10182), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9824), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8784), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9451));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2261 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .S0(N30297));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2262 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10232), .A(N30306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2263 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2264 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2265 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2266 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9605), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2267 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9977), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10232), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8951), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9605));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2268 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9729), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9335), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9207), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10182), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9977));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2269 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10202), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9846), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9729), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9296), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10054));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2270 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9195), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8830), .A(N26768), .B(N26766), .CI(N29464));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2271 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8758), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9565), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9789), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10295));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .S0(N30297));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9873), .A(N30306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2276 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2277 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .S0(N30297));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2278 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9488), .A(N30306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2279 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10042), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9674), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9488));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2280 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9027), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10012), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9873), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10042));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2281 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9761), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8841), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9824), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9027));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2282 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2283 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2287 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9247), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8876), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9755), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10154));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2289 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9905), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2290 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2291 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9068), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2296 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10008), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9638), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9368), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9068), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10294));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2297 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8991), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9247), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9905), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10008));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2298 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9497), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9105), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8991), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9335));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2299 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9231), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8861), .A(N26752), .B(N26750), .CI(N29460));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2300 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9962), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9231), .B(N29466), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8830));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2301 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8942), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10282), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9195), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9962));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2302 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7836), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7526), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7654), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2305 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7526), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7654));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2306 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8089), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7836), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7960));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8089), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2310 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[19]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2311 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2312 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9153), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9092), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[21]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2314 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9672), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8942), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10252), .CI(N30224));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2315 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8689), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9049), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9672));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2316 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8661), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9974), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10179), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8649), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8689));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9537), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2319 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2320 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8797), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2321 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8012), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2322 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8012), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2323 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9193), .A(N29392), .B(N28088));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9193), .B(N27939));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2325 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2326 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2327 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9597), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9205), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8797), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8966));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2328 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9563), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9400), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9537), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9597));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2329 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10293), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10144), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8661), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9169));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2330 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[29]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10293), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9563), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9360));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6510), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2335 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6346), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2336 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6620), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5977), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6158), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6346));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[11]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6510), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5859));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2338 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[29]), .B(N23050), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[29]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8792), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10305), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2344 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10153), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9792), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8792), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10305), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10006));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9581), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2349 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9966), .A0N(N29392), .A1N(N28088), .B0(N27939));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2350 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9966));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655), .A(N29392), .B(N28088));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2354 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9393), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2355 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9441), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9581), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9769), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9393));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6279), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2357 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2358 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2359 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6168), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6279), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6629), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5989), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6168));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2361 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6519), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2362 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6351), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2363 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9517), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5867), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6519), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6351));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2364 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6324), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2365 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6491), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5837), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6211), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6324), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6491), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5837), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6211));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6385), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9894), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6565), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6026), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6385));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2372 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9270), .A0(N30248), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30242));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2378 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9644), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2379 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9831), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9444), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9941), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8989), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9644));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2381 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8727), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8848), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2384 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2385 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9793), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2386 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9062), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8723), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8848), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9793));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2387 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9794), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9408), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9831), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9062), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8876));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2388 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8789), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9794), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9598), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8663));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2389 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10237), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9881), .A(N29452), .B(N26704), .CI(N29458));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2390 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9994), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8861), .B(N29462), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10237));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7909), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2392 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753));
NAND2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .AN(N28113), .B(N28313));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2394 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8978), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8650), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9585), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9994), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2395 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9711), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10282), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9270), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8978));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10031), .A0(N30242), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30250));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2397 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8721), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10040), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9711), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10031), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9280));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10131), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9778), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2404 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9407), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9024), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9959), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10131), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9778));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2405 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9175), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8815), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9441), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8721), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9024));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2406 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10120), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10153), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9974), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9175));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2407 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9145), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2409 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9367), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8988), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9407), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9145), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9205));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2410 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[28]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[27]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9367), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9940));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6472), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6472));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6393), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6297), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2417 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6005), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6111), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6393), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6297));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[10]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6367), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6005));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2419 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[28]), .B(N23008), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[28]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2423 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2424 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2425 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2426 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2427 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10188), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9829), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9953), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10040));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2432 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9480), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9192), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9321));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9383), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9017), .A0N(N28287), .A1N(N30226), .B0(N28088));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2436 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9017));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2438 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402), .A(N28287), .B(N30226));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2439 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8833), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2442 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9572), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2443 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8745), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8833), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9572));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2444 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9215), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8847), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9480), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8745), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9059));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2445 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9950), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9792), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10188), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9215));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2446 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[27]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9950), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8988), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9760));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2447 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2448 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6526), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5876), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6063), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6253), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6063), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6526), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5876), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6253));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[9]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5960));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2454 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[27]), .B(N22949), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[27]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2456 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6586), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6661), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6230), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6586), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5940));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2460 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6309), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9125), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6121), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6309));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10241), .A0(N30246), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30248));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2464 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2466 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9748), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9356), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10241), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10172));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2467 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9762), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9003), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2471 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2472 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9404), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2473 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .S0(N30297));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2474 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9099), .A(N30306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10048), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2477 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8884), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9404), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9099), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10048));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2479 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9683), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9203));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2480 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9969), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2481 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2483 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9866), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9482), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9969), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9252));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2484 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8850), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10190), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8884), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9866), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9674));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2485 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8816), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10156), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9638), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8850));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2486 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9533), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9143), .A(N26230), .B(N26228), .CI(N29450));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2488 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9268), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9533), .B(N30232), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9881));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2489 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5884), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2490 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6465), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6071), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6646), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6465), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6071));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2495 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6435));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5884), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19025));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9498), .A0(N30240), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30246));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2498 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9013), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9623), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9498));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2500 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2501 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8778), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9013), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9183));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2502 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10223), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9864), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9748), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9762), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8778));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2503 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2504 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8676), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2505 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2506 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8827), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715), .A(N30250), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2509 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9520), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8827), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9375));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2510 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9251), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8883), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10075), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9520), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9093));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2511 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9980), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9604), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9829), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10223), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9251));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2512 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[26]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9980), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8815), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9567));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6319), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6673), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2516 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6488), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6558), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5948), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6319), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6673), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6488));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6023), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6558), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6023), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6203));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2521 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[26]), .B(N23035), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[26]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2523 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9815), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .A(N30226));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669), .A(N28313));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133), .A(N30268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2533 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10189), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .S0(N30297));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8750), .A(N30306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2538 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8728), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10049), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8882), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9292), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8750));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2539 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9647), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9254), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10189), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8728));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2540 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9607), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9444), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8723), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9647));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2541 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9571), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9179), .A(N26254), .B(N26252), .CI(N26256));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2542 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10034), .A(N30232), .B(N23556));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2543 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10271), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9917), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9571), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10034), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9143));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6419), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6056), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6030), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6419), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6056), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6601), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2550 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5955), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6030), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6139), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8761), .A0(N30234), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30240));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2552 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10029), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8899), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10271), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8761));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2553 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9781), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9395), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9815), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9628), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10029));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2560 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8803), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8670), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9992));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2561 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10257), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9356), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9781), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8803));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8820), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8996), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2566 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9558), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8680), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8820), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8996));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2567 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9288), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8916), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10111), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9558), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9129));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2568 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10013), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9864), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10257), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9288));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2569 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[25]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10013), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8847), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9604));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5895), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6271), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6444), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6514), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5895), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6271), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6622), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6444));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2576 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6514), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5982), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6161));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2578 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[25]), .B(N22939), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[25]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9805), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2586 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9818), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9431), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9805), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9984), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9619));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9427), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196), .A(N30268), .B(N30266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9272), .A(N30232), .B(N23859));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2594 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2595 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9828), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2596 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9681), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2598 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9454), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9069), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9025), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9828), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9681));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2599 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8697), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9482), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9454), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10226));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2600 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8668), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8697), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9217));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2601 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10301), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9272), .B(N29622), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9179));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6019), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2604 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6377), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2605 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6282), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6019), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6666), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6377));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6553), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5903), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6553), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9745), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6282), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6196), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5903));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9731), .A0(N30238), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30234));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2611 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9305), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8930), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9917), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10301), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9731));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2612 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9047), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9427), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9236), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9305));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2613 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10287), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9818), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9047), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9395));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610), .A(N30250), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841), .A(N30248), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2618 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8838), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10174), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9663), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10158), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8665));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2619 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9328), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8947), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10139), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8838), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9164));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2620 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10047), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9899), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10287), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9328));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2621 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[24]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[23]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10047), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8883), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9643));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2622 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6474), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6578));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6655), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5933));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15742 (.Y(N30368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I15743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6112), .A(N30368));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6112));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5848), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6223), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6302), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5848), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6223), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6037), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6397));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6474), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6655), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6010), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6302));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2634 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[24]), .B(N22929), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[24]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9419), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9228), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2645 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9081), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9419), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9609), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9228));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259), .A(N30266), .B(N30264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8868), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10245), .A(N30232), .B(N23861));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2656 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9263), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8892), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10175), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9442));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .S0(N30296));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10080), .A(N30305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2665 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10023), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9657), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8690), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10224), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10080));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2666 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10197), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9840), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9263), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9975), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10023));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2667 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9417), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9035), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9254), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10197), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10015));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2668 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9379), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10245), .B(N29472), .CI(N29620));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6344), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6508), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5857), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2673 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5976), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6344), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6508), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5857));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9352), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6045));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8957), .A0(N30236), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30238));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2677 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9341), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9951), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9379), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8957));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2678 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10062), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9045), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8868), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9341));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2679 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9593), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9081), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10062), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8711));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9798), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902), .A(N30246), .B(N30240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9979), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2684 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9856), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9465), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9798), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9979));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2685 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8657), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9431), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9856), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10174));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2686 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10082), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9718), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9593), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8657));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2687 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[23]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10082), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8916), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9680));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5879), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5879));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5998), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6362), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5998), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6530), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6362));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[5]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5966), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6429));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2696 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[23]), .B(N23018), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[23]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513), .A(N30250), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2701 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2702 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8860), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2704 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9113), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8765), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9036), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9220), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8860));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8709), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651), .A(N30264), .B(N30262), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9501), .A(N30232), .B(N24239));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9865), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .S0(N30296));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9719), .A(N30305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2716 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9625), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9060), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9865), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9719));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9430), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8917), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2720 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8863), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8917));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2721 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9042), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8705), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9625), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8863), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8892));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2722 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9227), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8857), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9069), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10049), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9042));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2723 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10163), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9501), .B(N26646), .CI(N29470));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2724 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6572), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5926), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5926), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6471), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6186), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6572), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6110), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6471));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6296), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8975), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6186), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6296), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6651));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9947), .A0(N30230), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30236));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2733 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10130), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9767), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10163), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9947));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2734 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10100), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9735), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8709), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10207), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10130));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2735 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8870), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10211), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9113), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10100), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9697));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747), .A(N30248), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9411), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9603), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2740 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9887), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9505), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8963), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9411), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9603));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2741 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9631), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9241), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8740), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9887), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9465));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2742 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9362), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8870), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9631));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2743 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[22]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8947), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9718));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6596), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5866), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6323), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6052), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5866));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2749 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6415), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6415));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[4]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6596), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6323), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6209));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2752 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[22]), .B(N22989), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[22]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806), .A(N30246), .B(N30240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9029), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751), .A(N30260), .B(N30258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9464), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5993), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5873), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5993));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5873), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6173), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6358), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2764 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2765 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6173), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6358), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6524), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2766 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2767 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10310), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6061), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5958), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6252));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2768 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9173), .A0(N30228), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B1(N30230));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2769 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .S0(N30296));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2770 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9329), .A(N30305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2774 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9972), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9594), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8712), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9479));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2777 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8681), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9996), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9972), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10007), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10203));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2778 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9811), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8681), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9657), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8705));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2779 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9988), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9615), .A(N27102), .B(N27100), .CI(N29448));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9734), .A(N25457), .B(N24248));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2782 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9664), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2786 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .S0(N30296));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2787 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8946), .A(N30305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2788 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9337), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2789 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8986), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10258), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9337));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2790 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9397), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8986), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9234), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9996));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2791 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8832), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9734), .B(N29398), .CI(N29446));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8763), .A(N30232), .B(N24241));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2793 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9008), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8832), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8763), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9615));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2794 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9188), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8826), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9988), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9008));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2795 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9958), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9464), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9173), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8826));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2796 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8938), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10279), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9767), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9029), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9958));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704), .A(N30262), .B(N30260), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2798 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9851), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2799 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2800 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2801 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9151), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8795), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9851), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9188), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10025));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2802 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8905), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10247), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9151), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9735));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2805 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2806 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8853), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2807 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2808 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2809 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9924), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8853), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10200));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2810 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9669), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8765), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9924), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9505));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2811 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8685), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10001), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10211), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8905), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9669));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2812 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[21]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8685), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9970), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8984));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6085), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6015));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6278), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6191));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2818 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6450), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6371));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6118), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6480), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6308), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6118), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6480));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2823 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6085), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6278), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6450), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5899));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2824 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[21]), .B(N22959), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[21]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2825 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2827 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9842), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2828 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409), .A(N30250), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10016), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965), .B(N30228));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805), .A(N30258), .B(N30256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2832 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9076), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2833 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9776), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10149), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8675), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9076));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2834 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9742), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9351), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10016), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9776));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2835 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8743), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10279), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9742), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9543));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2836 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024), .A(N30234), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2837 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9210), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2838 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645), .A(N30248), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2839 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10193), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2840 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2841 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9661), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2842 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8695), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2844 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8974), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10193), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9661), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8695));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2845 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9705), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9315), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8795), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9210), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8974));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2846 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8715), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8743), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9705), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10247));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2847 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[20]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8715), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9241), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10001));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2848 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5972), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5852), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6613));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5883), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6434), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5883), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6434), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6263), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6150));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[2]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5972), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5852), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6341));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2857 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[20]), .B(N22969), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[20]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2858 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2860 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2861 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086), .A(N30238), .B(N30236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2862 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8843), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712), .A(N30246), .B(N30240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9833), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2865 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2867 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932), .A(N30234), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2869 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8800), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10135), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9267), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10010));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2870 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8773), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8843), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8800));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2876 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9094), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2877 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2878 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9897), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2879 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2880 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10041), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2881 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10095), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9730), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9094), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9897), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10041));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2882 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9757), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9364), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9594), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10095), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8658));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8960), .A(N30232), .B(N24250));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2884 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10143), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9784), .A(N29396), .B(N26726), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8960));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2885 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862), .A(N30256), .B(N30254), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8736), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2887 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9589), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10169), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10143), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8736));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2888 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9552), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9160), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9649), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9589));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2889 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9514), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10308), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9552), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9351));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2890 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9473), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9315), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8773), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9514));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2891 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[19]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9473), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9276), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10037));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2893 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6645), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5919));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2894 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6567), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2895 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6104), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6001), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6104));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5839), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2900 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6464), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6327), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5839), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6494));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2901 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6645), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6567), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6001), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6464));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2902 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[19]), .B(N22979), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[19]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2903 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2904 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6354), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2905 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2906 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6055), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5992));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2907 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6454), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6170), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2911 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6090), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6454), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6631), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6170));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2912 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[0]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6055), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6520));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2913 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142), .A(N30236), .B(N30230), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2914 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2915 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2916 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8893), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2919 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993), .A(N30238), .B(N30236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2920 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2921 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8652), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9964), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9448), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8893), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9640));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2922 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10284), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9930), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9389), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10187), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8652));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2923 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310), .A(N30250), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2924 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9071), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544), .A(N30248), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8897), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2931 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2932 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10215), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9858), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8897), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8746));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2933 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9108), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8958), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10215), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9730));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2934 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9949), .A(N30232), .B(N24268));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2935 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8785), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10117), .A(N26744), .B(N26742), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9949));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2936 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923), .A(N30254), .B(N30244), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2937 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2938 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9167), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8806), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9784), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8785), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10060));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2939 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9359), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8980), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9071), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9258), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9167));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2940 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9324), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10135), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9359), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9160));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2941 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10253), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9893), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10284), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9324));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2942 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[18]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10253), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10070), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9087));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2943 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989), .A(N23378), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[18]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12498), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2946 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205), .A(N30230), .B(N30228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2947 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9827), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2948 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837), .A(N30234), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053), .A(N30236), .B(N30230), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9249), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2954 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9936), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9066), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10236), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9249));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2955 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10114), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9198), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9827), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9936));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439), .A(N30248), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2960 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .S0(N30296));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9934), .A(N30305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2963 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9374), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9882), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9934));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507), .S0(N30295));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2965 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10288), .A(N30304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2966 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9243), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9374), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10288), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9858));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2967 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9177), .A(N30232), .B(N24653));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2968 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9884), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9499), .A(N26736), .B(N26734), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9177));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2969 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2970 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10074), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2971 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2972 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9130), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2973 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .S0(N30295));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9557), .A(N30304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2976 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8777), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2978 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10039), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9671), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9557), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9106), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8777));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2979 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10127), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9764), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9130), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10152), .A(N30232), .B(N24633));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2981 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10005), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9633), .A(N27094), .B(N27092), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10152));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046), .A(N30252), .B(N30250), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9300), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2984 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8901), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9499), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10005), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9300));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2985 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9298), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8924), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10052), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10227), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8901));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898), .A(N30238), .B(N30236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8725), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204), .A(N30250), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9879), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2990 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115), .A(N30230), .B(N30228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8879), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2992 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10265), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9879), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8879));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2993 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8752), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10085), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10265), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9562));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2994 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9901), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9750), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8980), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8752));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608), .A(N30246), .B(N30240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8886), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2997 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I2998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8729), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I2999 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8950), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8886), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8729));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9438), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3002 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983), .A(N30244), .B(N30252), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3004 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9529), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9136), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10117), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9884), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9694));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3005 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9722), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9330), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9438), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9529), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8806));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3006 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9131), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9964), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8950), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9722));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3007 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10076), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9714), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10114), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9131));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3008 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[16]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9901), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8943), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9714));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3009 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[17]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9123), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9893));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3010 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[17]));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12310), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[16]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[16]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3012 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12310));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3013 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10091), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .S0(N30295));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9165), .A(N30304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3016 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8968), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10091), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9165));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3017 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3018 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10112), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .S0(N30295));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8804), .A(N30304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10296), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736), .B(N30295));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10138), .A(N30304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3025 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9863), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9476), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10296), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10138));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3026 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9410), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9030), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9336), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9863));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3027 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9737), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9344), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10112), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9410));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3028 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9057), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8717), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9671), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8968), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9737));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3029 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9147), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8791), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9764), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8995), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9057));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104), .A(N24635), .B(N30242), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8928), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3032 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9022), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9633), .B(N29618), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8928));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3033 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020), .A(N30230), .B(N30228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3034 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9678), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3035 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339), .A(N30248), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3036 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804), .A(N30238), .B(N30236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3038 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3039 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9791), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9403), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9678), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9103), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9485));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3040 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9432), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9048), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9022), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9791));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3041 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9074), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8735), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8924), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9910), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9432));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3043 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3044 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961), .A(N30236), .B(N30230), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10046), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3046 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9665), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9494), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10046));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3047 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3048 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3049 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744), .A(N30234), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9870), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508), .A(N30246), .B(N30240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3053 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8713), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10220), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9870), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9686));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3054 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10056), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9136), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8713));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3055 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9492), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9101), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10056), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10290), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9330));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3056 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[14]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10085), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9074), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9101));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3057 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[15]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8780), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9492), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9524));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3058 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[15]));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12410), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[14]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[14]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9405), .A(N30232), .B(N30250));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3061 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170), .A(N30242), .B(N30248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3062 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10268), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3063 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9920), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9536), .A(N29616), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9405), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10268));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3064 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3065 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9293), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3066 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8813), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9920), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9293), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8688));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3067 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10177), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9820), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9269), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8813), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10032));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3068 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[13]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10177), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9691), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8735));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3069 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12104), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[13]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3070 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641), .A(N30234), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868), .A(N30236), .B(N30230), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3073 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9097), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3074 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8691), .A(N30232), .B(N24662));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3075 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240), .A(N24642), .B(N30246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3076 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9912), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3077 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9826), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9440), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8691), .B(N27231), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9912));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3078 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9701), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8921), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9097), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9826));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3079 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406), .A(N30246), .B(N30240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3083 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8932), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10274), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8757), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9285));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3084 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9566), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9701), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8932), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9403));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3085 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[12]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9048), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9820));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3086 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[12]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931), .A(N30230), .B(N30228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3090 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10088), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3091 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708), .A(N30238), .B(N30236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10262), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3093 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8845), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10186), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10088), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10262));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3094 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8741), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8845), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9536), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10274));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3095 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[11]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8741), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10150), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9172));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[11]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3097 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9635), .A(N30232), .B(N24642));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304), .A(N24644), .B(N25288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3099 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3100 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8767), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10104), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9635), .B(N27456), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9532));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542), .A(N30234), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3102 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9725), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10078), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3105 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9510), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9117), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10078));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3106 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9602), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9440), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8767), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9510));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3107 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[10]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[9]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9602), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9308), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10066));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11915), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[10]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3109 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8874), .A(N30232), .B(N30246));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369), .A(N30240), .B(N30234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3112 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10160), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9797), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8874), .B(N27448), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9139));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3113 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770), .A(N30236), .B(N30230), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9903), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3115 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10250), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9889), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10160), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9903), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10104));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3116 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[9]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10186), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10250), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9209));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3117 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12270), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[9]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834), .A(N30230), .B(N30228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3119 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606), .A(N30238), .B(N30236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9334), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9859), .A(N30232), .B(N30240));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436), .A(N25313), .B(N30238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3124 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8786), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3125 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8878), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10222), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9859), .B(N27640), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8786));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3126 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9182), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8819), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9527), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9334), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8878));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3127 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[8]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9117), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9182), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9889));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3128 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11996), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[8]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[8]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3129 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673), .A(N30236), .B(N30230), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3132 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9133), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3133 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9642), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8952), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9133));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3134 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[7]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9642), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9797), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8819));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12350), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[7]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3136 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9084), .A(N30232), .B(N30234));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3137 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9564), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3138 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504), .A(N25295), .B(N25297), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3139 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10122), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3140 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10072), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9710), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9084), .B(N27844), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10122));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10069), .A(N30232), .B(N30238));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3142 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570), .A(N30236), .B(N25852), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3144 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10281), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10069), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9759));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741), .A(N30230), .B(N30228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N30224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3147 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9090), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10292), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9710));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3148 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[6]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10222), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10072), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9090));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3149 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12069), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[6]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3150 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[5]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3151 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3152 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9942), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545), .B(N29556), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9311), .A(N30232), .B(N30236));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637), .A(N25852), .B(N25854), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9366), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3156 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9546), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9366));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3157 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[4]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9942), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9546));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3158 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[4]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3159 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[3]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10277), .A(N30232), .B(N30230));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3161 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[2]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10277), .B(N30226));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[2]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704), .A(N30228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3165 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12278), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[1]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[1]));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3166 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12112), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12230), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12278), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[2]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[2]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[3]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3168 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11958), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12509), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12112), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12376));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3169 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12346), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12151), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11958), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[4]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[4]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[5]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3171 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12101), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12432), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12346), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12291));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12421), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12069), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12101), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[6]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[6]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[7]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12083), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12350), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12421), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12207));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12320), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11996), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12083), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[8]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[8]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[9]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11920), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12270), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12320), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12128));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12061), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11915), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11920), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[10]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[10]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[11]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3180 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12210), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12185), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12061), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12052));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12281), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12467), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12210), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[12]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[12]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[13]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3183 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12348), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12104), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12281), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11973));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3184 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[14]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3185 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12519), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[15]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3186 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12266), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12243), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12519));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12250), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12410), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12348), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12266));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[16]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12444), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[17]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12169), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12161), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12444));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12014), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12169), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[18]), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12192), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12148), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12250), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12014));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12498), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12192), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3196 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3197 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3198 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3200 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3201 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3202 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3203 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3204 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3205 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3206 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3207 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3208 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3210 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3211 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3212 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3213 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3215 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3217 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3218 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3219 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3224 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3225 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3226 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3227 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182), .A(N29502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464), .A(N22618), .B(N29506));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3232 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3233 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3234 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3235 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3236 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3237 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3238 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3239 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3240 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3241 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12415), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3242 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3243 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12246), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12302), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391), .A1(N29510), .B0(N21795));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3248 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12356), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12302));
AOI31X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3249 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127), .A2(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12356));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3251 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3252 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107), .A(N29679), .B(N29681));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156), .A(N22305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3255 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273), .A(N21999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3256 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3257 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3260 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3261 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3262 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3263 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3264 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3265 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3266 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3269 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3270 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3271 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3276 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3277 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3278 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3279 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3280 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3281 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3282 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3283 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3287 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3289 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3290 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3291 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024), .A0(N22305), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464), .B0(N22309));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3296 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131), .A0(N21999), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024), .B0(N22003));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3297 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3298 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12418), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3299 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11976), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12418));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3300 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12030), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131), .B0(N20660));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3301 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12076), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12030));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3302 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12133), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12217), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12076));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[48]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12133), .B(N20538));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(N20492), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[48]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3305 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219), .B(N18660));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3306 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470), .A(N29667), .B(N29669));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999), .A(N21993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3310 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3311 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3312 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3314 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3315 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3316 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3319 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3320 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3321 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3322 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3323 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492), .A0(N21993), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383), .B0(N21988));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3325 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12328), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3326 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12387), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492), .B0(N21782));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3327 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12440), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12387));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3328 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12494), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11945), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12440));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3329 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11901), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3330 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[47]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12494), .B(N21075));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[47]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242), .A(N21765), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3335 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3336 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3338 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12299), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3344 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3349 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3350 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12055), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12103), .A0(N21765), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211), .B0(N21769));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12157), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12103));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3354 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12213), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12299), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12157));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3355 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12115), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[46]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12213), .B(N21090));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3357 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[46]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3358 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3359 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972), .A(N29566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3361 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12027), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3362 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3363 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3364 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3365 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12466), .A0(N29566), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941), .B0(N29510));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12516), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12466));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11943), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12027), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12516));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12335), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[45]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11943), .B(N21080));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[45]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3372 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12384), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3378 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3379 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12184), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12239), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12184));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3381 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12297), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12384), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12239));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11927), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[44]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12297), .B(N21085));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3384 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[44]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3385 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3386 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3387 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3388 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3389 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12100), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3390 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3392 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11914), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11969), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11914));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12023), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12100), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11969));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3395 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12138), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[43]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12023), .B(N21070));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[43]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12463), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12269), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3404 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12322), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12269));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3405 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12382), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12463), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12322));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3406 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12362), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3407 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[42]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12382), .B(N21100));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[42]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12047), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12097), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12181), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12047));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11950), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[41]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12097), .B(N21105));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[41]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11911), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3417 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12407), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12459), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11911), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12407));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3419 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12163), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[40]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12459), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12163));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[40]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3423 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3424 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3425 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3426 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12125), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3427 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12179), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12263), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12125));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12390), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[39]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12179), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12390));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[39]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3432 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12484), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11909), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11992), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12484));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11975), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[38]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11975));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3436 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[38]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3438 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3439 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12203), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12260), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12345), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12203));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12187), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3442 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[37]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12260), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12187));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3443 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[37]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3444 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3445 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11935), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3446 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11990), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12065), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11935));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3447 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12414), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3448 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[36]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12414));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[36]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12264), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11998), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[35]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12264), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11998));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[35]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3456 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12124), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12209), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[34]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12124), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12209));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[34]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3460 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12434), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[33]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12434));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[33]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3464 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12020), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[32]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12020));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3466 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[32]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3467 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3471 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12232), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3472 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12232));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3473 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[31]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3474 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12456), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[30]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12456));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[30]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12042), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3479 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12042));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3480 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[29]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3481 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12257), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12257));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3483 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[28]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3484 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3485 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3486 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13351), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13387), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13406), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13351), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13387));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3489 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13347), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3490 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13406), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13347));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12478), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[27]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12478));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[27]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12060), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3495 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12060));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[26]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3498 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13349), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13367), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13397), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13349));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3500 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13359), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3501 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3502 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13392), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13359), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13375));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3503 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13339), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13367), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13392));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3504 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13383), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3505 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13374), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13383), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3506 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13339), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13374));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12284), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12284));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[25]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3510 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13340), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3511 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3512 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13393), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13340), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13376));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13384), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13337), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13384), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13402));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3516 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13379), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13393), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13337));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13409), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13343), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13362), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13409), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13343));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13352), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3521 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13388), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13352), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13368));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3523 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13334), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13362), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13388));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13360), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13379), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13334));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13377), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13395), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13332), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13377), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13395));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13404), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13398), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13358), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13404), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13398));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13394), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13332), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13358));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13394));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3533 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13475), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13475), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13472), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[0]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3540 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3541 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3542 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[0]));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3543 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3550 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13492), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13540), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13492), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13490), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13540), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13591), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13490), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0]));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N701), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13591), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N670), .A0(N30278), .A1(N18886), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N701));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13185), .A(a_exp[7]), .B(a_exp[0]));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13187), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19047), .A(a_exp[6]), .B(a_exp[5]), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13187));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13185), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19047));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3576 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19054));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13221), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3578 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13225), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13221));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13208), .A(a_man[10]), .B(a_man[9]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13227), .A(a_man[6]), .B(a_man[5]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13216), .A(a_man[8]), .B(a_man[7]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13236), .A(N30313), .B(a_man[3]));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13227), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13216), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13236));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13230), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13240), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3586 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__24), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13219), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13230), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13240));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__24));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13288), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13292), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__17), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13292));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__17), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N670), .B(N30270), .S0(N30273));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3594 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3595 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3596 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3599 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3600 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13511), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13612), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3604 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3605 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13610), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13511), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13558), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13610), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N700), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13558), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669), .A0(N30281), .A1(N18971), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N700));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669), .B(N30270), .S0(N30272));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3619 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3621 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3622 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13628), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13576), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13628), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13522), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13576), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N699), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13522), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668), .A0(N30279), .A1(N19020), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N699));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668), .B(N30270), .S0(N30273));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13596), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13539), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13596), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13491), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13539), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N698), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13491), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667), .A0(N30282), .A1(N19000), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N698));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3645 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667), .B(N30270), .S0(N30276));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13510), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13611), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13510), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N697), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13611), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666), .A0(N30282), .A1(N19030), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N697));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666), .B(N30270), .S0(N30274));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13627), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3656 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13578), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13627), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N696), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13578), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665), .A0(N30279), .A1(N19010), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N696));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665), .B(N30270), .S0(N30275));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13595), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13542), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13595), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3665 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3666 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N695), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13542), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664), .A0(N30281), .A1(N18990), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N695));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664), .B(N30270), .S0(N30274));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13562), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13513), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13562), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3673 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13513));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663), .A0(N30283), .A1(N19040), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N694));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663), .B(N30270), .S0(N30275));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13630), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13630));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662), .A0(N30278), .A1(N19050), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N693));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662), .B(N30270), .S0(N30274));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13597), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13597));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661), .A0(N30280), .A1(N19099), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N692));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661), .B(N30270), .S0(N30275));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3684 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13564), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3685 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13564));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3686 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660), .A0(N30278), .A1(N19109), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N691));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3687 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660), .B(N30270), .S0(N30272));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13528), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13528));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659), .A0(N30284), .A1(N19119), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N690));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659), .B(N30270), .S0(N30272));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13498), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N689), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13498));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658), .A0(N30278), .A1(N19149), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N689));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658), .B(N30270), .S0(N30275));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13618), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13618));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657), .A0(N30280), .A1(N19060), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N688));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[9]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657), .B(N30270), .S0(N30274));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13584), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3701 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13584));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3702 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656), .A0(N30283), .A1(N19129), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N687));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656), .B(N30270), .S0(N30272));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3704 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13588));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655), .A0(N30280), .A1(N19159), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N686));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655), .B(N30270), .S0(N30273));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N685), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654), .A0(N30283), .A1(N19139), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N685));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654), .B(N30270), .S0(N30276));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N684), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653), .A0(N30282), .A1(N19070), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N684));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653), .B(N30270), .S0(N30273));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652), .A0(N30281), .A1(N19080), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N683));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652), .B(N30270), .S0(N30273));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N682), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651), .A0(N30282), .A1(N19233), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N682));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651), .B(N30270), .S0(N30276));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N681), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650), .A0(N30281), .A1(N19223), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N681));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650), .B(N30270), .S0(N30275));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3723 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3724 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649), .A0(N30280), .A1(N19275), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N680));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649), .B(N30270), .S0(N30274));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648), .A0(N30279), .A1(N19410), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N679));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[0]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648), .B(N30270), .S0(N30272));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647), .A(a_exp[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14019), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14019));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[30]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .AN(N30278), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13863), .A0(N20175), .A1(N30281), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13863));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646), .B(N18839), .S0(N18835));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13818), .A0(N20182), .A1(N30280), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13818));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3740 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645), .B(N18839), .S0(N18835));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13877), .A0(N19891), .A1(N30283), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13877));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[27]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644), .B(N18839), .S0(N18835));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13832), .A0(N19768), .A1(N30283), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13832));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643), .B(N18839), .S0(N18835));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13786), .A0(N19900), .A1(N30279), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13786));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3749 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642), .B(N18839), .S0(N18835));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13845), .A0(N19909), .A1(N30279), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13845));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641), .B(N18839), .S0(N18835));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13800), .A0(N20144), .A1(N30282), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13800));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[23]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640), .B(N18839), .S0(N18835));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5424));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N577), .A(a_sign), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N757));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13947), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13940), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13947), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3764 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13925), .A(N19633), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3765 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3766 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13969), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3767 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13939), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13957), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13969));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3768 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13939), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3769 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13934), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13955), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3770 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N578), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13943), .C(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13940), .D(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13934));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_4_I3771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N579), .AN(N18881), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N578), .C(N18678), .D(N18879));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_4_I3772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N579), .B(N18664), .S0(N30284));
reg x_reg_L0_30__I3803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_30__I3803_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[30];
	end
assign N9100 = x_reg_L0_30__I3803_QOUT;
reg x_reg_L1_0__I3805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__I3805_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[0];
	end
assign x[0] = x_reg_L1_0__I3805_QOUT;
reg x_reg_L1_1__I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__I3806_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[1];
	end
assign x[1] = x_reg_L1_1__I3806_QOUT;
reg x_reg_L1_2__I3807_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__I3807_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[2];
	end
assign x[2] = x_reg_L1_2__I3807_QOUT;
reg x_reg_L1_3__I3808_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__I3808_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[3];
	end
assign x[3] = x_reg_L1_3__I3808_QOUT;
reg x_reg_L1_4__I3809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__I3809_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[4];
	end
assign x[4] = x_reg_L1_4__I3809_QOUT;
reg x_reg_L1_5__I3810_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__I3810_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[5];
	end
assign x[5] = x_reg_L1_5__I3810_QOUT;
reg x_reg_L1_6__I3811_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__I3811_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[6];
	end
assign x[6] = x_reg_L1_6__I3811_QOUT;
reg x_reg_L1_7__I3812_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__I3812_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[7];
	end
assign x[7] = x_reg_L1_7__I3812_QOUT;
reg x_reg_L1_8__I3813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__I3813_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[8];
	end
assign x[8] = x_reg_L1_8__I3813_QOUT;
reg x_reg_L1_9__I3814_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__I3814_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[9];
	end
assign x[9] = x_reg_L1_9__I3814_QOUT;
reg x_reg_L1_10__I3815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__I3815_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[10];
	end
assign x[10] = x_reg_L1_10__I3815_QOUT;
reg x_reg_L1_11__I3816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__I3816_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[11];
	end
assign x[11] = x_reg_L1_11__I3816_QOUT;
reg x_reg_L1_12__I3817_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__I3817_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[12];
	end
assign x[12] = x_reg_L1_12__I3817_QOUT;
reg x_reg_L1_13__I3818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__I3818_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[13];
	end
assign x[13] = x_reg_L1_13__I3818_QOUT;
reg x_reg_L1_14__I3819_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__I3819_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[14];
	end
assign x[14] = x_reg_L1_14__I3819_QOUT;
reg x_reg_L1_15__I3820_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__I3820_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[15];
	end
assign x[15] = x_reg_L1_15__I3820_QOUT;
reg x_reg_L1_16__I3821_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__I3821_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[16];
	end
assign x[16] = x_reg_L1_16__I3821_QOUT;
reg x_reg_L1_17__I3822_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__I3822_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[17];
	end
assign x[17] = x_reg_L1_17__I3822_QOUT;
reg x_reg_L1_18__I3823_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__I3823_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[18];
	end
assign x[18] = x_reg_L1_18__I3823_QOUT;
reg x_reg_L1_19__I3824_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__I3824_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[19];
	end
assign x[19] = x_reg_L1_19__I3824_QOUT;
reg x_reg_L1_20__I3825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__I3825_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[20];
	end
assign x[20] = x_reg_L1_20__I3825_QOUT;
reg x_reg_L1_21__I3826_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__I3826_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[21];
	end
assign x[21] = x_reg_L1_21__I3826_QOUT;
reg x_reg_L1_22__I3827_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__I3827_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[22];
	end
assign x[22] = x_reg_L1_22__I3827_QOUT;
reg x_reg_L1_23__I3828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__I3828_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[23];
	end
assign x[23] = x_reg_L1_23__I3828_QOUT;
reg x_reg_L1_24__I3829_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__I3829_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[24];
	end
assign x[24] = x_reg_L1_24__I3829_QOUT;
reg x_reg_L1_25__I3830_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__I3830_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[25];
	end
assign x[25] = x_reg_L1_25__I3830_QOUT;
reg x_reg_L1_26__I3831_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__I3831_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[26];
	end
assign x[26] = x_reg_L1_26__I3831_QOUT;
reg x_reg_L1_27__I3832_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__I3832_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[27];
	end
assign x[27] = x_reg_L1_27__I3832_QOUT;
reg x_reg_L1_28__I3833_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__I3833_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[28];
	end
assign x[28] = x_reg_L1_28__I3833_QOUT;
reg x_reg_L1_29__I3834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__I3834_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[29];
	end
assign x[29] = x_reg_L1_29__I3834_QOUT;
reg x_reg_L1_30__I3835_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__I3835_QOUT <= N9100;
	end
assign x[30] = x_reg_L1_30__I3835_QOUT;
reg x_reg_L1_31__I3836_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I3836_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[31];
	end
assign x[31] = x_reg_L1_31__I3836_QOUT;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[29] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[49] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[30] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[4] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urX4TwjdoxhI : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



