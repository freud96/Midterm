/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:53 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42;
wire [22:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82;
wire [0:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195;
wire [20:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197;
wire [32:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5398,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5406,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5409,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5411,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5476,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5499,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5501,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5654,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5726,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5766,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5795,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5815,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5818,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5825,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5842,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5857,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5876,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5889,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5895,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5905,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5907,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5912,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6007,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6026,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6027,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6049,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6051,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6064,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6085,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6193,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6248,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7127,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7217,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7297,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7347,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7726,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7762,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7790,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7793,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7809,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7815,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7855,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7857,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7860,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7861,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7868,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7873,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7877,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7882,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7883,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7894,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7896,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7898,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7930,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7942,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7974,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7997,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7998,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8003,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8019,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8026,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8027,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8048,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8053,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8064,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8071,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8112,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8127,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8135,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8141,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8167,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8282,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8297,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8300,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8323,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8340,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8342,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8348,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8358,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8360,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8372,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8381,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8428,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8444,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8455,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8537,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8546,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8559,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8581,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8597,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8762,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9912,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9930,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9933,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9942,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9995,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9996,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9997,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10002,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10015,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10017,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10031,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10032,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10041,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10049,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10051,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10077,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10085,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10094,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10106,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10112,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10117,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10122,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10127,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10137,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10149,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10286,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10312,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10318,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10342,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10343,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10347,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10348,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10359,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10372,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10374,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10380,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10381,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10382,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10384,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10387,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10409,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10423,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10465,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10476,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10496,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10500,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10518,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11193,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11217,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11268,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11272,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11312,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11332,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11340,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11342,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11343,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11360,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11378,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11382,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11387,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11398,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11407,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11411,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11415,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11428,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11429,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11462,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11465,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11476,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11499,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11500,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11501,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11559,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11654,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11762,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11790,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11793,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11795,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11809,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11825,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11828,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11836,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11850,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11853,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11861,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11868,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11873,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11877,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11879,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11880,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11889,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11892,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11894,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11895,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11896,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11897,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11901,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11995,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11998,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12013,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12018,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12026,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12030,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12051,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12053,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12060,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12064,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12071,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12073,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12085,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12094,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12114,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12122,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12137,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12149,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12167,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12250,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12259,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12274,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12279,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12286,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12296,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12297,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12300,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12318,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12323,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12340,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12343,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12348,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12358,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12360,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12374,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12375,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12381,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12382,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12384,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12392,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12398,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12406,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12407,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12415,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12423,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12428,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12444,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12455,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12462,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12465,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12496,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12499,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12515,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12518,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12537,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12548,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12559,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12581,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12597,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12604,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12793,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12815,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12822,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12825,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12842,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12857,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12860,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12864,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12866,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12868,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14515,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14537,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14604,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14795,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14822,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14853,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14877,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14882,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14896,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14974,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15031,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15041,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15048,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15057,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15790,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15898,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43268,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43853,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43894,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43997,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44049,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44095,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44122,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44129;
wire N19976,N19980,N19983,N19994,N19998,N20199,N20253 
	,N20260,N20350,N20360,N20370,N20392,N20414,N20424,N20434 
	,N20444,N20454,N20471,N20481,N20491,N20501,N20537,N20547 
	,N20557,N20567,N20577,N20587,N20597,N20607,N20617,N20988 
	,N21042,N21116,N21208,N21231,N21450,N21461,N21468,N21766 
	,N21801,N22304,N22319,N22330,N22332,N22342,N22344,N22349 
	,N22351,N22356,N22358,N22361,N22366,N22368,N22373,N22378 
	,N22385,N22387,N22392,N22395,N22397,N22402,N22404,N22409 
	,N22411,N22416,N22421,N22423,N22430,N22432,N22437,N22439 
	,N22442,N22444,N22451,N22453,N22482,N22484,N22489,N22504 
	,N22508,N22510,N22512,N22516,N22518,N22520,N22524,N22526 
	,N22528,N22531,N22534,N22536,N22558,N22562,N22564,N22566 
	,N22569,N22571,N22581,N22583,N22593,N22598,N22600,N22644 
	,N22646,N22648,N23029,N23056,N23313,N23314,N23315,N23316 
	,N23317,N23318,N23319,N23320,N23321,N23322,N23323,N23324 
	,N23325,N23326,N23327,N23328,N23329,N23330,N23331,N23332 
	,N23333,N23334,N23335,N23336;
EDFFHQX1 x_reg_31__retimed_I13794 (.Q(N23056), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14990), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13781 (.Q(N23029), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43441), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13653 (.Q(N22648), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14700), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13652 (.Q(N22646), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14649), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13651 (.Q(N22644), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14896), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13631 (.Q(N22600), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13630 (.Q(N22598), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14959), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13628 (.Q(N22593), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14822), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13625 (.Q(N22583), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13624 (.Q(N22581), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14888), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13620 (.Q(N22571), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13619 (.Q(N22569), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14644), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13618 (.Q(N22566), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14783), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13617 (.Q(N22564), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13616 (.Q(N22562), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13615 (.Q(N22558), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14830), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13608 (.Q(N22536), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14655), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13607 (.Q(N22534), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15006), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13606 (.Q(N22531), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14634), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13605 (.Q(N22528), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13604 (.Q(N22526), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13603 (.Q(N22524), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13602 (.Q(N22520), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14537), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13601 (.Q(N22518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13600 (.Q(N22516), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13599 (.Q(N22512), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15039), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13598 (.Q(N22510), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14610), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13597 (.Q(N22508), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13596 (.Q(N22504), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14951), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13591 (.Q(N22489), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14787), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13589 (.Q(N22484), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14980), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13588 (.Q(N22482), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14859), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13586 (.Q(N22453), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15014), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13585 (.Q(N22451), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14564), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13582 (.Q(N22444), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14652), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13581 (.Q(N22442), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14525), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13580 (.Q(N22439), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14619), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13579 (.Q(N22437), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14739), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13577 (.Q(N22432), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14877), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13576 (.Q(N22430), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15000), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13573 (.Q(N22423), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15024), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13572 (.Q(N22421), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14899), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13570 (.Q(N22416), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14571), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13568 (.Q(N22411), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14958), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13567 (.Q(N22409), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14840), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13565 (.Q(N22404), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14589), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13564 (.Q(N22402), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15038), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13562 (.Q(N22397), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14782), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13561 (.Q(N22395), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14665), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13560 (.Q(N22392), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14669), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13558 (.Q(N22387), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14703), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13557 (.Q(N22385), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14826), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13554 (.Q(N22378), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14964), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13552 (.Q(N22373), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43811), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13550 (.Q(N22368), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14760), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13549 (.Q(N22366), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14643), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13547 (.Q(N22361), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14528), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13546 (.Q(N22358), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15079), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13545 (.Q(N22356), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14630), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13543 (.Q(N22351), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43804), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13542 (.Q(N22349), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43800), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13540 (.Q(N22344), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15061), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13539 (.Q(N22342), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14609), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13535 (.Q(N22332), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43432), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13534 (.Q(N22330), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43446), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13531 (.Q(N22319), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14881), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13526 (.Q(N22304), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14614), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13362 (.Q(N21801), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14543), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13349 (.Q(N21766), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13270 (.Q(N21468), .D(a_exp[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13267 (.Q(N21461), .D(a_exp[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13262 (.Q(N21450), .D(a_exp[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13187 (.Q(N21231), .D(a_exp[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13177 (.Q(N21208), .D(a_exp[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13151 (.Q(N21116), .D(a_exp[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13120 (.Q(N21042), .D(a_exp[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I13108 (.Q(N20988), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12961 (.Q(N20617), .D(a_man[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12957 (.Q(N20607), .D(a_man[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12953 (.Q(N20597), .D(a_man[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12949 (.Q(N20587), .D(a_man[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12945 (.Q(N20577), .D(a_man[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12941 (.Q(N20567), .D(a_man[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12937 (.Q(N20557), .D(a_man[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12933 (.Q(N20547), .D(a_man[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12929 (.Q(N20537), .D(a_man[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12914 (.Q(N20501), .D(a_man[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12910 (.Q(N20491), .D(a_man[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12906 (.Q(N20481), .D(a_man[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12902 (.Q(N20471), .D(a_man[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12895 (.Q(N20454), .D(a_man[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12891 (.Q(N20444), .D(a_man[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12887 (.Q(N20434), .D(a_man[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12883 (.Q(N20424), .D(a_man[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12879 (.Q(N20414), .D(a_man[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12870 (.Q(N20392), .D(a_man[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12861 (.Q(N20370), .D(a_man[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12857 (.Q(N20360), .D(a_man[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12853 (.Q(N20350), .D(a_man[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12816 (.Q(N20260), .D(a_man[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I12813 (.Q(N20253), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16612), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_26__retimed_I12789 (.Q(N20199), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I12700 (.Q(N19998), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I13923 (.Y(N23313), .A(N19998));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13929 (.Y(N23319), .A(N23313));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13928 (.Y(N23318), .A(N23313));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13927 (.Y(N23317), .A(N23313));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13926 (.Y(N23316), .A(N23313));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13925 (.Y(N23315), .A(N23313));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13924 (.Y(N23314), .A(N23313));
EDFFHQX1 x_reg_22__retimed_I12698 (.Q(N19994), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I13930 (.Y(N23320), .A(N19994));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13936 (.Y(N23326), .A(N23320));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13935 (.Y(N23325), .A(N23320));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13934 (.Y(N23324), .A(N23320));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13933 (.Y(N23323), .A(N23320));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13932 (.Y(N23322), .A(N23320));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13931 (.Y(N23321), .A(N23320));
EDFFHQX1 x_reg_20__retimed_I12693 (.Q(N19983), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I13937 (.Y(N23327), .A(N19983));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13938 (.Y(N23328), .A(N23327));
EDFFHQX1 x_reg_31__retimed_I12692 (.Q(N19980), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I13939 (.Y(N23329), .A(N19980));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13946 (.Y(N23336), .A(N23329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13945 (.Y(N23335), .A(N23329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13944 (.Y(N23334), .A(N23329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13943 (.Y(N23333), .A(N23329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13942 (.Y(N23332), .A(N23329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13941 (.Y(N23331), .A(N23329));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13940 (.Y(N23330), .A(N23329));
EDFFHQX1 x_reg_31__retimed_I12690 (.Q(N19976), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829), .E(bdw_enable), .CK(aclk));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I0 (.Y(bdw_enable), .A(astall));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15746), .A(a_exp[6]), .B(a_exp[5]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749), .A(a_exp[4]), .B(a_exp[3]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15737), .A(a_exp[2]), .B(a_exp[1]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15737));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I5 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22738), .A(a_exp[7]), .B(a_exp[0]), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15744));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I6 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15746), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22738));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I7 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15854), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I8 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15854));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I9 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15839), .A(a_sign), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I10 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829), .A(a_sign));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I11 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15832), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I12 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15798), .A(a_man[4]), .B(a_man[3]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I13 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15767), .A(a_man[10]), .B(a_man[9]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I14 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15777), .A(a_man[8]), .B(a_man[7]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I15 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15788), .A(a_man[6]), .B(a_man[5]));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I16 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15798), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15767), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15777), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15788));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I17 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956), .A(a_man[2]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I18 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15790), .A(a_man[0]), .B(a_man[1]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I19 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15790));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I20 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053), .A(a_man[22]), .B(a_man[21]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I21 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15763), .A(a_man[20]), .B(a_man[19]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I22 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15804), .A(a_man[12]), .B(a_man[11]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I23 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15773), .A(a_man[18]), .B(a_man[17]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I24 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15784), .A(a_man[16]), .B(a_man[15]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I25 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15794), .A(a_man[14]), .B(a_man[13]));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I26 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15796), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15773), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15784), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15794));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I27 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15763), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15796));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I28 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15771), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22746));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I29 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__24), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15780), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15769));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I30 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15839), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15832), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__24));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I31 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15863), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I32 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15867), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I33 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__17), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15863), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15867));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I34 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__17), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I35 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I36 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I37 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15898), .A(a_exp[5]), .B(a_exp[6]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I38 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15891), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15898));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I39 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639), .A(a_exp[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15891));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I40 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100), .A(a_exp[2]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I41 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103), .A(a_exp[1]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I42 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107), .A(a_exp[3]));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I43 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I44 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44070), .A(a_exp[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I45 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .A(a_exp[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44070));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I46 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103));
XOR2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I47 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7108));
XOR2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I48 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .A(a_exp[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I49 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236), .A(a_man[22]), .B(a_man[21]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I50 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I51 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .A(a_man[21]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I52 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177), .A(a_man[20]), .B(a_man[22]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I53 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I54 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802), .A(a_man[19]), .B(a_man[21]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I55 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I56 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I57 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5821), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I58 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816), .A(a_man[20]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I59 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5454), .A(a_man[12]), .B(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I60 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5406), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6083), .A(a_man[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5454));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I61 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5912), .A(a_man[14]), .B(a_man[16]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I62 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6211), .A(a_man[13]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I63 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5773), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .B(a_man[19]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6211));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I64 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5406), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5912), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5587));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I65 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5798), .A(a_man[15]), .B(a_man[17]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I66 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6103), .A(a_man[14]), .B(a_man[16]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I67 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703), .A(a_man[22]));
BUFX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I68 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I69 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6155), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6103), .B(a_man[20]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I70 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5773), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5798), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5966));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I71 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I72 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .A(a_man[19]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I73 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5944), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5748), .A(a_man[13]), .B(a_man[11]), .CI(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I74 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5887), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .B(a_man[17]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5944));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I75 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6028), .A(a_man[13]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I76 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5887), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6028), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6083));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I77 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I78 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I79 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541), .A(a_man[17]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I80 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5558), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I81 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .A(a_man[18]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I82 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6059), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5862), .A(a_man[12]), .B(a_man[10]), .CI(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I83 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5507), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5558), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6059));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I84 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6132), .A(a_man[12]), .B(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I85 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6132), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5699));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I86 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I87 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6163), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5975), .A(a_man[11]), .B(a_man[9]), .CI(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I88 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6004), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5810), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6243), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6163), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5862));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I89 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6185), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5748), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6004));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I90 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I91 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I92 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I93 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6051), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5854), .A(a_man[19]), .B(a_man[17]), .CI(a_man[22]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I94 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427), .A(a_man[20]), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6051));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I95 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I96 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040), .A(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I97 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5668), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5476), .A(a_man[21]), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I98 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5668), .B(a_man[16]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5854));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I99 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I100 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5992), .A(a_man[15]), .B(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I102 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5992), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6155));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I105 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5951), .A(a_man[22]), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I109 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5676), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5951), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659), .A(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I111 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5414), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6090), .A(a_man[13]), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5754), .A(a_man[22]), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I113 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5571), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6252), .A(a_man[7]), .B(a_man[21]), .CI(a_man[9]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I114 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5783), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5595), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5754), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5571), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I115 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5621), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5414), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5783));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I116 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5810), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5676), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5621));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I117 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147), .A(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I119 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5514), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6193), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I120 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5683), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5491), .A(a_man[6]), .B(a_man[20]), .CI(a_man[8]));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761), .A(a_man[13]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I122 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6064), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761), .B(a_man[11]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I123 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5895), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5708), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6064), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6252));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I124 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6115), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6090), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5514), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5895));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I125 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5485), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6115));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I126 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I127 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I128 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399), .A(a_man[12]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I129 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6173), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5985), .A(a_man[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I130 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5627), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5441), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6173));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I131 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5792), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5605), .A(a_man[5]), .B(a_man[19]), .CI(a_man[7]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I132 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6011), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5818), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5872), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5792), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5491));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I133 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5727), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6193), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6011));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I134 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5595), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5921));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I136 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878), .A(a_man[11]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I137 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5421), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6097), .A(a_man[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I138 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5736), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5544), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5421), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I139 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5905), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5715), .A(a_man[4]), .B(a_man[18]), .CI(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I140 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6123), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5905), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5985), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5605));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I141 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6221), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5441), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5736), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6123));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I142 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5708), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6221), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5535));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735));
CLKINVX8 DFT_compute_cynw_cm_float_sin_E8_M23_1_I147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496), .A(a_man[10]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I148 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5522), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43881), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I149 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5847), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5661), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5522), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I150 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6021), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43852), .A(a_man[3]), .B(a_man[17]), .CI(a_man[5]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I151 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6227), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6043), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6097), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6021), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5715));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I152 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5842), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5654), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5544), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5847), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6227));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I153 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5818), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6036));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I155 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43875), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43862), .A(a_man[2]), .B(a_man[16]), .CI(a_man[4]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I156 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5957), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43884), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43875));
CLKINVX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I157 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993), .A(a_man[9]));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I158 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43837), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43890), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I159 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5468), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43846), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43837), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43881), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43852));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I160 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5460), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6143), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5957), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5468));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I161 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5460), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5929), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5654));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5478), .A(a_man[22]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I165 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6237), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6054), .A(a_man[3]), .B(a_man[1]), .CI(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I166 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43841), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43894), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6237));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612), .A(a_man[8]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I168 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43845), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43831), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I169 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43870), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43862), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43845), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43890));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I170 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5953), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43841), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43884), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43870));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I171 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5953), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6043), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6143));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I173 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5969), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5775), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040));
ADDFHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I174 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6085), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5889), .A(a_man[14]), .B(a_man[21]), .CI(a_man[0]));
CLKINVX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105), .A(a_man[7]));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I176 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5590), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5408), .A(a_man[5]), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I177 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43849), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43834), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5969), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6085), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5590));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6156), .A(a_man[22]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I179 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43878), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5499), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6156), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6054), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43831));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I180 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43853), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43838), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43894), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43849), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43878));
ADDFHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I181 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43846), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43853), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43867));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I183 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494));
NOR2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I184 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I185 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5700), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I186 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5434), .A(a_man[20]), .B(a_man[13]));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760), .A(a_man[6]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I188 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6188), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43488), .A(a_man[4]), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I189 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43859), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5434), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6188));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I190 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43887), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5775), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5889));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I191 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43891), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43859), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43834), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43887));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I192 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43891), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43838));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43473), .A(a_man[20]), .B(a_man[13]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I195 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5914), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43482), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43473), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43517), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43488));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I196 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43526), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43511), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I197 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5656), .A(a_man[19]), .B(a_man[12]));
CLKINVX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I198 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212), .A(a_man[5]));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I199 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43498), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43481), .A(a_man[3]), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I200 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5530), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43526), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5656), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43498));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I201 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5685), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5493), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5530), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6108));
ADDFHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I202 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5685), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5499), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5874));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I203 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I204 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I205 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5990), .A(a_man[17]), .B(a_man[10]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I206 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5397), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I207 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43485), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5397));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I208 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5758), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5574), .A(a_man[11]), .B(a_man[18]), .CI(a_man[2]));
CLKINVX8 DFT_compute_cynw_cm_float_sin_E8_M23_1_I209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833), .A(a_man[4]));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I210 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6145), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I211 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43477), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5758), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6145));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I212 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551), .A(a_man[3]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I213 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5876), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I214 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43514), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5876), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5955));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I215 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43489), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43474), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43485), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43530), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43514));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43467), .A(a_man[19]), .B(a_man[12]));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I217 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43506), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43492), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43511), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43467), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43481));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I218 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6174), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43477), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43506), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43520));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I219 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43482), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43489), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43503));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I220 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6174), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5614), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5493));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102));
NOR2X6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I224 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I225 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I226 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6222), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906));
CLKINVX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I227 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560), .A(a_man[1]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I228 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5726), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I229 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5702), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5510), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580), .A(a_man[0]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5840), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I232 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6086), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5890), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5840), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I233 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5702), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5890));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I234 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6113), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5919), .A(a_man[0]), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I235 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5620), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5431), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I236 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5591), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5409), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5431), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5726), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I237 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5919), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5409));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I238 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5505), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I239 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6001), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5808), .A(a_man[1]), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I240 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5970), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5779), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6113), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5620), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5808));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I241 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5591), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6183), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5779));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I242 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I243 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6020), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5651), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I245 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6189), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761), .B(a_man[4]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I246 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5651), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6189), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5510));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I248 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5813), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5624), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399), .B(a_man[3]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I249 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5436), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6120), .A(a_man[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612));
BUFX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I251 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5436), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5624));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I252 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6007), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5813), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I255 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5924), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5731), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I256 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5538), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6225), .A(a_man[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I257 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5731), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5538), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I258 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5924), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I260 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6153), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I261 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6153));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I262 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I263 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I264 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5577), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I265 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I266 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5398), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I269 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I270 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I271 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6176), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5467), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6026), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6148));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6042), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I276 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6068), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5660), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6042));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I277 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5730), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5398), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6176), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6068));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I278 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I279 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5778), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5734), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5730), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5542));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I280 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5658), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5464), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I281 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5464), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I282 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6039), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5845), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I283 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5845), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5658), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5857), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5928), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I287 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5439), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5671), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5928), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5439));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I289 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5606), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5778), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5857), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5671));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I290 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6225));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I291 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420));
CLKAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6010));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5817), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I296 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6192));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I297 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5503), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5817), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44036));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I298 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6081), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5606), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5692), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5503));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I299 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5707), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I300 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6089), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I301 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5965), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5707), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6089));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I302 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5594), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5852), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5594), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5973));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I305 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5786), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5965), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5852));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I306 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5540), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5976), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6081), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5786));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5936), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6121), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5540), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5927));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5438), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I310 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I311 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5825), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5438), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5814));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I312 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6020), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5936), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5825));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5815), .A(a_man[9]), .B(a_man[2]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I314 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5404), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5815), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I315 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5886), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5695), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I316 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5481), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6159), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5505), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6001), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5695));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I317 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6079), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5970), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6159));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6009), .A(a_man[9]), .B(a_man[2]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I319 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5891), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5705), .A(a_man[3]), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I320 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6152), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5961), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6009), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5705), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I321 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5770), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I322 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5858), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5672), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5886), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5585), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5404));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I323 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5481), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5672));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I325 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5682), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I326 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5411), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6088), .A(a_man[4]), .B(a_man[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I327 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6047), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5851), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5891), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6088));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I328 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5664), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5473), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I329 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6239), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6056), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5770), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5473), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6152));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I330 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5858), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5851), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6056));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I331 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5781), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5592), .A(a_man[5]), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I332 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5932), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5592));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I333 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5549), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I334 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5744), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6231), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5664), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6047));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I335 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6239), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5740), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5555));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I336 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5410), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I338 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5410));
NOR2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5682), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5704), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5492), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6191), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5704));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I344 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5593), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6251), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6087), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5593));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5492), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6251));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5674), .A(a_man[14]), .B(a_man[7]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I349 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6093), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5900), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5674));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I350 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6199), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6014), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5484), .A(a_man[14]), .B(a_man[7]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I352 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6160), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5972), .A(a_man[6]), .B(a_man[13]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I353 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5556), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6241), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I354 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5711), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5484), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6160), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6241));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I355 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6023), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5826), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5900), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6199), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5711));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6025), .A(a_man[16]), .B(a_man[9]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I357 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5610), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5425), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I358 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6100), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5909), .A(a_man[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I359 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5488), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6025), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5425), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5909));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5941), .A(a_man[15]), .B(a_man[8]));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I361 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5829), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I362 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5980), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5788), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5941), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5829));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I363 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5746), .A(a_man[15]), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I364 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5600), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5417), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5746), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5556), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5642));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I365 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5523), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5788), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5600));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I366 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6023), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6169), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6207));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5795), .A(a_man[17]), .B(a_man[10]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I368 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43523), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5795), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6066), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5687));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6209), .A(a_man[16]), .B(a_man[9]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I370 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43495), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5678), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5610), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6209), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6100));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I371 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5907), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5718), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5678), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5980), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5488));
ADDFHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I372 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6061), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5718));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I374 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43527), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43495), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43470), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43523));
ADDFHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I375 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5907), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5946), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6098));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452));
ADDFHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I378 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43527), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43492), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43474));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I379 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I381 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830));
NOR2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I383 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5445), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6126), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I384 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6130), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5549), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5932));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I385 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5820), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5632), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5781), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5972));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I386 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5640), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5445), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5820));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I387 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5517), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5451));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I388 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5417), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5826));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I389 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I390 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I392 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5744), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5632), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5939));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I395 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6161), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673));
NOR2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5483), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5971), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5483));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5807), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I404 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5807));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I405 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I406 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I407 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6232), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6232));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I417 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I419 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5789), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5789));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I423 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I424 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I425 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I426 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6214), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I427 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6214));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I432 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5764), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5764));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I436 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I438 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I439 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6195), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I442 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6195));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I443 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I444 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I445 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I446 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I447 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I448 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5747), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5526), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5747));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5776), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5526));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5607), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5776));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6035), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5607));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6222), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6035));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I456 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053));
OA21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5821), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5633));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I460 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5978));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I464 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5442), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6124), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I466 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635), .S0(a_exp[0]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I467 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248), .A(a_exp[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103));
BUFX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I471 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I472 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I473 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I474 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6027), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5910));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6027));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6045), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6044), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6045));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I479 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I480 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I481 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5841), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I483 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I484 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I485 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I486 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6099), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I489 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5653), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6099));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I490 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5841), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5653));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5849), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5796), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I495 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5796));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5694), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5469), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5694));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I498 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5469), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6150), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I500 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631), .S0(a_exp[0]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I501 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I502 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I503 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I504 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5738), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5545), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I505 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5987), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I506 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
CLKMX2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[1]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I510 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I511 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315));
NAND3BX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I512 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43412), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43412));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7197), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I516 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5831), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5831), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5521), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I521 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5501), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5521));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I523 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6181), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5805), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6052));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5805), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5618), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627), .S0(a_exp[0]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6219), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I533 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5766), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6219));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5766), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5582), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5870), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6076), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5870));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I540 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5884), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I541 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5884), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I542 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I543 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7160), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7160));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N752));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I550 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44063), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5916), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6110), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5916), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7361), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44063), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7341), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N751), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7361));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N751));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I576 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5777), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I578 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7306), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7230), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7306));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N750));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I586 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7330), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N755));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I594 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I595 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I596 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7162), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I599 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7273), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I600 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N754), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7273));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N754));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I604 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I605 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7217), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7307), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22759), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7217));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N753));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I619 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I621 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I622 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8162), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8162));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I645 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I656 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I665 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I666 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8438), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I673 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8707), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8707));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I684 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I685 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I686 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I687 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8288), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I701 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I702 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I704 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574));
OR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7904), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7809), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7904));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7956), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8438), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8288), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7809));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[29]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I723 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I724 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8417), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657));
OR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I740 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I749 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8463), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8463));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8173), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7941));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8417), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8173));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843), .A(1'B0), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8723), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8723));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I764 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8484), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I765 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I766 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I767 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I768 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I769 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I770 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I774 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8444), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8238), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8484), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8098));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[27]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7867), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8444), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I777 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043), .A(1'B1), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[27]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I778 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I779 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14655), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I782 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5461), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I786 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I787 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6142), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I788 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5461), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6142));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I789 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6139), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5948), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I790 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6119), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I791 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6119), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621), .S0(a_exp[0]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I793 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I794 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I795 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I796 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6116), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I798 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6116));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I799 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I800 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5532), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6216), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I801 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I802 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5838), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5756));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5648), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I805 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5838), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5648), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I806 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I807 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I808 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I809 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7269), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I810 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7339), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I811 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7339));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I812 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N746));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5784), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I818 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5784));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5827), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5827));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6248), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I823 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I824 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5757), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I825 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5952), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5479), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5757));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6248), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I827 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I828 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7212), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I832 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7283), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I833 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7283));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I834 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N745));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I835 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12783), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I836 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I837 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7324), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I838 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7324));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I839 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7140), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I840 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7140));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I841 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N747));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I842 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12783), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I844 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11832), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I845 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I846 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I847 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I848 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8459), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8390), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8634));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7881), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8685), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I857 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7827), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7881), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8685));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I858 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8459), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7827));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I860 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7997), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I861 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I862 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7997), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I865 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I867 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I869 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8757));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I870 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7954), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7741));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8191), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7954));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12730), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I876 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I877 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5482), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I878 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5869), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5482));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I879 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I880 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5869), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5680), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I881 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I882 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7156), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I884 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7156), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I885 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7229));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I887 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N744));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I888 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I889 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I890 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I891 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5983), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I893 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I894 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I895 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7355), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7173), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7173));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N743));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[10]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I900 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I901 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22721), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I902 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22721));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I903 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I904 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12814), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I905 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I906 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11862), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I907 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11862), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I911 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I912 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I913 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I914 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I915 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I916 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I919 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I920 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I921 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8492), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I922 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8492));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I923 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8341));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I924 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7969), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7712), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7969));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I931 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I932 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I933 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I934 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I935 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I936 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8710), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8609));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I937 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N780), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8752), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8225), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8710));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I938 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N780));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I939 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I940 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I941 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11813), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I942 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44056), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I943 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I946 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I947 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7299), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44056), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I948 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7299), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7371));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22642));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I954 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I955 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44043), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5539), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I960 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5539));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I963 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288), .A(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I965 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7354), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I966 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I967 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I968 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I969 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I970 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7316), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I971 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7316));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I972 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N741));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I973 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12844), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12844), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I976 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I978 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11623), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12730), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11813), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11562));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I979 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7125), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7125));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I981 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N748), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7195));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N748));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I984 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I985 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7252));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N749));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I990 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11796), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I992 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11796), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I993 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I994 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897));
NAND2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7923), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I997 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7834), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7923), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I999 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1002 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7721), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8061), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1004 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1005 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1006 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8257), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1007 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8257));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1008 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8517));
CLKAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1009 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7834), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8690));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1010 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1012 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1013 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12199), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1016 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1017 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11953), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11559), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12199), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11389));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1018 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12684), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12330), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11623), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12345), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11559));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11897), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12237), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1025 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6069), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1026 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6069));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1027 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1028 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1029 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7189), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1032 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7146), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7189), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1033 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7146), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1034 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7261));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1035 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N740));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1036 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43255), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1038 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43245), .A(a_exp[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43255));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1039 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1040 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1041 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1043 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43287), .AN(a_exp[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43261));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1044 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43245), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43287));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1046 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43289), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1047 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43268), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43236), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43289), .B0(a_exp[0]));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1048 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43266), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
AOI211XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1049 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43251), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288), .C0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43266));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43271), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43268), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43251));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43233), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7134), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1053 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7347), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7134), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1054 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7347), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1055 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7206));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1056 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N739));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1057 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[6]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1058 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12875), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1061 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1062 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1063 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11428), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1064 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11312), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12661), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12237), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11428));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1065 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1066 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1067 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1068 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1069 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1070 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7791), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8116));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1073 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1074 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1075 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1076 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1077 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1078 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1079 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171));
NAND2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952));
NAND4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1083 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8759));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1084 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1085 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1086 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8046), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1090 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1091 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1093 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1094 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1095 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8419), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8313), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8563));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8131), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8046), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8419));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1097 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8618), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8131));
NAND3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N776), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7791), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8525), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7747));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1099 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N776));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1100 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1102 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11398), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11968), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11246));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1105 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8549), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8449));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1109 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7964), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1113 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8297), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7964));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8783), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8549), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8297));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1115 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1116 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1117 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1119 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7928), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8783), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7928));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1124 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1125 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12381), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1126 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1127 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12763), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1128 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1129 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11852), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1131 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11214), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11852), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11625));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1132 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12087), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11575), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12381), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11214));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1133 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1134 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1136 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1137 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8457), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1138 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8472), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8457));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1139 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8472));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1140 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1142 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7669), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7669), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7733));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8571), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7936));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1148 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1149 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1150 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7986), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1151 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1152 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8605), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8705), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8605), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8705));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8182), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7986), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7688));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1157 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8182));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1158 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1159 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1161 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1165 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1166 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12273), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1168 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5911), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1169 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5911), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1171 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7333), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7333), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7290), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7151));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N738));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44049), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1180 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1183 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44049), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1184 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1185 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1186 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5635), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5447), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7243), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7276), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7352));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22635));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1196 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11186), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1197 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11186), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1198 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1200 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1201 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12840), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12273), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11467));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1202 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12715), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12363), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11195), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12012), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12840));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1203 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12805), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12453), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12715), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12661), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11683));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1204 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12174), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11785), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12742), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12087), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12805));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1205 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[38]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[37]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11398), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12174));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1206 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1207 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1208 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1210 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1211 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8511), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1212 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1213 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8653), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1215 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8671), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8455), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8671));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1217 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1218 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8120), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8653), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8455), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1219 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7730), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8138));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8029), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1224 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[19]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8511), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7730), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8029));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1225 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0]));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1226 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1227 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9909), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1232 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1233 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9945), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10070));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1234 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1235 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1236 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9930), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1237 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1238 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10349), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1239 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1240 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1241 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10159), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10349), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9992), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10308));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1242 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9960), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10159));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1243 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10086), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1248 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10278), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1249 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10234), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10489), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10278));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10416), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1251 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10416), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10025));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1252 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10334), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10384), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1255 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1256 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10046), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9908), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10334), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10384), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10432));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1257 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10147), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1260 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9937), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1261 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9914), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1262 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10484), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10066), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9937), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9914));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1263 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10318), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10180), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10208), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10484));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1264 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10103), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10046), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10318));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1265 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1266 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10528), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1269 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1270 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10286), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1271 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10014), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10512), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10528), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10413), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10286));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10478), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1276 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10281), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10509), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10263), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10478));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1277 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10125), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10014), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10012), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10281));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1278 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9908), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10180));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1279 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1280 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10133), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1281 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10140), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1282 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10356), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1283 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10170), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10038), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10133), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10140), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10356));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10362), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1287 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10505), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1289 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10059), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9922), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10149), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10505));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1290 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10442), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10198), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9995), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10059));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1291 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9932), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10418), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10512), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10170), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10442));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1292 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9932), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10338), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9991));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1296 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1297 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10498), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1298 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1299 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10328), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10224), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10498), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9929));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1300 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10094), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10328), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10307));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1301 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10150), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10094));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1302 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10511), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10214), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1305 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10526), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1306 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9946), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10431), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10511), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10214), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10526));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10342), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1308 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9980), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10471), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10342), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9922));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1310 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10078), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1311 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10091), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1312 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10218), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10085), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10276), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10078), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10091));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10423), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1314 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9942), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1315 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1316 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10456), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9942), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10011));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10237), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1319 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10182), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10050), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10226), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10237));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1320 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10500), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10348), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10456), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10182), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10431));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1321 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10245), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10113), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10218), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10191), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10500));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1322 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9980), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10245), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9959));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1323 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1325 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1326 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1327 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1328 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5785), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1329 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5785));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1330 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5935), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7121), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1335 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7220), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1336 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7293), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7178), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N736), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7293));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1338 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N736));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1344 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10419), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10284), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10294), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9958), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9970));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1345 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10104), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9955), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9982), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10419));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10306), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10319), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1349 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1350 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6049), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6049), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7319), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1354 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7165), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7319), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1355 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7165), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43414), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7123), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1357 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43404), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43414));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1358 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43404));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1359 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[2]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1361 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10386), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10247), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10319), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9975));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1362 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1363 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6242), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1364 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1365 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7364), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7364), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7182), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7321), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7182));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N734));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1372 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[1]));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22602), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10305), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22602));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1376 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10310), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10305), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10062));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1377 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10339), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10353), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10310));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1378 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10024), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1379 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1381 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10040), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10538), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10024), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10154), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10090));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10439), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10421), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1384 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1385 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10075), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10439), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10421), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10329));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1386 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9993), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10488), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10284), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10040), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9935));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1387 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10029), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9971), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10339), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9993));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1388 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10371), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10075), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10050), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10321));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1389 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10136), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10085), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10371));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1390 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10348), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10002));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1391 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10471), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10113));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1392 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1395 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10049), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10324), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1398 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10004), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10049), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10518), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10324));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10409), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1404 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1405 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1406 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1407 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6075), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5475), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5848), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5848));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5475), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7163), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N608), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7163), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7309), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7209), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7127), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7267), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1417 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7127));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N733));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1419 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10168), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1422 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10271), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10409), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10368), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10168));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1423 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9961), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10445), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10004), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10087), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10271));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1424 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10228), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10096), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10172), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10538), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10247));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1425 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10260), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10206), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10228));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1426 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10260), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10238), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10527));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1427 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
ADDHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1431 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10052), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9912), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10054), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10396));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1432 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10223), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10126), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1435 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10322), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10126), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10230));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1436 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9923), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10410), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9948), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10052), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10322));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1438 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10382), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1439 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10137), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1440 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9973), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10460), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10102), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10382), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10137));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1442 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1443 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10483), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1444 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10288), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10155), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9953), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10483));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1445 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10239), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9912));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1446 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10192), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10063), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10503), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9973), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10239));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1447 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10516), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10361), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9923), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10192), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10445));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1448 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10516), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10488), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10128));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10031), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1456 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10109), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9939), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10111), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10031));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10015), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10118), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1460 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10466), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10326), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10015), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10118));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10211), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10380), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1464 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9951), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10436), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10211), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10380), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10280));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1465 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10507), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10351), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10109), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10466), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10436));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1466 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9934), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1467 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10301), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9934));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9947), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10205), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1471 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10414), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10494), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10205));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1472 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10335), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9947), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10275));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1473 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1474 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10041), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9933), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1476 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10068), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9928), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10036), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10041), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9933));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10388), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1479 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10221), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10089), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10388), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10164));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1480 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9986), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9928), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9951), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10221));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1481 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10196), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10477));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10130), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472));
ADDHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1483 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9903), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1484 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10097), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9965), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10389), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10414), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10068));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1485 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1486 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1489 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10173), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10042), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10470), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10203));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1490 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10311), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1493 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10447), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10312), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10311), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10219), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10487));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1494 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10363), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10335), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10042), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10312));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1495 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9986), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9965), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10231));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1496 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10491), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10447), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10155), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10173));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9964), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1498 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10401), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10502), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1500 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9938), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10422), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9964), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10401), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10502));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1501 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10127), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1502 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10112), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1503 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10209), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10077), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10127), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10112), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9903));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1504 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10129), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10422), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10077), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10097));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1505 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10363), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10341), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9994));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1506 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10017), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1510 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9997), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10496), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10017), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10290));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1511 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10476), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1512 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10359), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1514 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10265), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10476), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10359), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10373));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1515 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10376), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10242), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9997), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10265));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1516 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10376), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10089), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10351));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9927), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1520 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10523), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9920), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1521 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10021), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10189), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1523 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10425), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10021), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10189));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10443), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1528 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10232), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10100), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10443));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1529 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10081), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10195), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10232));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1530 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10292), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9941));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10469), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1532 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9916), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10425), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10469), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10496));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1533 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10132), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10081), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10402));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10035), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056));
NOR2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10171), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1537 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10316), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10177), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10267));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10535), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1540 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1541 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10393), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10448));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1542 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9967), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10098), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10393), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10177));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1543 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10100), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10316), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9967));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10379), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9999), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10347), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
ADDHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1550 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10122), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10246), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10347));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1551 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10122));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10468), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1556 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10084));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10266), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10354), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10134), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10480), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10266), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10354), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10134));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10404), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10314), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9919), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10480), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10404));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10079), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10188), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10314), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10058));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10327), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10464), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10468), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10079), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10327));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10142), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10110), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10464), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9978));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10446), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10379), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10142), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10244));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10051), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10035), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10446), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10534));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1576 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9976), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9916), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10242));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10303), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1578 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009));
CLKAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10255), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10303), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10166), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10438), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9972), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10166), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10438));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9972));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10385), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10051), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10255), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10123));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10385));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1586 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10440), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9957), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10169), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10440));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10092), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10357));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1592 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10529), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10374), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10185), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9938), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10209));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1593 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10162), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10460), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10106), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10491));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1594 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10129), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10374), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10032));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1595 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1596 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10473), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10410), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10138), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10529));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1597 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10063), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10331));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1599 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1600 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10473), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10361));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1604 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1605 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1619 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1621 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1622 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9988), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9988));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10289), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10479), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10289));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10387), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10479));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10076), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10387));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10372), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10207), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10076));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10146), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[32]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10372), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10146));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10243));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9996), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1645 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10463), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9996), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10241), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10463));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10117), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1656 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10420), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10117));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9936), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10420));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10241), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1659 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12770), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12051), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[32]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12770));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12051));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11613), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1665 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1666 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12416), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8591), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8144));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1673 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7993), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8247), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431));
NAND3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8322), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8573), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8107), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8322), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8573), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1684 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8247), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8107));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1685 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7972), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8591), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8287));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1686 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1687 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7854), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7877), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8054), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8344), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7854), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7877), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8054), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7972), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8344));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1694 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11894), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11506), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11613), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12416), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12556));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8348), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8038), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8348), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1701 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7761), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1702 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7829), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1704 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8385), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8303), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8385));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8659), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7829), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8303));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7781), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8659));
CLKAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8038), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7781));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12190), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12044), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1717 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12751), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12401), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12044), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11233));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12799), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11891), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1723 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11254), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12607), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12799), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11891), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11686));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1724 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12634), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12751), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11254), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12489));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1725 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11752), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12571), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11894), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12634));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12446), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11501), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11647), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1732 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12156), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11762), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12446), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11501), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11647));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11961), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12309), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11218), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1740 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8560), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8560));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7678), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7860), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7678), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7940));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1749 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7903), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8436), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7903), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8325));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754));
NOR3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7805), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8479));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8676), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8436), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7805));
NAND3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7701), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7860), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8676));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N771));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11803), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1764 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11379), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12722), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11803));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1765 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11792), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11407), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12156), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11379), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12607));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1766 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11657), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11792), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11506), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12280));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1767 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12516), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12149), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12363), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11370));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1768 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11858), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12453), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11752), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12516));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1769 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[37]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[36]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11785), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11858));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1770 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[37]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[19]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[37]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7898), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1774 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8428), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1777 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1778 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8610), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1779 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7911), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8610), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1782 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8358), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8358));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8319), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8753));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1786 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8319));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1787 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[18]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7898), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8428), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7911), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7691));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1788 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1789 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1790 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1791 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8788), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8367));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8652), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8788), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1793 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1794 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8512), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1795 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1796 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22714), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8512), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8652), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22714));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1798 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12260), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1799 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8141), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1800 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1801 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1802 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7950), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1805 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8053), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7950));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1806 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8053));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1807 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22705), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8141), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7910));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1808 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1809 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8608));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1810 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11492), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1811 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1812 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10493), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10465), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10493));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10325), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10465), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1818 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10055), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9915), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11925), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1823 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11532), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12866), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11492), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12149), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1824 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[36]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[35]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12260), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11532));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1825 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[36]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[18]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[36]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1827 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1828 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12834), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11926), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1832 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11729), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11351), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12834), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11926), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11755));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1833 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1834 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1835 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1836 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1837 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8152), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1838 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8039), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1839 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8401), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8039));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1840 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1841 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1842 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7764), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1844 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7764));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1845 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8020), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1846 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8020), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1847 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8351), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8740), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7994));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1848 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8778), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267));
NAND4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N770), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8152), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8401), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8351), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8778));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N770));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11418), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12083), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1857 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11512), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11418), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12083), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12229));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1858 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11160), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12526), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11729), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12589), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11512));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1860 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11995), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1861 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1862 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1865 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11844), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1867 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12100), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11702), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12341), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11844));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1869 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1870 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12484), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1876 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12821), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12466), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11536), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11680));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1877 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12284), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11901), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12100), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11269), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12821));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1878 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11932), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11762), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12722), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12284));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1879 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12547), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11160), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12401), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11932));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1880 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1881 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1882 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1884 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8355), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7975));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1885 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8650), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1887 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1888 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8276), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8565), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7683));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1889 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1890 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1891 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7946), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8276), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8178));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1893 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1894 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1895 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7843), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8422), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7843));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1900 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8082), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7918));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1901 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8558), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8082));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1902 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8762), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8422), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8558));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1903 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8527), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8762));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1904 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1905 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1906 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1907 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12871), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11826), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1911 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12650), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12871), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11963), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11826));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1912 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11870), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11484), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12620), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12756), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12650));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1913 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11289), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11351), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12849), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11870));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1914 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12668), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12314), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11289), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12526), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11542));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1915 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11568), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11407), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12184));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1916 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12427), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11280), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12547), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11568));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12869), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12869));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1919 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243));
XNOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1920 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1921 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1922 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1923 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1924 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7974), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8556), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7974), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8684), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8460), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1931 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8594), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1932 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8165), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8460), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8594));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1933 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8684), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8165));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1934 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8556), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22699));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1935 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12471), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1936 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11441), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12777), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12626), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12471), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12059));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1937 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[35]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[34]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12866), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12427), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11441));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1938 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1939 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8775), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1940 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8204), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8540), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8775));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1941 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1942 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1943 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7717), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1946 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8072), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1947 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8204), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7717), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8072));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1948 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[35]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[17]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[35]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8300), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1954 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8300));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1955 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7998), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8522), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1960 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7776), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7776));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1963 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7857), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7743), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8477), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8328), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7998), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7857));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1965 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8328));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1966 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1967 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8092), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1968 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1969 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7858), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1970 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1971 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8092), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7858), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8579));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1972 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[16]));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1973 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11708), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1976 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10403), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10403));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1978 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10131), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1979 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1981 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10264), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10175));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10285), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1984 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10152), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1985 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10285), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10152));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10264), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10381), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293));
XNOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10381), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105));
AO21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1990 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12339), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11708), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11185));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1992 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11460), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1993 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1994 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12262), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I1997 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12440), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11460), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12119), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12262));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I1999 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8490), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8729), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2002 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8242), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2004 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2005 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7798), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2006 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7968), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7798));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2007 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2008 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7871), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2009 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7709), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7871));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2010 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8069), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8490), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8729), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7968), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7709));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2012 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2013 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8299), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8069), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8299));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2016 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12408), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2017 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2018 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[1]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22556));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2025 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2026 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12474), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2027 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11459), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12791), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11304), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12474));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2028 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12613), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11702), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12440), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11459));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2029 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12065), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11664), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11901), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12613), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12642));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7815), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8677), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2032 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7976), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7815), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8677));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2033 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2034 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7976), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2035 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2036 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2038 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7762), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2039 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8042), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7762));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2040 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7887), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8042));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2041 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7887));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8212), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44103));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2043 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12677), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2044 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11692), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11319), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12314), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12065), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12677));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2046 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2047 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11342), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12269), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11959));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2048 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[34]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[33]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12339), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11342));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2049 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[34]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[16]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[34]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2053 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12279), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2054 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12279));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2055 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2056 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2057 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2058 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11685), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12792), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2061 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2062 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2063 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12334), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2064 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2065 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12001), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2066 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12299), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12334), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12001));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2067 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2068 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2069 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11268), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12792), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12299), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12658));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2070 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12518), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2073 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11570), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2074 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2075 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11720), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2076 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12265), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11880), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12518), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11570), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11720));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2077 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12228), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11843), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11268), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12265), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12075));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2078 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11640), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11484), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12466), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12228));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2079 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10343), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10199), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2083 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10495), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10199));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2084 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10343), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10495), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2085 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2086 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10080), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9940), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450));
MX2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10080), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9940), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11715), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2090 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11715), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2091 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12785), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11640), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2093 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11888), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2094 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12460), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12094), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11685), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12785), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11888));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2095 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8260), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2097 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8078), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8260), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8078));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2099 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8308));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2100 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8001), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8132));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2102 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2105 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8372), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8697), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8235), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8667), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8372));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8235));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11945), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2109 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7862), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8607), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7862), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8708), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8607));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2113 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7896), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2115 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8123), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2116 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8439), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7896), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8123));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2117 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7851), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8439));
CLKAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8708), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7851));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2119 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12035), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12107), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2124 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2125 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2126 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11306), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12657), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11188), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12151), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11920));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2127 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12043), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12035), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12107), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11306));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2128 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11235), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12791), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12291), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12043));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2129 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12407), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12034), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11235), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12256), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11261));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11310), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2132 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11833), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12407), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11310));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2133 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2134 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11499), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2136 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8681), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2137 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2138 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8641));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2139 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2140 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7797), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7708), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7797), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2142 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8782), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7708), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8601));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44095), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8782), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8102));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2148 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8681), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44095));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2149 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11172), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2150 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2151 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11493), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2152 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8576), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7789), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8386), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7789));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2157 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2158 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8249), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8630));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2159 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7878), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8576), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8249));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2161 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8147), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8229), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8538), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8056), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8309), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2165 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8772), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8056), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8309));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2166 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8538), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8772));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8495), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8370));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2168 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7878), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8495));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2169 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11638), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2171 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12300), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2173 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12082), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11493), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11638), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12300));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2174 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12765), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12415), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11880), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12082), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12619));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2175 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12011), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11843), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12765), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12588));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095));
XOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12830), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2180 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12830));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12491), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2183 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11417), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12758), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11172), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12011), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12491));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2184 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12581), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12221), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11499), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12435), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11417));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2185 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11476), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12813), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11319), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11833), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12581));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2186 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[33]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[32]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12460), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11476));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7763), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8112), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7763));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8258), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2196 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8293), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8010));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2197 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8293));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2198 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8599), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7971));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2200 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8151), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8234));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2201 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[15]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8112), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8545), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8599), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8151));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2202 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[33]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[15]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[33]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2203 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2204 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2205 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2206 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7726), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2207 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8784), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2208 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8468), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8784));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7682), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8468), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2210 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8420), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7726), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7682));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2211 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7793), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8420));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2212 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8507), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2213 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7945), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[14]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7793), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8507), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7945));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2215 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10000), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450));
XNOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10000), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2217 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2218 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10291), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2219 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10156), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43775), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43757), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43743), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43775));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2224 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10291), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10156), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2225 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2226 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11620));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2227 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12552), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11606), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2232 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2233 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12837), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12483), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12552), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11606), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11757));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2234 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2235 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2236 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2237 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12825), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2238 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2239 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12072), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2240 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11890), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11500), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12825), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12072));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2241 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11854), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11466), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12837), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11890), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12657));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2242 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2243 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12441), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11339), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2248 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2249 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7938), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8209));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2251 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7938));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2252 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8754), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7978));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8559), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2255 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8559), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2256 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7784), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8169));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2257 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8520), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7784), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831));
CLKAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8754), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8520));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2260 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2261 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11262), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2262 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12118), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11721), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11919), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11956), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11262));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2263 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12798), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12441), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11339), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12118));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2264 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11812), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11427), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11854), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12798), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11649));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2265 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12729), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12383), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11812), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11612));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2266 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2269 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12192), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12729), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12034), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12660));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2270 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2271 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8655), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2274 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7894), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8062));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2276 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8160), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2277 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2278 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2279 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2280 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8706), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7732), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2281 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7894), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8160), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8706));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2282 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8655), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44087));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2283 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12168), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2284 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11672), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2286 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2287 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12186), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7863), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2289 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2290 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7811), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7863), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8022));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2291 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8541), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7811));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8394), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8541), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8636), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8394), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8636));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2295 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2296 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2297 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12150), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11672), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12186), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12614));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2298 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2299 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11228), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2300 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2301 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12549), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2302 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12367), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12549));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2303 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2304 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12333), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2305 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2306 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11529), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2309 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12870), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12519), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12333), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11529), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11371));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2310 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12627), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12274), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12150), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12367), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12870));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2311 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12596), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11679), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12448));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2312 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12561), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12415), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12596), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11427));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2314 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12122), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2315 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11772), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11388), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12168), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12561), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12122));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2316 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12831), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2318 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11194), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11772), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12831), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12758));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2319 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11602), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11449), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12192), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11194));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2320 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[32]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11602), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12094), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12813));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2321 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[32]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[32]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2322 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2323 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2324 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12481), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2325 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2326 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12306), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2327 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12530), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12162), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12306), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12481), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12383));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2328 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12593), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2329 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12593), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2330 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43395), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43395));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2335 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2336 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11541), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2337 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2338 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11924), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2339 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12351), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11977), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12202), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11924));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2344 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8537), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8143), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8771), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8537));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8055), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2348 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8323), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2349 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2350 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8430), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8003), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8430), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8003));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8246));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2354 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7703));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2355 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8055), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8323), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8012));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8143), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44079));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2357 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11393), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2358 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11654), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12483), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11721), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11500));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2359 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11621), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11466), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11654), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12236));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2360 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2361 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11723), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2362 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11584), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11393), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11621), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11723));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2363 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11549), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11168), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12351), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11584), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11388));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2364 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11967), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12530), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11802), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11549));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2365 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[31]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[30]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12221), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11224));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8280), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8379), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8340), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8280), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8379), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2369 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8624), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8770), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8624));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8340), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8770));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2372 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8086), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8086), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8006));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7965), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8103));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8196), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7965));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2378 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[31]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[13]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[31]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2379 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2381 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2382 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2384 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8356), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2385 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8356));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2386 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8071), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2387 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8466), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2388 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8027), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8466));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2389 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8469), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8071), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8027), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2390 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8469));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8218), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8701));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2392 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788), .A(1'B1), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[26]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8088), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2395 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8362), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7799), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8088), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8362), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7873), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2401 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7735), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2402 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8243), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8426), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7735));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2403 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[25]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7799), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7873), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8243));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2404 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541), .A(1'B1), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[25]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2405 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2406 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2407 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2408 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[42]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8647), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8036), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8647), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7890), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7672), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7890));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8302), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2417 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8410), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7672), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8302));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7779), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8658), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8410));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2419 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8036), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7779));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2420 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[24]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[41]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[42]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2423 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7786), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2424 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8326), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7786));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2425 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2426 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2427 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8127), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8474), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8127), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8474));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2432 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2433 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7855), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7698), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7855), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2436 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8190), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7953), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7698));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[23]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8326), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8190));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2438 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2439 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11730), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2442 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[41]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[40]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11730));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2443 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[41]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[23]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[41]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2444 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2445 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2446 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2447 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2448 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7886), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8396));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8255), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8597), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8255));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8210), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8597));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2453 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7919), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[22]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7886), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8210), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7919));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2456 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11886), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2460 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12695), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2462 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12479), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11771), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12695));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2463 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[40]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[39]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11352), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11886), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12479));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2464 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[40]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[22]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[40]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2466 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8101), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2467 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7839), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2468 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7839));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7819), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8175));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2470 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8664), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2471 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8523), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8664), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2472 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8101), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7819), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8523));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2473 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[39]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[38]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12116), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11953), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12684));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2474 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[39]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[21]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[39]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2475 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2478 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2479 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2480 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2481 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2483 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8295), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8065), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8447));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2484 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8779), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7750), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8622), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8295));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2485 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8779));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2486 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[38]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[20]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[38]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2489 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2490 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12115), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2495 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43770), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43770));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43769), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2498 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2499 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43769), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2500 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43747), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2501 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229));
MX2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2502 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43755), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43747), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2503 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11523), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2504 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2505 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2506 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2510 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12403), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12029), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12582), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11957), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12609));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2511 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2512 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12475), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2513 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11793), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2516 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8310), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8561), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8418), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8310), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8561));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8580), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2521 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7838), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8580));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2522 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7942), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7838));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2523 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8418), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7942));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2524 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2525 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8504), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2526 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8075), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8504), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8174), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8075), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8213));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7790), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8174));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8045), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7790));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12254), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2533 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12185), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11795), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11793), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11298), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12254));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2534 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11927), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12403), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12475), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12185));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12717), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12862), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2540 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2541 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11187), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12551), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12717), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12862), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12108));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2542 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12663), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11756), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11187), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12519));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2543 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12423), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12053), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12663), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12274));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2546 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2547 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11710), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2548 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2549 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12648), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2550 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11453), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12788), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11710), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12648), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11563));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2554 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12224), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2555 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12437), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12068), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12224));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7748), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2559 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7748), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8485));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8446), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8099), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8336));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2563 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8620), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2564 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8004), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2565 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8620), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8004));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8134), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7706), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8134));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8585), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7706));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7817), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8446), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8679));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7868), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8064), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7868));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7817), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8064));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2575 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11871), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2576 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2577 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12508), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2578 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12223), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11836), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12368), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11871), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12508));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2579 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11962), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11569), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11453), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12437), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12223));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2580 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11687), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11314), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11962), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11994), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11535));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2581 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11434), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12775), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11275), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12053));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2582 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12388), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12018), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12423), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11434));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7883), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2584 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8167), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7883));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2585 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8461), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2586 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7782), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8461), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8206));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2590 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8167), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7782), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8275));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12386), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11344), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2594 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11395), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12736), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12386), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11239), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11344));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2595 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11360), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12388), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11395));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2596 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2599 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2600 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11718), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2602 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12170), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11161), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11531), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11718));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2603 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12136), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11740), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11201), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11977));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2604 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12318), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11939), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11360), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12136));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2605 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[30]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[29]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12555), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11577));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7693));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8033), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7935), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2610 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8345), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7824), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8161), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8345), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7824), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2615 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8656), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8161));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2616 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8033), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8656));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2617 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[30]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[12]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[30]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2619 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12692), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12340), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12029), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11795), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12551));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2621 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11993), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2622 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12669), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2624 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11704), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11328), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11993), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12669));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11411), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11180), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2630 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8470), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2631 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8265), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8028));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8703));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8546), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7983), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8219));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8084), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8546));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7684), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8158));
AND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8568), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7684));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2645 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2647 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12257), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11873), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11180), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11485), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12752));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2648 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11227), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12584), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11411), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12257));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11837), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11333), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2655 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11488), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12822), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11837), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11333), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12292));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2656 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12004), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11605), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11488), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12068), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12788));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2657 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11725), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11346), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11227), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12004), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11569));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2658 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12455), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12089), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12308), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12692), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11725));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7982));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8232), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7788), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2665 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8581), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2666 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8315), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8581));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8232), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7788), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8315));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8416), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8437), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8058), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8416));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11619), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2673 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12209), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11821), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12455), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11619), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12690));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12505), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12505), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22]));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514));
CLKINVX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22582));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12344), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2684 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2685 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11207), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12775), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12344), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12525));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2686 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11174), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12209), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12018), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11207));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2687 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10235), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10235), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10099), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12350), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12350));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2695 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11472), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12807), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11314), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12089));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12868), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11337), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2701 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11987), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11472), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12868), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11337));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2702 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11948), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12736), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11780));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2703 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12857), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12502), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12703), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11174), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11948));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2704 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[29]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[28]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12857), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11168), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11939));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8324), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8673), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7738), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8324), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8189), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8365));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7695), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[11]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8673), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8189), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7695));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2714 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[29]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[11]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[29]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12155), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11969), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2723 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12515), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2724 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11249), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12155), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11969), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12515));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7723), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8642));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8602), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8503));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8019), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8113), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8019));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7723), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8602), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8113));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[8]));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12592), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11595), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11748), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12723), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2740 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12705), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11748), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12723));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12143), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11451), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8342), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7960));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2749 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8342));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8454), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7744));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8427), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8052), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8427), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8052), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7801), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7801), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8732), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7874));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8590), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7711));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8454), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8198));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12819), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2764 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11525), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11451), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12402), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12819));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2765 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11264), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12616), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12143), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11525));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2766 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12725), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12375), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11264), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11836), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12584));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2767 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12493), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12340), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11346));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2768 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2769 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2770 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12245), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12592), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12493), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12338));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2771 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12710), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11249), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12245), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11821));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2774 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11979), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11979));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2777 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2778 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2779 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11387), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2782 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11910), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2786 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12506), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12679), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11910), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12542));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2787 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12038), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12822), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12506), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11873));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2788 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2789 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11521), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2790 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2791 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11362), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2793 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12323), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2794 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11782), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11521), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11362), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12323));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2795 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2796 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12030), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2798 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12740), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12389), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11329), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12030));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2799 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2800 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11217), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2801 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2802 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12789), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12179), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2805 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12538), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11217), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12789), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12179));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2806 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12293), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11913), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11782), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12740), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12538));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2807 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12759), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12410), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12293), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11328), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12616));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2808 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11765), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11382), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11605), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12038), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12759));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2809 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10047), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2810 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10047));
NAND2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2811 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[18]));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2812 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11301), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12653), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12859), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12138), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12352));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11786), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12319), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2818 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11823), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11436), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11786), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12319), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12711));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12467), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11949), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2823 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2824 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2825 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12573), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2827 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12568), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12211), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11634), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12573));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2828 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11558), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12467), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12568));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12858), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2832 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12438), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2833 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11552), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2834 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2835 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12066), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2836 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12604), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12247), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11552), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12066));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2837 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11591), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11211), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12858), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12438), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12604));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2838 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12327), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11396), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12389), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11591));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2839 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12076), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11558), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12327), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11913));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2840 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11805), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11421), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11642), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11301), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12076));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2841 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12527), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12158), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12375), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11805));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2842 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11508), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12842), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11765), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11387), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12527));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2844 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2845 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12024), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11508), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12686));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2846 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11747), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11363), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12024), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12566), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11589));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2847 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12678), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12326), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12710), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11747));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2848 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[28]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[27]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12678), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11740), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12502));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8226));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8557), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8498), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7673), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8557), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8498));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8686), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[10]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7673), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8686), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2857 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[28]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[10]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[28]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2858 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2860 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11576), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2861 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2862 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11763), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12148), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2865 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11283), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12637), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11763), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12148));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2867 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7728), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2869 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8133), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7728), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2870 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8421), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8589));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8262), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8421));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8237), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8262), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2876 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7844), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2877 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8133), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8237), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8550), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7844));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2878 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11850), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2879 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12281), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11896), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11960), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11850), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12124));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2880 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12745), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12395), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11283), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12281), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11859));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2881 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2882 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12731), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2884 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11566), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2885 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11544), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11163), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12731), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11382), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11566));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2887 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12329), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2888 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2889 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11193), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2890 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8552), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2891 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8731), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8068), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8731));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2893 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8381), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2894 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8452), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2895 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7930), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8381), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8452));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8787), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8552), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8068), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7930), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8787));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[6]));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2900 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12797), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2901 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2902 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11378), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2903 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12315), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11934), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11193), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12797), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11378));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2904 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12061), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11659), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11544), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12329), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12315));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2905 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11788), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11401), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12061), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12601), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11626));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2906 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12511), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12142), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12357), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12745), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11788));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2907 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[27]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[26]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12511), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11556), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12326));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7999), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8273), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2911 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7861), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8273), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7899), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2912 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8330), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7861), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2913 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2914 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[9]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2915 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[27]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[9]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[27]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2916 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2919 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2920 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11754), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2921 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2922 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2923 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10315), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258));
CLKMX2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2924 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10315), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11256), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2931 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12398), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12503), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11256), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12216));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2932 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2933 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2934 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2935 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2936 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2937 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12358), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2938 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11628), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11251), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11557), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11402), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12358));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2939 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12360), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12398), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11628), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11436));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2940 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11335), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12682), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12360), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12172), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11176));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2941 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12794), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12443), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12653), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11335));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2942 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2943 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[18]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2946 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12558), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12194), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12794), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12410), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12200));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2947 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11322), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12158), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11754), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12558));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2948 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12779), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12430), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12842), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11322), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11896));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11955), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12382), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2954 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11184), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2955 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11579), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11197), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12382), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11421), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11184));
AND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7852), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8709), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2960 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7991), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7991));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7690), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7852), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8709), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8321));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2963 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[5]));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12078), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2965 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2966 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12721), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2967 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2968 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2969 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12346), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12078), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12721), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12557));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2970 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12096), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11695), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11955), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11579), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12346));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2971 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11827), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12637), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11659));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2972 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12541), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12779), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12395), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11827));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2973 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[26]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[25]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11363), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12142));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8722), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8678), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8722));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2976 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7765), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8678));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8063), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2978 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8153), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2979 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8021), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8063), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8153), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8741), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8021));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2981 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7888), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7765), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8741));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8402), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[8]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7888), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8402), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2984 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[26]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[8]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[26]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2985 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8026), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8510), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8277), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8026), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8510));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8180), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2990 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7729), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7794), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2992 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8763), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8180), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7729), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7794));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2993 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8277), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8763));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2994 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I2995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11368), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2997 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11985), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I2999 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12611), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3002 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11445), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12782), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11666), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12611));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11775), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3004 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12253), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11868), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11775));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3005 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12531), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3006 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3007 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11828), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3008 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12433), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12531), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11828));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3009 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11404), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12748), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11445), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12433), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12247));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3010 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11364), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12712), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12211), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11211), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11404));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12595), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3012 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12111), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11716), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11951), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11364), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12595));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3013 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11847), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11463), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12111), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11675), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12443));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11561), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3016 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11354), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11368), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11847), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11561));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3017 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12815), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12462), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11163), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11934));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3018 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11811), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12009), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12548), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3025 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12591), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11811), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12009), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12548));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3026 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3027 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11173), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3028 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3029 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12746), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3032 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3033 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11292), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3034 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11258), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12612), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11442), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11868), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11292));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3035 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12218), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11830), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11173), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12746), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11258));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3036 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12182), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11790), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12026), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11251), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12218));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11853), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3038 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12145), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12182), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11989), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11853));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3039 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12829), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12477), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12145), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12682), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11716));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3040 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8735), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3041 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3043 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7757), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3044 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7715), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7757));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22659), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8735), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7715));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3046 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7915), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3047 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8388), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3048 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7915), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8388));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3049 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22659), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8494));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11303), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12374), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3053 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11616), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12829), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11303), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12374));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3054 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12130), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12591), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12194), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11616));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3055 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43997), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12670), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12130), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11695));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3056 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12574), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43964), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12815), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12430), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43997));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3057 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[25]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[24]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11401), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12178));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3058 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[25]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[25]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3061 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8205), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3062 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8282), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8205));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3063 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8166), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8282));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3064 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8166));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3065 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8730), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3066 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7710), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8730), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3067 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8453), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7710));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3068 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8009), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3069 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8104), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8009));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3070 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7823), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8453), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8104), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8070), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7823));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3073 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12714), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3074 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3075 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3076 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3077 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3078 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12384), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12014), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12714), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12191), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11178));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3079 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12851), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12497), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11971), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11197), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12384));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11614), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3083 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11429), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3084 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3085 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12394), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3086 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12537), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3090 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12033), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12394), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11590), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12537));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3091 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11220), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12062), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12033), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12782));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12800), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3093 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11182), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12748), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11220), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12800));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3094 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12864), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12512), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11182), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12712), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11750));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3095 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11884), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11495), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11614), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11429), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12864));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7783), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3097 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7830), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7885), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3099 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8661), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7885));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3100 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8519), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7830), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8661), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3101 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7783), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8519), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3102 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12297), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3105 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3108 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12623), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12297), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12183), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12000));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3109 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11391), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12732), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11884), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11463), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12623));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3113 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11801), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3114 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11652), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11272), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12365), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11801), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12477));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3115 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12164), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11652), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12231), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11236));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3116 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43976), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43960), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12697), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11391), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12164));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3117 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43957), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12462), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12851), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43976));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3118 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[24]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43994), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43935), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43957), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43964));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3119 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[24]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[24]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3121 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12764), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3124 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11863), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3125 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3126 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3127 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3128 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11840), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11456), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11863), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12733), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12025));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3129 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3130 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12252), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3132 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3133 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3134 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3136 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3137 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12586), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12226), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11208), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12780), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12643));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3138 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12754), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12405), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11840), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12252), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12586));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3139 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11998), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11599), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11830), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12754), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12578));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3140 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11958), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11564), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11790), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11998), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12545));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3142 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3143 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11922), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11958), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12764), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11234));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3145 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12539), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11791), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3148 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8008), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3149 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8008));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3150 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8582));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3151 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8440), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3152 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7810), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8233), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8440), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7810));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3155 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7958), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22651));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11526), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3157 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3158 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3159 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12659), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12303), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11791), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11526), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11601));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3160 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12418), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12047), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11922), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12539), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12659));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3161 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3162 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11419), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3165 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11682), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11307), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11419), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12512));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3166 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11430), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12768), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11682), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11495), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12267));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3167 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11169), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12533), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12418), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12014), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11430));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3168 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43938), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11732), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12497), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11169));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3169 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43987), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43973), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43938), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43982), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43944));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3171 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7917), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8360), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7917));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44116), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8360), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43954), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44116));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8301), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7990), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7990));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43941), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8301), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7882));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43985), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43954), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43941));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3180 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43985), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43994));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3183 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3184 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3185 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14822), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3186 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12431), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3192 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12196), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11809), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12431), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11627), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12567));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12013), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11479), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3196 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11425), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12761), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12013), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11479));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3197 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11610), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12196), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11425), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11456));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3198 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11800), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11415), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11636), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12612), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11610));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3199 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12081), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3200 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12719), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12371), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11800), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12081), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11599));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3201 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3202 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12406), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3203 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3204 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11215), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3205 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11538), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12371), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12406), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11215));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3206 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3207 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12414), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3208 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3209 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12587), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3210 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12688), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12719), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12414), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12587));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3211 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8076), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3212 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8562), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3213 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3214 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3215 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8403), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8294));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3216 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7979), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8743), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8403), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3217 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8533), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201));
NOR4BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3218 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8562), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7979), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8533));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3219 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12507), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3220 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3221 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11408), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3222 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3223 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3224 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11722), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11340), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11408), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11225));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3225 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12276), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11892), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11538), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12336), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11340));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3226 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3227 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12045), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3228 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11305), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3229 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3230 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11904), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3231 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11237), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3232 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3233 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12060), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3234 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12535), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12167), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11904), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11237), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12060));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3235 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3236 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12286), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3237 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11199), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12559), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12286), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12761));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3238 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12379), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12008), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11199), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12226), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11231));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3239 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12554), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11305), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12405), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12379));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3240 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3241 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3242 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3243 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11758), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11376), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12554), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12230));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3244 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3245 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11784), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3246 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8702), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3247 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3248 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8724), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8702), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8183));
NAND3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3249 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8473), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3250 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8136), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3251 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8335), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8724), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8473), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8136));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3252 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8529), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3253 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8529));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3254 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8335), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7749));
OAI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3255 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11746), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3256 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3257 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3258 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3259 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12580), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3260 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12522), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12153), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11746), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12750), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12580));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3261 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11502), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12838), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11758), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11784), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12522));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3262 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3263 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12744), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3264 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3265 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12570), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3266 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3267 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11267), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3268 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3269 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12461), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3270 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3271 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11660), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3272 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3273 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12602), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3274 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12656), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12296), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12461), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11660), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12602));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3275 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3276 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11247), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3277 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3278 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12816), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3279 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12232), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3280 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3281 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11514), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3282 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11917), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11527), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12232), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11514));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3283 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11555), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11171), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11247), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12816), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11917));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3284 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12321), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12167), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12656), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11171));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3285 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11528), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3286 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11973), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11555), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11809), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12559));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3287 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12700), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12348), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12321), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11528), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11582));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3288 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3289 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3290 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12161), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11768), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12700), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11267), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11458));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3291 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12125), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11728), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12744), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12570), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12161));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3292 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3293 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11648), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3294 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12706), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3295 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11572), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11191), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11648), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11415), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12706));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3296 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3297 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11397), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3298 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12301), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3299 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11385), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12728), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11973), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12301), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12008));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3300 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3301 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11845), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3302 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12343), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11966), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12188), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11385), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11845));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3303 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12311), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11929), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11572), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11397), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12343));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3304 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12091), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12872), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11929));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3305 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12056), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11655), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11892), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12838), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12091));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3306 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12239), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11502), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11307), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12276));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3307 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3308 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11592), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3309 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3310 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3311 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12486), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11592), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12757), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11564));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3312 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11468), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12802), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11530), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12486), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12303));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3313 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3314 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3315 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12449), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12085), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12688), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12176), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11722));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3316 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3317 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3318 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3319 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12400), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3320 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3321 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3322 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11349), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12220), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12400), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12036));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3323 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11316), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11349), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11376), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12153));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3324 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11277), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12629), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12121), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12311), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11316));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3325 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11242), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12597), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12085), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11277));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3326 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[19]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[18]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12056), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11856), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12597));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3327 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8547), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3328 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8645), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3329 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8352), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3330 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8694), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8645), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8352), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3331 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8694));
NAND4BBXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3332 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7943), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8547), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7680));
AND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3333 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8464), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3334 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[1]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8464), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3335 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12204), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11816), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12449), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11272), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11468));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3336 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11203), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12047), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12768), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12239));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3337 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[20]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11816), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11242), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12563));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3338 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[1]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[19]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3339 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7812), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3340 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8059), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7812), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3341 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3342 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8719), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7859));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3343 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8395), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8059), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8719), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3344 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8542), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3345 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3346 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7920), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3347 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[2]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8395), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8542), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7920));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3348 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43947), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11551), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11774), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12732), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12204));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3349 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[21]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11203), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12533), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11551));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3350 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[20]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[20]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3351 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14601), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3352 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7785), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3353 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8434), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3354 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8413), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8434));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3355 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8040), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8413), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3356 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8755), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3357 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3358 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8612), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7785), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8755), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8662));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3359 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8612));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3360 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43967), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43960), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43947), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43990));
ADDFHXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3361 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[21]), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[21]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3362 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3363 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14601), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847));
NOR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3364 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3365 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7916), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3366 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8734), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7916), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3367 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43949), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8734));
NAND4XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3368 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43993), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43963), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43949));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3369 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43967), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43993), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43973));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3370 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3371 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577));
NAND2X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3372 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14522), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3373 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3374 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3375 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3376 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3377 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11639), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3378 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3379 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3380 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11834), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3381 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11166), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12529), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12028), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11639), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11834));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3382 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12846), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12496), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11166), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11191), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11966));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3383 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3384 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3385 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3386 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12392), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3387 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11937), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11547), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12728), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12392));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3388 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3389 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12793), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3390 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3391 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11632), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3392 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12499), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12134), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12348), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12793), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11632));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3393 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3394 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3395 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3396 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3397 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12097), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3398 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11462), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3399 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3400 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11284), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3401 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12772), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12420), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12097), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11462), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11284));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3402 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11678), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11302), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11527), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12772), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12296));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3403 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11331), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12676), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12509), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11678), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11946));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3404 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11737), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11357), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12621), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11331), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3405 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12673), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12316), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12499), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11737), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11768));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3406 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11900), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11509), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12693), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11937), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12673));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3407 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12810), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12458), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12846), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11900));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3408 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[18]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12810), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12629), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11655));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3409 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8669), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3410 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8048), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435));
NOR3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3411 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8486), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8048));
NAND4BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3412 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7961), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8669), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8486), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3413 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8135), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3414 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8135));
NOR4BBX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3415 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8586), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371), .BN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8621));
NAND3BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3416 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[0]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7961), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8586));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3417 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[0]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3418 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14673), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[18]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3419 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3420 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14673), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3421 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3422 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11260), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3423 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3424 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11448), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3425 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3426 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11825), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3427 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11519), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12854), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11260), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11448), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11825));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3428 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3429 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12263), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3430 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12444), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3431 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3432 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3433 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11954), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11560), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12444), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11696));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3434 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3435 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12852), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3436 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11820), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11433), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12852), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12420));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3437 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11749), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3438 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12445), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11302), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11820), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11749));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3439 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12105), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11707), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12263), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12445), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12676));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3440 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3441 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12022), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3442 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12288), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11906), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12105), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12022), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11357));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3443 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11698), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11325), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12529), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11519), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12288));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3444 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12639), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12283), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12496), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11728), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11698));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3445 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[17]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[16]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12639), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11688), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12458));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3446 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[17]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3447 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3448 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12615), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3449 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3450 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12784), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3451 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3452 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11439), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3453 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11877), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11491), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12615), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12784), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11439));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3454 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3455 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11253), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3456 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3457 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12442), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3458 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3459 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12636), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3460 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3461 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12498), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3462 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3463 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12128), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3464 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11676), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3465 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3466 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11321), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3467 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12599), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12242), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12128), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11676), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11321));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3468 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12685), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12331), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12636), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12498), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12599));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3469 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12709), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3470 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12565), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11433), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12685), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12709));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3471 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11465), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12796), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12079), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12565), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3472 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12824), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12472), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11253), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12442), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11465));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3473 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11295), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12647), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12824), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12134));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3474 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12464), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11547), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12316));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3475 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[16]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[15]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12464), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11509), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12283));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3476 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14882), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[16]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3477 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11986), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3478 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11719), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11336), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12331), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11560), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11986));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3479 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3480 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11494), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3481 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11588), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11205), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12206), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11719), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11494));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3482 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3483 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3484 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11673), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3485 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3486 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12250), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3487 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3488 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3489 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11733), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3490 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11533), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12651), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11733));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3491 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3492 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12671), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3493 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3494 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11355), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3495 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11914), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3496 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12860), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3497 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3498 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3499 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12428), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12058), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12860), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12696));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3500 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11991), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11593), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11355), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11914), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12428));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3501 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12305), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11923), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12867), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12671), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11991));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3502 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11624), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11244), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12242), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11533), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12305));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3503 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12480), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12114), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11624), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11336));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3504 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12355), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12480), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12250), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11673));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3505 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12016), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11618), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11588), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12796), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12355));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3506 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11645), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11266), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11491), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12472), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12016));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3507 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3508 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12073), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3509 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3510 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11879), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3511 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3512 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3513 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12234), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11849), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12073), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11879), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12608));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3514 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3515 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12255), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3516 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44110), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3517 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44110));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3518 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3519 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12436), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3520 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3521 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12776), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3522 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11238), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12594), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12255), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12436), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12776));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3523 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12618), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12259), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11707), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12234), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11238));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3524 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12071), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11670), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12854), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11906));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3525 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[14]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11645), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12647), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11670));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3526 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[15]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[14]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11325), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12071), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12099));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3527 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[15]));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3528 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14534), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[14]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[14]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3529 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3530 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11486), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3531 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3532 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11663), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3533 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12271), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11887), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11486), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11663), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12114));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3534 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3535 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12826), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3536 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3537 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11861), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3538 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3539 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11299), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3540 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11498), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12833), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12826), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11861), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11299));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3541 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12140), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12271), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11498), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11983));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3542 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3543 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11869), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3544 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3545 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12064), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3546 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11361), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12708), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11869), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12064), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11205));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3547 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12735), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12385), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11361), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11849), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12594));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3548 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[12]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12140), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11618), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12385));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3549 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[13]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12735), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12259), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11266));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3550 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15031), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[12]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3551 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[13]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3552 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14627), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15031), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3553 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3554 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11309), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12662), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11923), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12208), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3555 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3556 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3557 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3558 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3559 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11399), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12743), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11309), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12649), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11290));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3560 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11209), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3561 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3562 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12473), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3563 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12391), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12023), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11244), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11209), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12473));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3564 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11273), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11399), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12391), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12833));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3565 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[11]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11273), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12708), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11745));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3566 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14777), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[11]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3567 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3568 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12820), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3569 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3570 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12290), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3571 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3572 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12109), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3573 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3574 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3575 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12088), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11684), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12290), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12109), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12641));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3576 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12175), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11783), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12023), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12820), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12088));
ADDFXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3577 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[10]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[9]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12175), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11887), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12625));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3578 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[10]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3579 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3580 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12465), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3581 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11435), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3582 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3583 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3584 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12716), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12364), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11435), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11593), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11711));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3585 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12806), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12452), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12662), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12465), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12716));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3586 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[9]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12743), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12806), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11783));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3587 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14853), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[9]));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3588 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14887), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14853));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3589 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12422), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3590 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11438), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12778), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12422), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12058), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3591 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3592 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11911), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3593 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3594 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12101), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3595 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11753), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11367), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11438), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12101), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11911));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3596 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[8]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11684), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11753), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12452));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3597 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14604), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[8]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[8]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3598 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3599 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3600 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3601 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11332), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3602 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3603 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11522), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3604 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12214), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11824), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11701), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11332), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11522));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3605 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[7]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12364), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11367));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3606 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14924), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[7]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3607 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3608 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3609 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12628), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3610 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12841), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12490), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12628), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3611 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3612 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12324), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3613 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3614 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12504), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3615 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11895), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12490), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12324), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12504));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3616 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[5]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12841), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11895));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3617 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11653), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3618 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12137), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3619 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3620 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3621 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12632), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11653), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12137), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12680));
ADDFX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3622 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[6]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12778), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12632), .CI(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11824));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3623 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[6]));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3624 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14623), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[5]), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[5]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3625 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14745), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3626 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3627 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3628 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11889), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3629 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12835), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3630 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11343), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12835), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]));
ADDHX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3631 (.CO(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[3]), .S(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11889), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11343));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3632 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[3]));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3633 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14733), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[2]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3634 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3635 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3636 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[1]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[1]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3637 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[2]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3638 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[3]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3639 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14615), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14697), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14944));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3640 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15041), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14733), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14690), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14615));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3641 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14625), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[4]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3642 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14572), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14745), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15041), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14625));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3643 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14871), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[5]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3644 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14551), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[6]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3645 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15069), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14871), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14551));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3646 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14529), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14623), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14572), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15069));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3647 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14797), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[7]));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3648 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14807), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14924), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14529), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14797));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3649 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15055), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[8]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[8]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3650 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15016), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14604), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14807), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15055));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3651 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14724), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[9]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3652 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14974), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[10]));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3653 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14940), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14724), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14974));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3654 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14763), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14940));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3655 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14751), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14887), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15016), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14763));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3656 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14658), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[11]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3657 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14565), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14751), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14777), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14658));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3658 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14904), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[12]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3659 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14582), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[13]));
AO21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3660 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15075), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14904), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14582));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3661 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15057), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14627), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14565), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15075));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3662 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14834), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[14]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3663 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15083), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[15]));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3664 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14977), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14834), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15083));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3665 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14965), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14534), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15057), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14977));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3666 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14756), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[16]));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3667 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14635), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14882), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14965), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14756));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3668 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14621), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14635));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3669 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14867), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[17]));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3670 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14992), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14621), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14867));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3671 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[18]));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3672 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14792), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3673 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14545), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14792));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3674 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3675 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15048), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3676 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14719), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3677 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15048), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14719));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3678 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14971), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3679 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14651), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3680 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14971), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14651));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3681 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3682 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3683 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14634), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3684 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3685 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628));
AOI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3686 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3687 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3688 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3689 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076));
OAI21X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3690 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3691 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3692 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3693 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3694 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3695 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3696 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3697 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3698 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3699 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3700 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3701 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3702 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3703 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3704 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3705 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3706 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3707 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14812), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3708 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14812));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3709 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3710 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3711 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3712 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3713 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3714 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3715 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14515), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3716 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14515));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3717 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3718 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3719 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3720 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3721 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3722 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14795), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3723 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14922), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14795));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3724 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15001), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14922));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3725 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14566), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15001));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3726 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14700), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14566));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3727 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837), .A0(N22593), .A1(N22531), .B0(N22648));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3728 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3729 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3730 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3731 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15006), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985));
AOI2BB1X4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3732 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43813), .A0N(N22536), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837), .B0(N22534));
CLKINVX8 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3733 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43813));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3734 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14738), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3735 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14543), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14738));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3736 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3737 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[48]), .A(N21801), .B(N23056), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3738 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22752), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[48]), .B(N21766));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3739 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22752));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3740 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219), .B(N19980));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3741 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14787), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3742 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3743 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3744 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14783), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3745 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808), .A0(N22562), .A1(N22564), .B0(N22566));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3746 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[28]), .A(N22489), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3747 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[28]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3748 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3749 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14826), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3750 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14703), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3751 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[29]), .A(N22385), .B(N22387), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3752 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[29]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3753 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3754 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14938), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3755 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14589), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14938));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3756 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15038), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3757 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3758 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14896), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3759 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14951), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3760 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14644), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3761 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14771), .A0(N22571), .A1(N22566), .B0(N22569));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3762 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908), .A0(N22644), .A1(N22504), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14771));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3763 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[40]), .A(N22404), .B(N22402), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3764 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[40]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3765 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3766 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3767 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14858), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3768 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14858), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3769 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14600), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3770 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14600));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3771 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14840), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3772 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[41]), .A(N22411), .B(N22409), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3773 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[41]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3774 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3775 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3776 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14760), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3777 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3778 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3779 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3780 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3781 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3782 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3783 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3784 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43441), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3785 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3786 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3787 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3788 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14610), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3789 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43426), .A(N22510));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3790 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3791 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3792 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15039), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3793 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3794 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14752), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3795 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14888), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14752));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3796 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43433), .A0(N22583), .A1(N22512), .B0(N22581));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3797 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585), .A0(N23029), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43426), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43433));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3798 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[43]), .A(N22368), .B(N22366), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3799 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[43]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3800 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14881), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3801 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[42]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585), .B(N22319));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3802 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[42]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3803 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3804 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3805 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14669), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3806 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[46]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837), .B(N22392));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3807 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[46]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3808 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3809 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14739), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3810 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14619), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3811 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[47]), .A(N22437), .B(N22439), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3812 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[47]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3813 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3814 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3815 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14555), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3816 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14564), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14555));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3817 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15014), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3818 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[44]), .A(N22451), .B(N22453), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3819 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[44]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3820 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3821 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14588), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3822 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14588));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3823 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3824 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43432), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3825 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43438), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3826 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43446), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43438));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3827 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3828 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43448), .A(N22332), .B(N22330), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3829 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43448));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3830 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3831 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3832 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3833 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3834 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3835 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14782), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3836 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14665), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3837 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[39]), .A(N22397), .B(N22395), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908));
NOR2BX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3838 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[39]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3839 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14528), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3840 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[38]), .A(N22361), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3841 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[38]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3842 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3843 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3844 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3845 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3846 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14557), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3847 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14982), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3848 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14980), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14982));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3849 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14859), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3850 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3851 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3852 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14649), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3853 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3854 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14830), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3855 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14537), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3856 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14959), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3857 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14521), .A0(N22600), .A1(N22520), .B0(N22598));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3858 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662), .A0(N22646), .A1(N22558), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14521));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3859 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44122), .A(N22484), .B(N22482), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3860 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[37]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44122));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3861 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[37]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3862 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3863 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14753), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3864 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14609), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14753));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3865 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15061), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3866 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[36]), .A(N22342), .B(N22344), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3867 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[36]));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3868 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3869 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3870 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3871 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43800), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3872 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43804), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3873 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43808), .A(N22349), .B(N22351), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3874 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43808));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3875 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43811), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3876 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43817), .A(N22373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3877 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43817));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3878 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3879 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14571), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3880 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063), .A0(N22524), .A1(N22526), .B0(N22528));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3881 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[32]), .A(N22416), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3882 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[32]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3883 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3884 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15000), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3885 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14877), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3886 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[33]), .A(N22430), .B(N22432), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3887 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[33]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3888 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3889 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3890 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3891 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3892 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14630), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3893 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15079), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3894 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929), .A0(N22508), .A1(N22510), .B0(N22512));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3895 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[31]), .A(N22356), .B(N22358), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3896 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[31]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3897 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14964), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3898 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[30]), .A(N22378), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3899 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[30]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NOR2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3900 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3901 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3902 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3903 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3904 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14652), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3905 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14525), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3906 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732), .A(N22531));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3907 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[25]), .A(N22444), .B(N22442), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3908 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[25]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3909 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15920), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0]));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3910 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14614), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949));
OA21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3911 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687), .A0(N22516), .A1(N22518), .B0(N22520));
XNOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3912 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[26]), .A(N22304), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3913 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[26]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3914 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3915 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15024), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986));
XNOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3916 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14899), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3917 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[27]), .A(N22423), .B(N22421), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3918 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[27]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3919 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15959), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3920 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15978), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15920), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15959));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3921 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15945), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3922 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15967), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15945));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3923 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15987), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3924 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15917), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15967), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15987));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3925 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15962), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15978), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15917));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3926 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15994), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3927 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15923), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3928 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15941), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15994), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15923));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3929 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15931), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3930 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15950), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3931 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15972), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15931), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15950));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3932 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15913), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15941), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15972));
AOI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3933 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15962), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15913));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3934 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15960), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3935 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15980), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3936 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15911), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15960), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15980));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3937 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15970), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3938 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15989), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15970), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3939 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15983), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22]));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3940 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15937), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15989), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15983));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3941 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15949), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15911), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15937));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3942 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15949));
OAI21X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3943 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3944 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[0]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541));
CLKINVX4 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3945 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[0]));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3946 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3947 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3948 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43353), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3949 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43361), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3950 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43346), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43353), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43361));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3951 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15982), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3952 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15928), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3953 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43367), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15982), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15928));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3954 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15938), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3955 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15958), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3956 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43337), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15938), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15958));
AOI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3957 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43706), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43367), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43337));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3958 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43345), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3959 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43715), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43345), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3960 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43706), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43715));
MXI2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3961 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[1]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43346), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542));
CLKINVX6 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3962 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[1]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3963 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3964 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0]));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3965 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3966 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3967 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43708), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3968 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43717), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926));
OAI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3969 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43689), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43708), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43717));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3970 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43696), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693));
OAI21X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3971 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43689), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43696));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3972 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43713), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542));
CLKXOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3973 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[2]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43713));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3974 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[2]));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3975 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3976 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3977 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3978 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3979 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16087), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3980 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16139), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16087), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3981 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3982 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3983 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3984 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3985 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16107), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16139), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3986 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16062), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3987 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969));
INVXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3988 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544));
OAI2BB1X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3989 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16062), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44129));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3990 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16063), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3991 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[4]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16063), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952));
INVX3 DFT_compute_cynw_cm_float_sin_E8_M23_1_I3992 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[4]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3993 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16170), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16107), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3994 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3995 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3996 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3997 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3998 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I3999 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4000 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4001 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16144), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4002 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16144), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4003 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16065), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4004 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16069), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16065));
XOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4005 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[3]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16069), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544));
INVX2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4006 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[3]));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4007 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N701), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16170), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4008 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N670), .A0(N23330), .A1(N20260), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N701));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4009 (.Y(x[22]), .A0(N23314), .A1(N23328), .B0(N23321), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N670));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4010 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4011 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4012 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4013 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4014 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4015 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4016 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4017 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16208), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4018 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16108), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16208), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4019 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4020 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4021 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4022 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16229), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16108), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4023 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16133), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16229), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4024 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4025 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4026 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4027 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MX2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4028 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4029 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4030 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16113), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4031 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16113), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4032 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N700), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16133), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4033 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584), .A0(N23335), .A1(N20547), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N700));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4034 (.Y(x[21]), .A0(N23316), .A1(N23328), .B0(N23323), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4035 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4036 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4037 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4038 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16230), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4039 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4040 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16195), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16230), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4041 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16099), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16195), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4042 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4043 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4044 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16234), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4045 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16234), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4046 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N699), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16099), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4047 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668), .A0(N23331), .A1(N20392), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N699));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4048 (.Y(x[20]), .A0(N23319), .A1(N23328), .B0(N23326), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4049 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4050 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4051 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16196), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4052 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4053 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16161), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16196), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4054 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16221), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16161), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4055 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4056 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4057 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16201), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4058 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16201), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4059 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N698), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16221), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4060 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667), .A0(N23332), .A1(N20454), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N698));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4061 (.Y(x[19]), .A0(N23318), .A1(N23328), .B0(N23325), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4062 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4063 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4064 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16124), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4065 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16189), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16124), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4066 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16166), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4067 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16166), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4068 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N697), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16189), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4069 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666), .A0(N23333), .A1(N20350), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N697));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4070 (.Y(x[18]), .A0(N23314), .A1(N23328), .B0(N23321), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4071 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4072 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16091), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4073 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16155), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16091), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4074 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16130), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4075 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16130), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4076 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N696), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16155), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4077 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665), .A0(N23336), .A1(N20537), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N696));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4078 (.Y(x[17]), .A0(N23315), .A1(N23328), .B0(N23322), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665));
NOR2BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4079 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4080 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16212), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4081 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16120), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16212), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4082 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16096), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4083 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16096), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4084 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N695), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16120), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4085 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664), .A0(N23330), .A1(N20444), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N695));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4086 (.Y(x[16]), .A0(N23318), .A1(N23328), .B0(N23325), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4087 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16181), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4088 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16207), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16181), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4089 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16218), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4090 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16218), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4091 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N694), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16207), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4092 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663), .A0(N23335), .A1(N20557), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N694));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4093 (.Y(x[15]), .A0(N23317), .A1(N23328), .B0(N23324), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4094 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4095 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N693), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4096 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662), .A0(N23331), .A1(N20414), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N693));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4097 (.Y(x[14]), .A0(N23317), .A1(N23328), .B0(N23324), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4098 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4099 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N692), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4100 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661), .A0(N23333), .A1(N20360), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N692));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4101 (.Y(x[13]), .A0(N23314), .A1(N23328), .B0(N23321), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4102 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4103 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N691), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4104 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660), .A0(N23335), .A1(N20434), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N691));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4105 (.Y(x[12]), .A0(N23319), .A1(N23328), .B0(N23326), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4106 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4107 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N690), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4108 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659), .A0(N23333), .A1(N20481), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N690));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4109 (.Y(x[11]), .A0(N23319), .A1(N23328), .B0(N23326), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4110 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4111 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N689), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4112 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658), .A0(N23334), .A1(N20471), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N689));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4113 (.Y(x[10]), .A0(N23316), .A1(N23328), .B0(N23323), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4114 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4115 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N688), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4116 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657), .A0(N23334), .A1(N20424), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N688));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4117 (.Y(x[9]), .A0(N23315), .A1(N23328), .B0(N23322), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4118 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4119 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N687), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4120 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656), .A0(N23333), .A1(N20587), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N687));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4121 (.Y(x[8]), .A0(N23319), .A1(N23328), .B0(N23326), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4122 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N686), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4123 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655), .A0(N23332), .A1(N20577), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N686));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4124 (.Y(x[7]), .A0(N23314), .A1(N23328), .B0(N23321), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4125 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N685), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4126 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654), .A0(N23334), .A1(N20370), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N685));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4127 (.Y(x[6]), .A0(N23317), .A1(N23328), .B0(N23324), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4128 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N684), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4129 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653), .A0(N23332), .A1(N20491), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N684));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4130 (.Y(x[5]), .A0(N23316), .A1(N23328), .B0(N23323), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4131 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N683), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4132 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652), .A0(N23330), .A1(N20567), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N683));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4133 (.Y(x[4]), .A0(N23317), .A1(N23328), .B0(N23324), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4134 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N682), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4135 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651), .A0(N23330), .A1(N20501), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N682));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4136 (.Y(x[3]), .A0(N23315), .A1(N23328), .B0(N23322), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4137 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N681), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4138 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650), .A0(N23334), .A1(N20597), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N681));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4139 (.Y(x[2]), .A0(N23316), .A1(N23328), .B0(N23323), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4140 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N680), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4141 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649), .A0(N23332), .A1(N20607), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N680));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4142 (.Y(x[1]), .A0(N23318), .A1(N23328), .B0(N23325), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4143 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N679), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4144 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648), .A0(N23331), .A1(N20617), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N679));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4145 (.Y(x[0]), .A0(N23318), .A1(N23328), .B0(N23325), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4146 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487));
AND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4147 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647), .A(a_exp[7]), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4148 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[30]), .A0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759), .A1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4149 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16468), .A0(N21461), .A1(N23333), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452));
NAND2BXL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4150 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426), .AN(N23330), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4151 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16468), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4152 (.Y(x[29]), .A0(N23319), .A1(N20199), .B0(N23326), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646));
AOI21XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4153 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16422), .A0(N21468), .A1(N23332), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4154 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16422), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4155 (.Y(x[28]), .A0(N23314), .A1(N20199), .B0(N23321), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645));
INVX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4156 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N675), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[4]));
AOI22X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4157 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16482), .A0(N21042), .A1(N23335), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N675));
NAND2X2 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4158 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16482));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4159 (.Y(x[27]), .A0(N23318), .A1(N20199), .B0(N23325), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4160 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16436), .A0(N21116), .A1(N23335), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[3]));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4161 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16436));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4162 (.Y(x[26]), .A0(N23315), .A1(N20199), .B0(N23322), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4163 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16391), .A0(N21231), .A1(N23331), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[2]));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4164 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16391));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4165 (.Y(x[25]), .A0(N23315), .A1(N20199), .B0(N23322), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4166 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16449), .A0(N21208), .A1(N23331), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4167 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16449));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4168 (.Y(x[24]), .A0(N23316), .A1(N20199), .B0(N23323), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641));
AOI22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4169 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16405), .A0(N21450), .A1(N23334), .B0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4170 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16405), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426));
AO22XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4171 (.Y(x[23]), .A0(N23317), .A1(N20199), .B0(N23324), .B1(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640));
OR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4172 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16540), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4173 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16578), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4174 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16560), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4175 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16547), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16578), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16560));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4176 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16545), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16540), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16547));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4177 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16570), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658));
NOR3XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4178 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16542), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4179 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16575), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16570), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16542));
OR4X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4180 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16530), .A(N20988), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640));
NOR3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4181 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16565), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16530));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4182 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16534), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4183 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16557), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16565), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16534));
NOR3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4184 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16576), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16557), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4185 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16568), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4186 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16535), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16576), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16568));
NOR3X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4187 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16556), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652));
NOR2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4188 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16572), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584));
NAND2X1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4189 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16558), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16556), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16572));
OR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4190 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16563), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16535), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16558));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4191 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16532), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16575), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16563));
NAND2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4192 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7297), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
NOR2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4193 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7297), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4194 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N577), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829), .B(a_sign), .S0(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757));
NOR3BX1 DFT_compute_cynw_cm_float_sin_E8_M23_1_I4195 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16612), .AN(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N577), .B(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487), .C(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82));
OAI2BB1XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4196 (.Y(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16607), .A0N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16545), .A1N(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16532), .B0(N20253));
MXI2XL DFT_compute_cynw_cm_float_sin_E8_M23_1_I4197 (.Y(x[31]), .A(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16607), .B(N19976), .S0(N23336));
EDFFHQX1 x_reg_30__I4228 (.Q(x[30]), .D(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[30]), .E(bdw_enable), .CK(aclk));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[0] = x[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[1] = x[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[2] = x[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[3] = x[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[4] = x[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[5] = x[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[6] = x[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[7] = x[7];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[8] = x[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[9] = x[9];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[10] = x[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[11] = x[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[12] = x[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[13] = x[13];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[14] = x[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[15] = x[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[16] = x[16];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[17] = x[17];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[18] = x[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[19] = x[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[20] = x[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[21] = x[21];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[22] = x[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[23] = x[23];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[24] = x[24];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[25] = x[25];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[26] = x[26];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[27] = x[27];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[28] = x[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[29] = x[29];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[31] = x[31];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[18] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[19] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[20] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[34] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[35] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[49] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[30] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urb1TQjeqhlA : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



