/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:21:38 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__21,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire  inst_cellmath__46;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__66,
	inst_cellmath__67,
	inst_cellmath__68,
	inst_cellmath__69,
	inst_cellmath__82;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [20:0] inst_cellmath__197;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__200,
	inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire  inst_cellmath__219;
wire N491,N492,N493,N494,N548,N549,N550 
	,N551,N552,N583,N585,N594,N595,N597,N598 
	,N599,N600,N601,N602,N603,N604,N605,N606 
	,N607,N608,N609,N610,N611,N612,N613,N614 
	,N615,N616,N617,N618,N619,N620,N621,N622 
	,N623,N624,N625,N626,N627,N628,N629,N630 
	,N631,N632,N633,N634,N635,N636,N637,N638 
	,N639,N640,N641,N642,N643,N644,N645,N646 
	,N647,N648,N649,N650,N651,N652,N653,N654 
	,N655,N656,N657,N658,N659,N661,N662,N663 
	,N664,N665,N666,N667,N668,N669,N670,N671 
	,N672,N673,N674,N675,N676,N677,N678,N679 
	,N680,N681,N682,N683,N684,N685,N686,N687 
	,N688,N689,N690,N691,N692,N693,N694,N695 
	,N696,N697,N698,N699,N700,N701,N702,N703 
	,N704,N705,N706,N707,N708,N709,N710,N711 
	,N712,N713,N714,N715,N716,N717,N718,N719 
	,N720,N721,N722,N723,N724,N725,N726,N727 
	,N728,N729,N730,N731,N732,N733,N734,N735 
	,N736,N737,N738,N739,N741,N742,N743,N744 
	,N745,N746,N747,N748,N749,N750,N751,N752 
	,N753,N754,N755,N756,N757,N758,N759,N760 
	,N761,N762,N763,N764,N3807,N3808,N3809,N3810 
	,N3815,N3816;
cynw_cm_float_cos_inst_blk01_cellmath__39_bdw1157874770_bdw cynw_cm_float_cos_I0 (.inst_blk01_cellmath__39_out0({N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597}), .inst_blk01_cellmath__39_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_cos_inst_cellmath__42_0_bdw1157874770_bdw cynw_cm_float_cos_I1 (.inst_cellmath__42_0_out0({inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6], inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__42_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__48_bdw1157874770_bdw cynw_cm_float_cos_I2 (.inst_cellmath__48_out0({N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684}), .inst_cellmath__48_in0({inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__48_in1({N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623}));
cynw_cm_float_cos_inst_cellmath__58__24__bdw1157874770_bdw cynw_cm_float_cos_I3 (.inst_cellmath__58__24__out0({N493, N492}), .inst_cellmath__58__24__in0({N708, N707}));
cynw_cm_float_cos_inst_cellmath__61_0_bdw1157874770_bdw cynw_cm_float_cos_I4 (.inst_cellmath__61_0_out0({inst_cellmath__61[22], inst_cellmath__61[21], inst_cellmath__61[20], inst_cellmath__61[19], inst_cellmath__61[18], inst_cellmath__61[17], inst_cellmath__61[16], inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__61_0_in0({N492}), .inst_cellmath__61_0_in1({N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684}));
INVXL cynw_cm_float_cos_I360 (.Y(N3807), .A(inst_cellmath__61[6]));
INVXL cynw_cm_float_cos_I361 (.Y(N3808), .A(N3807));
INVXL cynw_cm_float_cos_I362 (.Y(N3809), .A(inst_cellmath__61[10]));
INVXL cynw_cm_float_cos_I363 (.Y(N3810), .A(N3809));
INVXL cynw_cm_float_cos_I5 (.Y(inst_cellmath__115__W1[0]), .A(inst_cellmath__61[16]));
cynw_cm_float_cos_inst_cellmath__195__80__2WWMM_2WWMM_bdw1157874770_bdw cynw_cm_float_cos_I6 (.inst_cellmath__195__80__2WWMM_2WWMM_out0({inst_cellmath__195[29], inst_cellmath__195[28], inst_cellmath__195[27], inst_cellmath__195[26], inst_cellmath__195[25], inst_cellmath__195[24], inst_cellmath__195[23], inst_cellmath__195[22], inst_cellmath__195[21], inst_cellmath__195[20], inst_cellmath__195[19], inst_cellmath__195[18], inst_cellmath__195[17], inst_cellmath__195[16], inst_cellmath__195[15], inst_cellmath__195[14], inst_cellmath__195[13], inst_cellmath__195[12], inst_cellmath__195[11], inst_cellmath__195[10], inst_cellmath__195[9], inst_cellmath__195[8], inst_cellmath__195[7], inst_cellmath__195[6], inst_cellmath__195[5], inst_cellmath__195[4], inst_cellmath__195[3], inst_cellmath__195[2], inst_cellmath__195[1], inst_cellmath__195[0], inst_cellmath__197[19], inst_cellmath__197[18], inst_cellmath__197[17], inst_cellmath__197[16], inst_cellmath__197[15], inst_cellmath__197[14], inst_cellmath__197[13], inst_cellmath__197[12], inst_cellmath__197[11], inst_cellmath__197[10], inst_cellmath__197[9], inst_cellmath__197[8], inst_cellmath__197[7], inst_cellmath__197[6], inst_cellmath__197[5], inst_cellmath__197[4], inst_cellmath__197[3], inst_cellmath__197[2], inst_cellmath__197[1], inst_cellmath__197[0], N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742}), .inst_cellmath__195__80__2WWMM_2WWMM_in0({inst_cellmath__61[22], inst_cellmath__61[21], inst_cellmath__61[20], inst_cellmath__61[19], inst_cellmath__61[18], inst_cellmath__61[17]}));
cynw_cm_float_cos_inst_cellmath__198_0_bdw1157874770_bdw cynw_cm_float_cos_I7 (.inst_cellmath__198_0_out0({inst_cellmath__198[32], inst_cellmath__198[31], inst_cellmath__198[30], inst_cellmath__198[29], inst_cellmath__198[28], inst_cellmath__198[27], inst_cellmath__198[26], inst_cellmath__198[25], inst_cellmath__198[24], inst_cellmath__198[23], inst_cellmath__198[22], inst_cellmath__198[21], inst_cellmath__198[20], inst_cellmath__198[19], inst_cellmath__198[18], inst_cellmath__198[17], inst_cellmath__198[16], inst_cellmath__198[15], inst_cellmath__198[14], inst_cellmath__198[13], inst_cellmath__198[12], inst_cellmath__198[11], inst_cellmath__198[10], inst_cellmath__198[9], inst_cellmath__198[8], inst_cellmath__198[7], inst_cellmath__198[6], inst_cellmath__198[5], inst_cellmath__198[4], inst_cellmath__198[3], inst_cellmath__198[2], inst_cellmath__198[1], inst_cellmath__198[0]}), .inst_cellmath__198_0_in0({inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__198_0_in1({inst_cellmath__115__W1[0]}));
cynw_cm_float_cos_inst_cellmath__203_0_bdw1157874770_bdw cynw_cm_float_cos_I8 (.inst_cellmath__203_0_out0({inst_cellmath__203__W1[46], inst_cellmath__203__W1[45], inst_cellmath__203__W1[44], inst_cellmath__203__W1[43], inst_cellmath__203__W1[42], inst_cellmath__203__W1[41], inst_cellmath__203__W1[40], inst_cellmath__203__W1[39], inst_cellmath__203__W1[38], inst_cellmath__203__W1[37], inst_cellmath__203__W1[36], inst_cellmath__203__W1[35], inst_cellmath__203__W1[34], inst_cellmath__203__W1[33], inst_cellmath__203__W1[32], inst_cellmath__203__W1[31], inst_cellmath__203__W1[30], inst_cellmath__203__W1[29], inst_cellmath__203__W1[28], inst_cellmath__203__W1[27], inst_cellmath__203__W1[26], inst_cellmath__203__W1[25], inst_cellmath__203__W1[24], inst_cellmath__203__W1[23], inst_cellmath__203__W1[22], inst_cellmath__203__W1[21], inst_cellmath__203__W1[20], inst_cellmath__203__W1[19], inst_cellmath__203__W1[18], inst_cellmath__203__W1[17], inst_cellmath__203__W1[16], inst_cellmath__203__W1[15], inst_cellmath__203__W1[14], inst_cellmath__203__W1[13], inst_cellmath__203__W1[12], inst_cellmath__203__W1[11], inst_cellmath__203__W1[10], inst_cellmath__203__W1[9], inst_cellmath__203__W1[8], inst_cellmath__203__W1[7], inst_cellmath__203__W1[6], inst_cellmath__203__W1[5], inst_cellmath__203__W1[4], inst_cellmath__203__W1[3], inst_cellmath__203__W1[2], inst_cellmath__203__W1[1], inst_cellmath__203__W1[0]}), .inst_cellmath__203_0_out1({inst_cellmath__203__W0[46], inst_cellmath__203__W0[45], inst_cellmath__203__W0[44], inst_cellmath__203__W0[43], inst_cellmath__203__W0[42], inst_cellmath__203__W0[41], inst_cellmath__203__W0[40], inst_cellmath__203__W0[39], inst_cellmath__203__W0[38], inst_cellmath__203__W0[37], inst_cellmath__203__W0[36], inst_cellmath__203__W0[35], inst_cellmath__203__W0[34], inst_cellmath__203__W0[33], inst_cellmath__203__W0[32], inst_cellmath__203__W0[31], inst_cellmath__203__W0[30], inst_cellmath__203__W0[29], inst_cellmath__203__W0[28], inst_cellmath__203__W0[27], inst_cellmath__203__W0[26], inst_cellmath__203__W0[25], inst_cellmath__203__W0[24], inst_cellmath__203__W0[23], inst_cellmath__203__W0[22], inst_cellmath__203__W0[21], inst_cellmath__203__W0[20], inst_cellmath__203__W0[19], inst_cellmath__203__W0[18], inst_cellmath__203__W0[17], inst_cellmath__203__W0[16], inst_cellmath__203__W0[15], inst_cellmath__203__W0[14], inst_cellmath__203__W0[13], inst_cellmath__203__W0[12], inst_cellmath__203__W0[11], inst_cellmath__203__W0[10], inst_cellmath__203__W0[9], inst_cellmath__203__W0[8], inst_cellmath__203__W0[7], inst_cellmath__203__W0[6], inst_cellmath__203__W0[5], inst_cellmath__203__W0[4], inst_cellmath__203__W0[3], inst_cellmath__203__W0[2], inst_cellmath__203__W0[1], inst_cellmath__203__W0[0]}), .inst_cellmath__203_0_in0({inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], N3810, inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], N3808, inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__203_0_in1({inst_cellmath__198[32], inst_cellmath__198[31], inst_cellmath__198[30], inst_cellmath__198[29], inst_cellmath__198[28], inst_cellmath__198[27], inst_cellmath__198[26], inst_cellmath__198[25], inst_cellmath__198[24], inst_cellmath__198[23], inst_cellmath__198[22], inst_cellmath__198[21], inst_cellmath__198[20], inst_cellmath__198[19], inst_cellmath__198[18], inst_cellmath__198[17]}), .inst_cellmath__203_0_in2({inst_cellmath__197[19], inst_cellmath__197[18], inst_cellmath__197[17], inst_cellmath__197[16], inst_cellmath__197[15], inst_cellmath__197[14], inst_cellmath__197[13], inst_cellmath__197[12], inst_cellmath__197[11], inst_cellmath__197[10], inst_cellmath__197[9], inst_cellmath__197[8], inst_cellmath__197[7], inst_cellmath__197[6], inst_cellmath__197[5], inst_cellmath__197[4], inst_cellmath__197[3], inst_cellmath__197[2], inst_cellmath__197[1], inst_cellmath__197[0]}), .inst_cellmath__203_0_in3({N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742}), .inst_cellmath__203_0_in4({inst_cellmath__115__W1[0]}));
cynw_cm_float_cos_inst_cellmath__201_0_bdw1157874770_bdw cynw_cm_float_cos_I9 (.inst_cellmath__201_0_out0({inst_cellmath__201[49], inst_cellmath__201[48], inst_cellmath__201[47], inst_cellmath__201[46], inst_cellmath__201[45], inst_cellmath__201[44], inst_cellmath__201[43], inst_cellmath__201[42], inst_cellmath__201[41], inst_cellmath__201[40], inst_cellmath__201[39], inst_cellmath__201[38], inst_cellmath__201[37], inst_cellmath__201[36], inst_cellmath__201[35], inst_cellmath__201[34], inst_cellmath__201[33], inst_cellmath__201[32], inst_cellmath__201[31], inst_cellmath__201[30], inst_cellmath__201[29], inst_cellmath__201[28], inst_cellmath__201[27], inst_cellmath__201[26], inst_cellmath__201[25], inst_cellmath__201[24], inst_cellmath__201[23], inst_cellmath__201[22], inst_cellmath__201[21], inst_cellmath__201[20], inst_cellmath__201[19], inst_cellmath__201[18], inst_cellmath__201[17], inst_cellmath__201[16], inst_cellmath__201[15], inst_cellmath__201[14], inst_cellmath__201[13], inst_cellmath__201[12], inst_cellmath__201[11], inst_cellmath__201[10], inst_cellmath__201[9], inst_cellmath__201[8], inst_cellmath__201[7], inst_cellmath__201[6], inst_cellmath__201[5], inst_cellmath__201[4], inst_cellmath__201[3], inst_cellmath__201[2], inst_cellmath__201[1], inst_cellmath__201[0]}), .inst_cellmath__201_0_in0({inst_cellmath__203__W1[46], inst_cellmath__203__W1[45], inst_cellmath__203__W1[44], inst_cellmath__203__W1[43], inst_cellmath__203__W1[42], inst_cellmath__203__W1[41], inst_cellmath__203__W1[40], inst_cellmath__203__W1[39], inst_cellmath__203__W1[38], inst_cellmath__203__W1[37], inst_cellmath__203__W1[36], inst_cellmath__203__W1[35], inst_cellmath__203__W1[34], inst_cellmath__203__W1[33], inst_cellmath__203__W1[32], inst_cellmath__203__W1[31], inst_cellmath__203__W1[30], inst_cellmath__203__W1[29], inst_cellmath__203__W1[28], inst_cellmath__203__W1[27], inst_cellmath__203__W1[26], inst_cellmath__203__W1[25], inst_cellmath__203__W1[24], inst_cellmath__203__W1[23], inst_cellmath__203__W1[22], inst_cellmath__203__W1[21], inst_cellmath__203__W1[20], inst_cellmath__203__W1[19], inst_cellmath__203__W1[18], inst_cellmath__203__W1[17], inst_cellmath__203__W1[16], inst_cellmath__203__W1[15], inst_cellmath__203__W1[14], inst_cellmath__203__W1[13], inst_cellmath__203__W1[12], inst_cellmath__203__W1[11], inst_cellmath__203__W1[10], inst_cellmath__203__W1[9], inst_cellmath__203__W1[8], inst_cellmath__203__W1[7], inst_cellmath__203__W1[6], inst_cellmath__203__W1[5], inst_cellmath__203__W1[4], inst_cellmath__203__W1[3], inst_cellmath__203__W1[2], inst_cellmath__203__W1[1], inst_cellmath__203__W1[0]}), .inst_cellmath__201_0_in1({inst_cellmath__203__W0[46], inst_cellmath__203__W0[45], inst_cellmath__203__W0[44], inst_cellmath__203__W0[43], inst_cellmath__203__W0[42], inst_cellmath__203__W0[41], inst_cellmath__203__W0[40], inst_cellmath__203__W0[39], inst_cellmath__203__W0[38], inst_cellmath__203__W0[37], inst_cellmath__203__W0[36], inst_cellmath__203__W0[35], inst_cellmath__203__W0[34], inst_cellmath__203__W0[33], inst_cellmath__203__W0[32], inst_cellmath__203__W0[31], inst_cellmath__203__W0[30], inst_cellmath__203__W0[29], inst_cellmath__203__W0[28], inst_cellmath__203__W0[27], inst_cellmath__203__W0[26], inst_cellmath__203__W0[25], inst_cellmath__203__W0[24], inst_cellmath__203__W0[23], inst_cellmath__203__W0[22], inst_cellmath__203__W0[21], inst_cellmath__203__W0[20], inst_cellmath__203__W0[19], inst_cellmath__203__W0[18], inst_cellmath__203__W0[17], inst_cellmath__203__W0[16], inst_cellmath__203__W0[15], inst_cellmath__203__W0[14], inst_cellmath__203__W0[13], inst_cellmath__203__W0[12], inst_cellmath__203__W0[11], inst_cellmath__203__W0[10], inst_cellmath__203__W0[9], inst_cellmath__203__W0[8], inst_cellmath__203__W0[7], inst_cellmath__203__W0[6], inst_cellmath__203__W0[5], inst_cellmath__203__W0[4], inst_cellmath__203__W0[3], inst_cellmath__203__W0[2], inst_cellmath__203__W0[1], inst_cellmath__203__W0[0]}), .inst_cellmath__201_0_in2({inst_cellmath__195[29], inst_cellmath__195[28], inst_cellmath__195[27], inst_cellmath__195[26], inst_cellmath__195[25], inst_cellmath__195[24], inst_cellmath__195[23], inst_cellmath__195[22], inst_cellmath__195[21], inst_cellmath__195[20], inst_cellmath__195[19], inst_cellmath__195[18], inst_cellmath__195[17], inst_cellmath__195[16], inst_cellmath__195[15], inst_cellmath__195[14], inst_cellmath__195[13], inst_cellmath__195[12], inst_cellmath__195[11], inst_cellmath__195[10], inst_cellmath__195[9], inst_cellmath__195[8], inst_cellmath__195[7], inst_cellmath__195[6], inst_cellmath__195[5], inst_cellmath__195[4], inst_cellmath__195[3], inst_cellmath__195[2], inst_cellmath__195[1], inst_cellmath__195[0]}));
cynw_cm_float_cos_inst_cellmath__200_0_bdw1157874770_bdw cynw_cm_float_cos_I10 (.inst_cellmath__200_0_out0({inst_cellmath__200[48], inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0], inst_cellmath__200[24], inst_cellmath__200[23], inst_cellmath__200[22], inst_cellmath__200[21], inst_cellmath__200[20], inst_cellmath__200[19], inst_cellmath__200[18], inst_cellmath__200[17], inst_cellmath__200[16], inst_cellmath__200[15], inst_cellmath__200[14], inst_cellmath__200[13], inst_cellmath__200[12], inst_cellmath__200[11], inst_cellmath__200[10], inst_cellmath__200[9], inst_cellmath__200[8], inst_cellmath__200[7], inst_cellmath__200[6], inst_cellmath__200[5], inst_cellmath__200[4], inst_cellmath__200[3], inst_cellmath__200[2], inst_cellmath__200[1], inst_cellmath__200[0]}), .inst_cellmath__200_0_in0({inst_cellmath__201[49], inst_cellmath__201[48], inst_cellmath__201[47], inst_cellmath__201[46], inst_cellmath__201[45], inst_cellmath__201[44], inst_cellmath__201[43], inst_cellmath__201[42], inst_cellmath__201[41], inst_cellmath__201[40], inst_cellmath__201[39], inst_cellmath__201[38], inst_cellmath__201[37], inst_cellmath__201[36], inst_cellmath__201[35], inst_cellmath__201[34], inst_cellmath__201[33], inst_cellmath__201[32], inst_cellmath__201[31], inst_cellmath__201[30], inst_cellmath__201[29], inst_cellmath__201[28], inst_cellmath__201[27], inst_cellmath__201[26], inst_cellmath__201[25], inst_cellmath__201[24], inst_cellmath__201[23], inst_cellmath__201[22], inst_cellmath__201[21], inst_cellmath__201[20], inst_cellmath__201[19], inst_cellmath__201[18], inst_cellmath__201[17], inst_cellmath__201[16], inst_cellmath__201[15], inst_cellmath__201[14], inst_cellmath__201[13], inst_cellmath__201[12], inst_cellmath__201[11], inst_cellmath__201[10], inst_cellmath__201[9], inst_cellmath__201[8], inst_cellmath__201[7], inst_cellmath__201[6], inst_cellmath__201[5], inst_cellmath__201[4], inst_cellmath__201[3], inst_cellmath__201[2], inst_cellmath__201[1], inst_cellmath__201[0]}));
cynw_cm_float_cos_inst_cellmath__17_0_bdw1157874770_bdw cynw_cm_float_cos_I11 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__46__15__bdw1157874770_bdw cynw_cm_float_cos_I12 (.inst_cellmath__46__15__out0({N491}), .inst_cellmath__46__15__in0({inst_cellmath__42[7], inst_cellmath__42[6]}));
cynw_cm_float_cos_inst_cellmath__46_0_bdw1157874770_bdw cynw_cm_float_cos_I13 (.inst_cellmath__46_0_out0(inst_cellmath__46), .inst_cellmath__46_0_in0({N491}), .inst_cellmath__46_0_in1({inst_cellmath__42[8]}));
cynw_cm_float_cos_inst_cellmath__21_0_bdw1157874770_bdw cynw_cm_float_cos_I14 (.inst_cellmath__21_0_out0(inst_cellmath__21), .inst_cellmath__21_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__83__62__bdw1157874770_bdw cynw_cm_float_cos_I15 (.inst_cellmath__83__62__out0({N494}), .inst_cellmath__83__62__in0(inst_cellmath__46), .inst_cellmath__83__62__in1(inst_cellmath__21), .inst_cellmath__83__62__in2(inst_cellmath__17));
cynw_cm_float_cos_inst_cellmath__19_0_bdw1157874770_bdw cynw_cm_float_cos_I16 (.inst_cellmath__19_0_out0(inst_cellmath__19), .inst_cellmath__19_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__24_0_bdw1157874770_bdw cynw_cm_float_cos_I17 (.inst_cellmath__24_0_out0(inst_cellmath__24), .inst_cellmath__24_0_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_cos_inst_cellmath__69_0_bdw1157874770_bdw cynw_cm_float_cos_I18 (.inst_cellmath__69_0_out0(inst_cellmath__69), .inst_cellmath__69_0_in0(inst_cellmath__24), .inst_cellmath__69_0_in1(inst_cellmath__19));
cynw_cm_float_cos_inst_cellmath__82_0_bdw1157874770_bdw cynw_cm_float_cos_I19 (.inst_cellmath__82_0_out0(inst_cellmath__82), .inst_cellmath__82_0_in0(inst_cellmath__69), .inst_cellmath__82_0_in1(inst_cellmath__19));
cynw_cm_float_cos_inst_cellmath__66_0_bdw1157874770_bdw cynw_cm_float_cos_I20 (.inst_cellmath__66_0_out0(inst_cellmath__66), .inst_cellmath__66_0_in0(inst_cellmath__24), .inst_cellmath__66_0_in1(inst_cellmath__19), .inst_cellmath__66_0_in2(a_sign));
cynw_cm_float_cos_inst_cellmath__67_0_bdw1157874770_bdw cynw_cm_float_cos_I21 (.inst_cellmath__67_0_out0(inst_cellmath__67), .inst_cellmath__67_0_in0(inst_cellmath__24), .inst_cellmath__67_0_in1(inst_cellmath__19), .inst_cellmath__67_0_in2(a_sign));
cynw_cm_float_cos_inst_cellmath__68_0_bdw1157874770_bdw cynw_cm_float_cos_I22 (.inst_cellmath__68_0_out0(inst_cellmath__68), .inst_cellmath__68_0_in0(inst_cellmath__67), .inst_cellmath__68_0_in1(inst_cellmath__66));
cynw_cm_float_cos_inst_cellmath__228__231__bdw1157874770_bdw cynw_cm_float_cos_I23 (.inst_cellmath__228__231__out0({N741}), .inst_cellmath__228__231__in0({N494}), .inst_cellmath__228__231__in1(inst_cellmath__82), .inst_cellmath__228__231__in2(inst_cellmath__68));
cynw_cm_float_cos_inst_cellmath__219_0_bdw1157874770_bdw cynw_cm_float_cos_I24 (.inst_cellmath__219_0_out0(inst_cellmath__219), .inst_cellmath__219_0_in0({inst_cellmath__61[22]}), .inst_cellmath__219_0_in1({inst_cellmath__200[48]}));
cynw_cm_float_cos_inst_cellmath__211__182__bdw1157874770_bdw cynw_cm_float_cos_I25 (.inst_cellmath__211__182__out0({N552, N551, N550, N549, N548}), .inst_cellmath__211__182__in0({inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0]}));
cynw_cm_float_cos_inst_cellmath__215_0_bdw1157874770_bdw cynw_cm_float_cos_I26 (.inst_cellmath__215_0_out0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}), .inst_cellmath__215_0_in0({N552, N551, N550, N549, N548}));
cynw_cm_float_cos_inst_cellmath__220__188__bdw1157874770_bdw cynw_cm_float_cos_I27 (.inst_cellmath__220__188__out0({N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661}), .inst_cellmath__220__188__in0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}), .inst_cellmath__220__188__in1({inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0]}));
cynw_cm_float_cos_inst_cellmath__221__195__bdw1157874770_bdw cynw_cm_float_cos_I28 (.inst_cellmath__221__195__out0({N659, N658, N657, N656, N655, N654, N653}), .inst_cellmath__221__195__in0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}));
cynw_cm_float_cos_inst_cellmath__220_2WWMM_bdw1157874770_bdw cynw_cm_float_cos_I29 (.inst_cellmath__220_2WWMM_out0({N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709}), .inst_cellmath__220_2WWMM_in0({N659, N658, N657, N656, N655, N654, N653}), .inst_cellmath__220_2WWMM_in1({N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661}), .inst_cellmath__220_2WWMM_in2(inst_cellmath__219));
INVXL cynw_cm_float_cos_I368 (.Y(N3815), .A(N733));
INVXL cynw_cm_float_cos_I369 (.Y(N3816), .A(N3815));
cynw_cm_float_cos_inst_cellmath__223__208__bdw1157874770_bdw cynw_cm_float_cos_I30 (.inst_cellmath__223__208__out0({N583}), .inst_cellmath__223__208__in0({N715, N714, N713, N712, N711, N710, N709}), .inst_cellmath__223__208__in1({N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717}));
cynw_cm_float_cos_inst_cellmath__223__199__bdw1157874770_bdw cynw_cm_float_cos_I31 (.inst_cellmath__223__199__out0({x[31]}), .inst_cellmath__223__199__in0(inst_cellmath__82), .inst_cellmath__223__199__in1({N493}), .inst_cellmath__223__199__in2({inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6]}), .inst_cellmath__223__199__in3({N583}));
cynw_cm_float_cos_inst_cellmath__224__213__bdw1157874770_bdw cynw_cm_float_cos_I32 (.inst_cellmath__224__213__out0({N585}), .inst_cellmath__224__213__in0({N494}), .inst_cellmath__224__213__in1(inst_cellmath__68));
cynw_cm_float_cos_inst_cellmath__224__212__bdw1157874770_bdw cynw_cm_float_cos_I33 (.inst_cellmath__224__212__out0({N595}), .inst_cellmath__224__212__in0(inst_cellmath__82), .inst_cellmath__224__212__in1({N585}));
cynw_cm_float_cos_inst_cellmath__225__215__bdw1157874770_bdw cynw_cm_float_cos_I34 (.inst_cellmath__225__215__out0({N594}), .inst_cellmath__225__215__in0(inst_cellmath__82), .inst_cellmath__225__215__in1(inst_cellmath__68));
cynw_cm_float_cos_inst_cellmath__228_0_bdw1157874770_bdw cynw_cm_float_cos_I35 (.inst_cellmath__228_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__228_0_in0({N741}), .inst_cellmath__228_0_in1({N594}), .inst_cellmath__228_0_in2({N595}), .inst_cellmath__228_0_in3({N715, N714, N713, N712, N711, N710, N709}));
cynw_cm_float_cos_inst_cellmath__231_0_bdw1157874770_bdw cynw_cm_float_cos_I36 (.inst_cellmath__231_0_out0({x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__231_0_in0(inst_cellmath__82), .inst_cellmath__231_0_in1({N741}), .inst_cellmath__231_0_in2({N739, N738, N737, N736, N735, N734, N3816, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717}), .inst_cellmath__231_0_in3({inst_cellmath__210[21]}));
assign inst_cellmath__197[20] = 1'B1;
assign inst_cellmath__200[25] = inst_cellmath__210[0];
assign inst_cellmath__200[26] = inst_cellmath__210[1];
assign inst_cellmath__200[27] = inst_cellmath__210[2];
assign inst_cellmath__200[28] = inst_cellmath__210[3];
assign inst_cellmath__200[29] = inst_cellmath__210[4];
assign inst_cellmath__200[30] = inst_cellmath__210[5];
assign inst_cellmath__200[31] = inst_cellmath__210[6];
assign inst_cellmath__200[32] = inst_cellmath__210[7];
assign inst_cellmath__200[33] = inst_cellmath__210[8];
assign inst_cellmath__200[34] = inst_cellmath__210[9];
assign inst_cellmath__200[35] = inst_cellmath__210[10];
assign inst_cellmath__200[36] = inst_cellmath__210[11];
assign inst_cellmath__200[37] = inst_cellmath__210[12];
assign inst_cellmath__200[38] = inst_cellmath__210[13];
assign inst_cellmath__200[39] = inst_cellmath__210[14];
assign inst_cellmath__200[40] = inst_cellmath__210[15];
assign inst_cellmath__200[41] = inst_cellmath__210[16];
assign inst_cellmath__200[42] = inst_cellmath__210[17];
assign inst_cellmath__200[43] = inst_cellmath__210[18];
assign inst_cellmath__200[44] = inst_cellmath__210[19];
assign inst_cellmath__200[45] = inst_cellmath__210[20];
assign inst_cellmath__200[46] = inst_cellmath__210[21];
assign inst_cellmath__200[47] = inst_cellmath__210[22];
assign inst_cellmath__200[49] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_blk01_cellmath__39_bdw1157874770_bdw (
	inst_blk01_cellmath__39_out0,
	inst_blk01_cellmath__39_in0
	); /* architecture "gate_level" */ 
output [55:0] inst_blk01_cellmath__39_out0;
input [22:0] inst_blk01_cellmath__39_in0;
wire N354,N360,N362,N366,N368,N370,N372 
	,N374,N376,N378,N380,N382,N384,N386,N388 
	,N390,N392,N394,N396,N1066,N1067,N1070,N1071 
	,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079 
	,N1082,N1083,N1084,N1085,N1088,N1089,N1090,N1091 
	,N1094,N1095,N1096,N1097,N1098,N1099,N1102,N1103 
	,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111 
	,N1114,N1115,N1116,N1117,N1118,N1119,N1122,N1123 
	,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131 
	,N1132,N1133,N1136,N1137,N1138,N1139,N1140,N1141 
	,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149 
	,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157 
	,N1158,N1159,N1160,N1161,N1162,N1163,N1166,N1167 
	,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177 
	,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185 
	,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193 
	,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201 
	,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209 
	,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217 
	,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225 
	,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233 
	,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241 
	,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249 
	,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257 
	,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265 
	,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273 
	,N1274,N1275,N1278,N1279,N1282,N1283,N1286,N1287 
	,N1294,N1295,N1298,N1299,N1300,N1301,N1302,N1303 
	,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311 
	,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319 
	,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327 
	,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335 
	,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343 
	,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351 
	,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359 
	,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367 
	,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375 
	,N1376,N1377,N1378,N1379,N1380,N1381,N1384,N1385 
	,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393 
	,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401 
	,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409 
	,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417 
	,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425 
	,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433 
	,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441 
	,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449 
	,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457 
	,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465 
	,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473 
	,N1474,N1475,N1476,N1477,N1482,N1483,N1484,N1485 
	,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493 
	,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501 
	,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1511 
	,N1521,N1531,N1535,N1536,N1547,N1561,N1565,N1566 
	,N1583,N1611,N1613,N1617,N1618,N1621,N1622,N1661 
	,N1663,N1665,N1684,N1687,N1690,N1693,N1696,N1699 
	,N1702,N1705,N1708,N1711,N1714,N1717,N1734,N1736 
	,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744 
	,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752 
	,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760 
	,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768 
	,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776 
	,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784 
	,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792 
	,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800 
	,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808 
	,N1809,N1810,N1811,N1814,N1818,N1819,N1826,N1830 
	,N1831,N1834,N1835,N1842,N1843,N1846,N1847,N1850 
	,N1851,N1858,N1859,N1862,N1863,N1866,N1867,N1874 
	,N1875,N1878,N1879,N1882,N1883,N1890,N1891,N1894 
	,N1895,N1898,N1899,N1906,N1907,N1910,N1911,N1914 
	,N1915,N1922,N1923,N1926,N1927,N1930,N1931,N1938 
	,N1939,N1942,N1943,N1946,N1947,N1952,N1953,N1954 
	,N1955,N1964,N1966,N1968,N1974,N1975,N2002,N2004 
	,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012 
	,N2013,N2014,N2015,N2020,N2022,N2024,N2025,N2026 
	,N2027,N2028,N2029,N2030,N2031,N2040,N2042,N2044 
	,N2046,N2154,N2157,N2160,N2163,N2166,N2175,N2178 
	,N2187,N2190,N2199,N2202,N2211,N2214,N2223,N2226 
	,N2235,N2238,N2259,N2262,N2278,N2279,N2281,N2282 
	,N2284,N2285,N2287,N2288,N2290,N2291,N2293,N2294 
	,N2296,N2297,N2299,N2300,N2302,N2303,N2305,N2306 
	,N2308,N2309,N2311,N2312,N2314,N2315,N2317,N2318 
	,N2320,N2321,N2323,N2324,N2326,N2327,N2329,N2330 
	,N2332,N2333,N2335,N2336,N2338,N2339,N2341,N2342 
	,N2344,N2345,N2347,N2348,N2350,N2351,N2353,N2354 
	,N2356,N2357,N2583,N2599,N2601,N2610,N2612,N2628 
	,N2630,N2639,N2641,N2657,N2659,N2668,N2670,N2686 
	,N2688,N2697,N2699,N2715,N2717,N2726,N2728,N2744 
	,N2746,N2755,N2757,N2773,N2775,N2784,N2786,N2795 
	,N2797,N2806,N2808,N2817,N2819,N2828,N2830,N2846 
	,N2848,N3018,N3022,N3024,N3069,N3070,N3075,N3078 
	,N3087,N3092,N3093,N3096,N3098,N3099,N3113,N3121 
	,N3131,N3141,N3151,N3159,N3167,N3174,N3175,N3178 
	,N3179,N3191,N3210,N3211,N3212,N3213,N3214,N3215 
	,N3216,N3217,N3218,N3223,N3228,N3234,N3240,N3246 
	,N3252,N3258,N3264,N3266,N3278,N3279,N3282,N3289 
	,N3296,N3303,N3310,N3317,N3324,N3331,N3338,N3345 
	,N3352,N5103;
INVX2 inst_blk01_cellmath__39_I5 (.Y(N1482), .A(inst_blk01_cellmath__39_in0[0]));
CLKINVX12 inst_blk01_cellmath__39_I6 (.Y(N354), .A(inst_blk01_cellmath__39_in0[1]));
CLKINVX4 inst_blk01_cellmath__39_I7 (.Y(N1484), .A(inst_blk01_cellmath__39_in0[2]));
CLKINVX4 inst_blk01_cellmath__39_I8 (.Y(N1381), .A(inst_blk01_cellmath__39_in0[3]));
CLKINVX6 inst_blk01_cellmath__39_I9 (.Y(N360), .A(inst_blk01_cellmath__39_in0[4]));
CLKINVX6 inst_blk01_cellmath__39_I10 (.Y(N362), .A(inst_blk01_cellmath__39_in0[5]));
CLKINVX16 inst_blk01_cellmath__39_I11 (.Y(N1295), .A(inst_blk01_cellmath__39_in0[6]));
CLKINVX6 inst_blk01_cellmath__39_I12 (.Y(N366), .A(inst_blk01_cellmath__39_in0[7]));
INVX3 inst_blk01_cellmath__39_I13 (.Y(N368), .A(inst_blk01_cellmath__39_in0[8]));
CLKINVX4 inst_blk01_cellmath__39_I14 (.Y(N370), .A(inst_blk01_cellmath__39_in0[9]));
CLKINVX8 inst_blk01_cellmath__39_I15 (.Y(N372), .A(inst_blk01_cellmath__39_in0[10]));
INVX2 inst_blk01_cellmath__39_I16 (.Y(N374), .A(inst_blk01_cellmath__39_in0[11]));
INVX2 inst_blk01_cellmath__39_I17 (.Y(N376), .A(inst_blk01_cellmath__39_in0[12]));
INVX3 inst_blk01_cellmath__39_I18 (.Y(N378), .A(inst_blk01_cellmath__39_in0[13]));
INVX3 inst_blk01_cellmath__39_I19 (.Y(N380), .A(inst_blk01_cellmath__39_in0[14]));
INVXL inst_blk01_cellmath__39_I20 (.Y(N382), .A(inst_blk01_cellmath__39_in0[15]));
BUFX2 inst_blk01_cellmath__39_I1836 (.Y(N3018), .A(N382));
INVX2 inst_blk01_cellmath__39_I21 (.Y(N384), .A(inst_blk01_cellmath__39_in0[16]));
INVX3 inst_blk01_cellmath__39_I22 (.Y(N386), .A(inst_blk01_cellmath__39_in0[17]));
INVX2 inst_blk01_cellmath__39_I23 (.Y(N388), .A(inst_blk01_cellmath__39_in0[18]));
INVX2 inst_blk01_cellmath__39_I24 (.Y(N390), .A(inst_blk01_cellmath__39_in0[19]));
INVXL inst_blk01_cellmath__39_I25 (.Y(N392), .A(inst_blk01_cellmath__39_in0[20]));
BUFX2 inst_blk01_cellmath__39_I1837 (.Y(N3022), .A(N392));
INVX2 inst_blk01_cellmath__39_I26 (.Y(N394), .A(inst_blk01_cellmath__39_in0[21]));
INVXL inst_blk01_cellmath__39_I27 (.Y(N396), .A(inst_blk01_cellmath__39_in0[22]));
BUFX2 inst_blk01_cellmath__39_I1838 (.Y(N3024), .A(N396));
XNOR2X1 hap1_A_I1412 (.Y(N1066), .A(inst_blk01_cellmath__39_in0[9]), .B(inst_blk01_cellmath__39_in0[2]));
OR2XL hap1_A_I1413 (.Y(N1067), .A(inst_blk01_cellmath__39_in0[9]), .B(inst_blk01_cellmath__39_in0[2]));
ADDFX1 inst_blk01_cellmath__39_I332 (.CO(N1071), .S(N1070), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[10]), .CI(N354));
ADDFXL inst_blk01_cellmath__39_I333 (.CO(N1073), .S(N1072), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[11]), .CI(N1484));
ADDFX1 inst_blk01_cellmath__39_I334 (.CO(N1075), .S(N1074), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[12]), .CI(N1381));
ADDFX1 inst_blk01_cellmath__39_I335 (.CO(N1077), .S(N1076), .A(inst_blk01_cellmath__39_in0[6]), .B(inst_blk01_cellmath__39_in0[13]), .CI(N360));
XNOR2X1 hap1_A_I1414 (.Y(N1078), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[7]));
OR2XL hap1_A_I1415 (.Y(N1079), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[7]));
ADDHX1 inst_blk01_cellmath__39_I337 (.CO(N1083), .S(N1082), .A(N1482), .B(N362));
XNOR2X1 hap1_A_I1416 (.Y(N1084), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[8]));
OR2XL hap1_A_I1417 (.Y(N1085), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[8]));
ADDFHXL inst_blk01_cellmath__39_I339 (.CO(N1089), .S(N1088), .A(N1295), .B(N354), .CI(N372));
XNOR2X1 hap1_A_I1418 (.Y(N1090), .A(inst_blk01_cellmath__39_in0[16]), .B(inst_blk01_cellmath__39_in0[9]));
OR2XL hap1_A_I1419 (.Y(N1091), .A(inst_blk01_cellmath__39_in0[16]), .B(inst_blk01_cellmath__39_in0[9]));
ADDFX1 inst_blk01_cellmath__39_I341 (.CO(N1095), .S(N1094), .A(N1484), .B(inst_blk01_cellmath__39_in0[0]), .CI(N366));
ADDHX1 inst_blk01_cellmath__39_I342 (.CO(N1097), .S(N1096), .A(N374), .B(N396));
XNOR2X1 hap1_A_I1420 (.Y(N1098), .A(inst_blk01_cellmath__39_in0[17]), .B(inst_blk01_cellmath__39_in0[10]));
OR2XL hap1_A_I1421 (.Y(N1099), .A(inst_blk01_cellmath__39_in0[17]), .B(inst_blk01_cellmath__39_in0[10]));
ADDFXL inst_blk01_cellmath__39_I344 (.CO(N1103), .S(N1102), .A(N368), .B(inst_blk01_cellmath__39_in0[1]), .CI(N1381));
ADDHX1 inst_blk01_cellmath__39_I345 (.CO(N1105), .S(N1104), .A(N376), .B(N392));
ADDFX1 inst_blk01_cellmath__39_I346 (.CO(N1107), .S(N1106), .A(inst_blk01_cellmath__39_in0[11]), .B(inst_blk01_cellmath__39_in0[18]), .CI(inst_blk01_cellmath__39_in0[2]));
ADDFXL inst_blk01_cellmath__39_I347 (.CO(N1109), .S(N1108), .A(N370), .B(N360), .CI(N378));
XNOR2X1 hap1_A_I1422 (.Y(N1110), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[12]));
OR2XL hap1_A_I1423 (.Y(N1111), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[12]));
ADDFHXL inst_blk01_cellmath__39_I349 (.CO(N1115), .S(N1114), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[0]), .CI(N362));
ADDHX1 inst_blk01_cellmath__39_I350 (.CO(N1117), .S(N1116), .A(N372), .B(N380));
XNOR2X1 hap1_A_I1424 (.Y(N1118), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[13]));
OR2XL hap1_A_I1425 (.Y(N1119), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[13]));
ADDFX1 inst_blk01_cellmath__39_I352 (.CO(N1123), .S(N1122), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[1]), .CI(N1295));
ADDHX1 inst_blk01_cellmath__39_I353 (.CO(N1125), .S(N1124), .A(N374), .B(N382));
ADDFX1 inst_blk01_cellmath__39_I354 (.CO(N1127), .S(N1126), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[21]), .CI(inst_blk01_cellmath__39_in0[0]));
ADDFX1 inst_blk01_cellmath__39_I355 (.CO(N1129), .S(N1128), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[2]), .CI(N366));
ADDHX1 inst_blk01_cellmath__39_I356 (.CO(N1131), .S(N1130), .A(N376), .B(N384));
XNOR2X1 hap1_A_I1426 (.Y(N1132), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[15]));
OR2XL hap1_A_I1427 (.Y(N1133), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[15]));
ADDFX1 inst_blk01_cellmath__39_I358 (.CO(N1137), .S(N1136), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[1]), .CI(inst_blk01_cellmath__39_in0[6]));
ADDFXL inst_blk01_cellmath__39_I359 (.CO(N1139), .S(N1138), .A(N378), .B(N386), .CI(N368));
ADDFX1 inst_blk01_cellmath__39_I360 (.CO(N1141), .S(N1140), .A(inst_blk01_cellmath__39_in0[2]), .B(inst_blk01_cellmath__39_in0[16]), .CI(inst_blk01_cellmath__39_in0[4]));
ADDFXL inst_blk01_cellmath__39_I361 (.CO(N1143), .S(N1142), .A(N380), .B(inst_blk01_cellmath__39_in0[7]), .CI(N370));
ADDFX1 inst_blk01_cellmath__39_I362 (.CO(N1145), .S(N1144), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[17]), .CI(inst_blk01_cellmath__39_in0[5]));
ADDHX1 inst_blk01_cellmath__39_I363 (.CO(N1147), .S(N1146), .A(inst_blk01_cellmath__39_in0[8]), .B(N372));
ADDFX1 inst_blk01_cellmath__39_I364 (.CO(N1149), .S(N1148), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[18]), .CI(inst_blk01_cellmath__39_in0[6]));
ADDHX1 inst_blk01_cellmath__39_I365 (.CO(N1151), .S(N1150), .A(inst_blk01_cellmath__39_in0[9]), .B(N374));
ADDFX1 inst_blk01_cellmath__39_I366 (.CO(N1153), .S(N1152), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[19]), .CI(inst_blk01_cellmath__39_in0[7]));
ADDHX1 inst_blk01_cellmath__39_I367 (.CO(N1155), .S(N1154), .A(inst_blk01_cellmath__39_in0[10]), .B(N376));
ADDFX1 inst_blk01_cellmath__39_I368 (.CO(N1157), .S(N1156), .A(inst_blk01_cellmath__39_in0[6]), .B(inst_blk01_cellmath__39_in0[20]), .CI(inst_blk01_cellmath__39_in0[8]));
ADDHX1 inst_blk01_cellmath__39_I369 (.CO(N1159), .S(N1158), .A(inst_blk01_cellmath__39_in0[11]), .B(N378));
ADDFX1 inst_blk01_cellmath__39_I370 (.CO(N1161), .S(N1160), .A(inst_blk01_cellmath__39_in0[7]), .B(inst_blk01_cellmath__39_in0[21]), .CI(inst_blk01_cellmath__39_in0[9]));
XNOR2X1 hap1_A_I1428 (.Y(N1162), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[8]));
OR2XL hap1_A_I1429 (.Y(N1163), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[8]));
XNOR2X1 hap1_A_I1430 (.Y(N1166), .A(inst_blk01_cellmath__39_in0[5]), .B(N1482));
OR2XL hap1_A_I1431 (.Y(N1167), .A(inst_blk01_cellmath__39_in0[5]), .B(N1482));
ADDFX1 inst_blk01_cellmath__39_I373 (.CO(N1171), .S(N1170), .A(N354), .B(inst_blk01_cellmath__39_in0[6]), .CI(N3018));
ADDFX1 inst_blk01_cellmath__39_I374 (.CO(N1173), .S(N1172), .A(inst_blk01_cellmath__39_in0[0]), .B(inst_blk01_cellmath__39_in0[7]), .CI(N1484));
ADDHX1 inst_blk01_cellmath__39_I375 (.CO(N1175), .S(N1174), .A(N384), .B(N378));
ADDFX1 inst_blk01_cellmath__39_I376 (.CO(N1177), .S(N1176), .A(inst_blk01_cellmath__39_in0[1]), .B(inst_blk01_cellmath__39_in0[8]), .CI(N1381));
ADDFX1 inst_blk01_cellmath__39_I377 (.CO(N1179), .S(N1178), .A(N380), .B(N386), .CI(N374));
ADDFX1 inst_blk01_cellmath__39_I378 (.CO(N1181), .S(N1180), .A(N360), .B(N1482), .CI(N388));
ADDFX1 inst_blk01_cellmath__39_I379 (.CO(N1183), .S(N1182), .A(N376), .B(N3018), .CI(N1066));
ADDFX1 inst_blk01_cellmath__39_I380 (.CO(N1185), .S(N1184), .A(N390), .B(N362), .CI(N384));
ADDFX1 inst_blk01_cellmath__39_I381 (.CO(N1187), .S(N1186), .A(N1067), .B(N378), .CI(N1070));
ADDFX1 inst_blk01_cellmath__39_I382 (.CO(N1189), .S(N1188), .A(N386), .B(N1295), .CI(N3022));
ADDFX1 inst_blk01_cellmath__39_I383 (.CO(N1191), .S(N1190), .A(N1071), .B(N380), .CI(N1072));
ADDFX1 inst_blk01_cellmath__39_I384 (.CO(N1193), .S(N1192), .A(N388), .B(N366), .CI(N394));
ADDFX1 inst_blk01_cellmath__39_I385 (.CO(N1195), .S(N1194), .A(N1073), .B(N3018), .CI(N1074));
ADDFX1 inst_blk01_cellmath__39_I386 (.CO(N1197), .S(N1196), .A(N3024), .B(N368), .CI(N390));
ADDFX1 inst_blk01_cellmath__39_I387 (.CO(N1199), .S(N1198), .A(N1075), .B(N384), .CI(N1076));
ADDFX1 inst_blk01_cellmath__39_I388 (.CO(N1201), .S(N1200), .A(N386), .B(N370), .CI(N3022));
ADDFX1 inst_blk01_cellmath__39_I389 (.CO(N1203), .S(N1202), .A(N1082), .B(N1077), .CI(N1078));
ADDFX1 inst_blk01_cellmath__39_I390 (.CO(N1205), .S(N1204), .A(N388), .B(N394), .CI(N1079));
ADDFX1 inst_blk01_cellmath__39_I391 (.CO(N1207), .S(N1206), .A(N1084), .B(N1083), .CI(N1088));
ADDFHXL inst_blk01_cellmath__39_I392 (.CO(N1209), .S(N1208), .A(N1085), .B(N390), .CI(N1089));
ADDFX1 inst_blk01_cellmath__39_I393 (.CO(N1211), .S(N1210), .A(N1090), .B(N1096), .CI(N1094));
ADDFX1 inst_blk01_cellmath__39_I394 (.CO(N1213), .S(N1212), .A(N1097), .B(N1091), .CI(N1095));
ADDFX1 inst_blk01_cellmath__39_I395 (.CO(N1215), .S(N1214), .A(N1098), .B(N1104), .CI(N1102));
ADDFX1 inst_blk01_cellmath__39_I396 (.CO(N1217), .S(N1216), .A(N1099), .B(N394), .CI(N1105));
ADDFX1 inst_blk01_cellmath__39_I397 (.CO(N1219), .S(N1218), .A(N1106), .B(N1103), .CI(N1108));
ADDFXL inst_blk01_cellmath__39_I398 (.CO(N1221), .S(N1220), .A(N1107), .B(N3024), .CI(N1109));
ADDFX1 inst_blk01_cellmath__39_I399 (.CO(N1223), .S(N1222), .A(N1116), .B(N1110), .CI(N1114));
ADDFX1 inst_blk01_cellmath__39_I400 (.CO(N1225), .S(N1224), .A(N1117), .B(N1111), .CI(N1115));
ADDFX1 inst_blk01_cellmath__39_I401 (.CO(N1227), .S(N1226), .A(N1118), .B(N1124), .CI(N1122));
ADDFX1 inst_blk01_cellmath__39_I402 (.CO(N1229), .S(N1228), .A(N1125), .B(N1119), .CI(N1123));
ADDFX1 inst_blk01_cellmath__39_I403 (.CO(N1231), .S(N1230), .A(N1126), .B(N1130), .CI(N1128));
ADDFHXL inst_blk01_cellmath__39_I404 (.CO(N1233), .S(N1232), .A(N1127), .B(N1131), .CI(N1129));
ADDFX1 inst_blk01_cellmath__39_I405 (.CO(N1235), .S(N1234), .A(N1136), .B(N1132), .CI(N1138));
ADDFX1 inst_blk01_cellmath__39_I406 (.CO(N1237), .S(N1236), .A(N1133), .B(N388), .CI(N1137));
ADDFX1 inst_blk01_cellmath__39_I407 (.CO(N1239), .S(N1238), .A(N1140), .B(N1139), .CI(N1142));
ADDFX1 inst_blk01_cellmath__39_I408 (.CO(N1241), .S(N1240), .A(N390), .B(N3018), .CI(N1141));
ADDFX1 inst_blk01_cellmath__39_I409 (.CO(N1243), .S(N1242), .A(N1143), .B(N1146), .CI(N1144));
ADDFX1 inst_blk01_cellmath__39_I410 (.CO(N1245), .S(N1244), .A(N3022), .B(N384), .CI(N1147));
ADDFX1 inst_blk01_cellmath__39_I411 (.CO(N1247), .S(N1246), .A(N1150), .B(N1145), .CI(N1148));
ADDFX1 inst_blk01_cellmath__39_I412 (.CO(N1249), .S(N1248), .A(N394), .B(N386), .CI(N1151));
ADDFX1 inst_blk01_cellmath__39_I413 (.CO(N1251), .S(N1250), .A(N1154), .B(N1149), .CI(N1152));
ADDFX1 inst_blk01_cellmath__39_I414 (.CO(N1253), .S(N1252), .A(N3024), .B(N388), .CI(N1155));
ADDFX1 inst_blk01_cellmath__39_I415 (.CO(N1255), .S(N1254), .A(N1158), .B(N1153), .CI(N1156));
ADDFX1 inst_blk01_cellmath__39_I416 (.CO(N1257), .S(N1256), .A(N390), .B(inst_blk01_cellmath__39_in0[12]), .CI(N380));
ADDFX1 inst_blk01_cellmath__39_I417 (.CO(N1259), .S(N1258), .A(N1157), .B(N1159), .CI(N1160));
ADDFX1 inst_blk01_cellmath__39_I418 (.CO(N1261), .S(N1260), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[10]), .CI(N3018));
ADDFX1 inst_blk01_cellmath__39_I419 (.CO(N1263), .S(N1262), .A(N1161), .B(N3022), .CI(N1162));
ADDFX1 inst_blk01_cellmath__39_I420 (.CO(N1265), .S(N1264), .A(inst_blk01_cellmath__39_in0[11]), .B(inst_blk01_cellmath__39_in0[9]), .CI(inst_blk01_cellmath__39_in0[14]));
ADDFX1 inst_blk01_cellmath__39_I421 (.CO(N1267), .S(N1266), .A(N394), .B(N384), .CI(N1163));
ADDFX1 inst_blk01_cellmath__39_I422 (.CO(N1269), .S(N1268), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[10]), .CI(inst_blk01_cellmath__39_in0[15]));
ADDHX1 inst_blk01_cellmath__39_I423 (.CO(N1271), .S(N1270), .A(N386), .B(N3024));
ADDFX1 inst_blk01_cellmath__39_I424 (.CO(N1273), .S(N1272), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[11]), .CI(inst_blk01_cellmath__39_in0[16]));
XNOR2X1 hap1_A_I1432 (.Y(N1274), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[14]));
OR2XL hap1_A_I1433 (.Y(N1275), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[14]));
XNOR2X1 hap1_A_I1434 (.Y(N1278), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[15]));
OR2XL hap1_A_I1435 (.Y(N1279), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[15]));
XNOR2X1 hap1_A_I1436 (.Y(N1282), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[16]));
OR2XL hap1_A_I1437 (.Y(N1283), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[16]));
XNOR2X1 hap1_A_I1438 (.Y(N1286), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[17]));
OR2XL hap1_A_I1439 (.Y(N1287), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[17]));
INVXL inst_blk01_cellmath__39_I430 (.Y(N1294), .A(N1295));
ADDHX1 inst_blk01_cellmath__39_I431 (.CO(N1299), .S(N1298), .A(N366), .B(N360));
ADDHX1 inst_blk01_cellmath__39_I432 (.CO(N1301), .S(N1300), .A(N368), .B(N362));
ADDFX1 inst_blk01_cellmath__39_I433 (.CO(N1303), .S(N1302), .A(N370), .B(inst_blk01_cellmath__39_in0[0]), .CI(N1295));
ADDFX1 inst_blk01_cellmath__39_I434 (.CO(N1305), .S(N1304), .A(N372), .B(inst_blk01_cellmath__39_in0[1]), .CI(N366));
ADDFX1 inst_blk01_cellmath__39_I435 (.CO(N1307), .S(N1306), .A(N374), .B(inst_blk01_cellmath__39_in0[2]), .CI(N368));
ADDFX1 inst_blk01_cellmath__39_I436 (.CO(N1309), .S(N1308), .A(N376), .B(inst_blk01_cellmath__39_in0[3]), .CI(N370));
ADDFX1 inst_blk01_cellmath__39_I437 (.CO(N1311), .S(N1310), .A(N378), .B(inst_blk01_cellmath__39_in0[4]), .CI(N372));
ADDFX1 inst_blk01_cellmath__39_I438 (.CO(N1313), .S(N1312), .A(N374), .B(N380), .CI(N368));
ADDFX1 inst_blk01_cellmath__39_I439 (.CO(N1315), .S(N1314), .A(N376), .B(N370), .CI(N1167));
ADDFX1 inst_blk01_cellmath__39_I440 (.CO(N1317), .S(N1316), .A(N1174), .B(N372), .CI(N1171));
ADDFX1 inst_blk01_cellmath__39_I441 (.CO(N1319), .S(N1318), .A(N1173), .B(N1175), .CI(N1176));
ADDFX1 inst_blk01_cellmath__39_I442 (.CO(N1321), .S(N1320), .A(N1179), .B(N1177), .CI(N1180));
ADDFX1 inst_blk01_cellmath__39_I443 (.CO(N1323), .S(N1322), .A(N1184), .B(N1181), .CI(N1183));
ADDFX1 inst_blk01_cellmath__39_I444 (.CO(N1325), .S(N1324), .A(N1188), .B(N1185), .CI(N1187));
ADDFXL inst_blk01_cellmath__39_I445 (.CO(N1327), .S(N1326), .A(N1192), .B(N1189), .CI(N1191));
ADDFXL inst_blk01_cellmath__39_I446 (.CO(N1329), .S(N1328), .A(N1196), .B(N1193), .CI(N1195));
ADDFHXL inst_blk01_cellmath__39_I447 (.CO(N1331), .S(N1330), .A(N1200), .B(N1197), .CI(N1199));
ADDFX1 inst_blk01_cellmath__39_I448 (.CO(N1333), .S(N1332), .A(N1204), .B(N1201), .CI(N1203));
ADDFXL inst_blk01_cellmath__39_I449 (.CO(N1335), .S(N1334), .A(N1208), .B(N1205), .CI(N1207));
ADDFXL inst_blk01_cellmath__39_I450 (.CO(N1337), .S(N1336), .A(N1212), .B(N1209), .CI(N1211));
ADDFXL inst_blk01_cellmath__39_I451 (.CO(N1339), .S(N1338), .A(N1216), .B(N1213), .CI(N1215));
ADDFXL inst_blk01_cellmath__39_I452 (.CO(N1341), .S(N1340), .A(N1220), .B(N1217), .CI(N1219));
ADDFHXL inst_blk01_cellmath__39_I453 (.CO(N1343), .S(N1342), .A(N1223), .B(N1221), .CI(N1224));
ADDFHXL inst_blk01_cellmath__39_I454 (.CO(N1345), .S(N1344), .A(N1227), .B(N1225), .CI(N1228));
ADDFHXL inst_blk01_cellmath__39_I455 (.CO(N1347), .S(N1346), .A(N1232), .B(N1229), .CI(N1231));
ADDFXL inst_blk01_cellmath__39_I456 (.CO(N1349), .S(N1348), .A(N1236), .B(N1233), .CI(N1235));
ADDFHXL inst_blk01_cellmath__39_I457 (.CO(N1351), .S(N1350), .A(N1240), .B(N1237), .CI(N1239));
ADDFXL inst_blk01_cellmath__39_I458 (.CO(N1353), .S(N1352), .A(N1244), .B(N1241), .CI(N1243));
ADDFXL inst_blk01_cellmath__39_I459 (.CO(N1355), .S(N1354), .A(N1248), .B(N1245), .CI(N1247));
ADDFX1 inst_blk01_cellmath__39_I460 (.CO(N1357), .S(N1356), .A(N1252), .B(N1249), .CI(N1251));
ADDFXL inst_blk01_cellmath__39_I461 (.CO(N1359), .S(N1358), .A(N1253), .B(N1256), .CI(N1255));
ADDFX1 inst_blk01_cellmath__39_I462 (.CO(N1361), .S(N1360), .A(N1260), .B(N1257), .CI(N1259));
ADDFX1 inst_blk01_cellmath__39_I463 (.CO(N1363), .S(N1362), .A(N1264), .B(N1261), .CI(N1263));
ADDFX1 inst_blk01_cellmath__39_I464 (.CO(N1365), .S(N1364), .A(N1270), .B(N1265), .CI(N1268));
ADDFX1 inst_blk01_cellmath__39_I465 (.CO(N1367), .S(N1366), .A(N1271), .B(N388), .CI(N1269));
ADDFX1 inst_blk01_cellmath__39_I466 (.CO(N1369), .S(N1368), .A(N390), .B(inst_blk01_cellmath__39_in0[17]), .CI(N1273));
ADDFX1 inst_blk01_cellmath__39_I467 (.CO(N1371), .S(N1370), .A(N3022), .B(inst_blk01_cellmath__39_in0[18]), .CI(N1275));
ADDFX1 inst_blk01_cellmath__39_I468 (.CO(N1373), .S(N1372), .A(N394), .B(inst_blk01_cellmath__39_in0[19]), .CI(N1279));
ADDFX1 inst_blk01_cellmath__39_I469 (.CO(N1375), .S(N1374), .A(N3024), .B(inst_blk01_cellmath__39_in0[20]), .CI(N1283));
ADDFX1 inst_blk01_cellmath__39_I470 (.CO(N1377), .S(N1376), .A(inst_blk01_cellmath__39_in0[21]), .B(inst_blk01_cellmath__39_in0[18]), .CI(N384));
ADDFX1 inst_blk01_cellmath__39_I471 (.CO(N1379), .S(N1378), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[17]), .CI(inst_blk01_cellmath__39_in0[22]));
INVXL inst_blk01_cellmath__39_I472 (.Y(N1380), .A(N1381));
ADDHX1 inst_blk01_cellmath__39_I473 (.CO(N1385), .S(N1384), .A(N360), .B(N354));
ADDHX1 inst_blk01_cellmath__39_I474 (.CO(N1387), .S(N1386), .A(N362), .B(N1484));
ADDFX1 inst_blk01_cellmath__39_I475 (.CO(N1389), .S(N1388), .A(N1482), .B(N1381), .CI(N1294));
ADDFX1 inst_blk01_cellmath__39_I476 (.CO(N1391), .S(N1390), .A(N1295), .B(N354), .CI(N1298));
ADDFX1 inst_blk01_cellmath__39_I477 (.CO(N1393), .S(N1392), .A(N1299), .B(N1484), .CI(N1300));
ADDFX1 inst_blk01_cellmath__39_I478 (.CO(N1395), .S(N1394), .A(N1301), .B(N1381), .CI(N1302));
ADDFX1 inst_blk01_cellmath__39_I479 (.CO(N1397), .S(N1396), .A(N1303), .B(N360), .CI(N1304));
ADDFX1 inst_blk01_cellmath__39_I480 (.CO(N1399), .S(N1398), .A(N1305), .B(N362), .CI(N1306));
ADDFX1 inst_blk01_cellmath__39_I481 (.CO(N1401), .S(N1400), .A(N1307), .B(N1295), .CI(N1308));
ADDFX1 inst_blk01_cellmath__39_I482 (.CO(N1403), .S(N1402), .A(N1309), .B(N366), .CI(N1310));
ADDFX1 inst_blk01_cellmath__39_I483 (.CO(N1405), .S(N1404), .A(N1166), .B(N1311), .CI(N1312));
ADDFX1 inst_blk01_cellmath__39_I484 (.CO(N1407), .S(N1406), .A(N1170), .B(N1313), .CI(N1314));
ADDFX1 inst_blk01_cellmath__39_I485 (.CO(N1409), .S(N1408), .A(N1315), .B(N1172), .CI(N1316));
ADDFX1 inst_blk01_cellmath__39_I486 (.CO(N1411), .S(N1410), .A(N1317), .B(N1178), .CI(N1318));
ADDFX1 inst_blk01_cellmath__39_I487 (.CO(N1413), .S(N1412), .A(N1182), .B(N1319), .CI(N1320));
ADDFX1 inst_blk01_cellmath__39_I488 (.CO(N1415), .S(N1414), .A(N1186), .B(N1321), .CI(N1322));
ADDFHXL inst_blk01_cellmath__39_I489 (.CO(N1417), .S(N1416), .A(N1323), .B(N1190), .CI(N1324));
ADDFHXL inst_blk01_cellmath__39_I490 (.CO(N1419), .S(N1418), .A(N1325), .B(N1194), .CI(N1326));
ADDFHXL inst_blk01_cellmath__39_I491 (.CO(N1421), .S(N1420), .A(N1327), .B(N1198), .CI(N1328));
ADDFHXL inst_blk01_cellmath__39_I492 (.CO(N1423), .S(N1422), .A(N1329), .B(N1202), .CI(N1330));
ADDFX1 inst_blk01_cellmath__39_I493 (.CO(N1425), .S(N1424), .A(N1331), .B(N1206), .CI(N1332));
ADDFHXL inst_blk01_cellmath__39_I494 (.CO(N1427), .S(N1426), .A(N1333), .B(N1210), .CI(N1334));
ADDFHXL inst_blk01_cellmath__39_I495 (.CO(N1429), .S(N1428), .A(N1335), .B(N1214), .CI(N1336));
ADDFHXL inst_blk01_cellmath__39_I496 (.CO(N1431), .S(N1430), .A(N1337), .B(N1218), .CI(N1338));
ADDFHX1 inst_blk01_cellmath__39_I497 (.CO(N1433), .S(N1432), .A(N1339), .B(N1222), .CI(N1340));
ADDFHX1 inst_blk01_cellmath__39_I498 (.CO(N1435), .S(N1434), .A(N1341), .B(N1226), .CI(N1342));
ADDFHXL inst_blk01_cellmath__39_I499 (.CO(N1437), .S(N1436), .A(N1343), .B(N1230), .CI(N1344));
ADDFHX1 inst_blk01_cellmath__39_I500 (.CO(N1439), .S(N1438), .A(N1345), .B(N1234), .CI(N1346));
ADDFHXL inst_blk01_cellmath__39_I501 (.CO(N1441), .S(N1440), .A(N1347), .B(N1238), .CI(N1348));
ADDFHX1 inst_blk01_cellmath__39_I502 (.CO(N1443), .S(N1442), .A(N1349), .B(N1242), .CI(N1350));
ADDFX1 inst_blk01_cellmath__39_I503 (.CO(N1445), .S(N1444), .A(N1351), .B(N1246), .CI(N1352));
ADDFX1 inst_blk01_cellmath__39_I504 (.CO(N1447), .S(N1446), .A(N1353), .B(N1250), .CI(N1354));
ADDFHX1 inst_blk01_cellmath__39_I505 (.CO(N1449), .S(N1448), .A(N1355), .B(N1254), .CI(N1356));
ADDFHXL inst_blk01_cellmath__39_I506 (.CO(N1451), .S(N1450), .A(N1357), .B(N1258), .CI(N1358));
ADDFXL inst_blk01_cellmath__39_I507 (.CO(N1453), .S(N1452), .A(N1359), .B(N1262), .CI(N1360));
ADDFX1 inst_blk01_cellmath__39_I508 (.CO(N1455), .S(N1454), .A(N1361), .B(N1266), .CI(N1362));
ADDFX1 inst_blk01_cellmath__39_I509 (.CO(N1457), .S(N1456), .A(N1364), .B(N1267), .CI(N1363));
ADDFX1 inst_blk01_cellmath__39_I510 (.CO(N1459), .S(N1458), .A(N1366), .B(N1272), .CI(N1365));
ADDFX1 inst_blk01_cellmath__39_I511 (.CO(N1461), .S(N1460), .A(N1367), .B(N1274), .CI(N1368));
ADDFX1 inst_blk01_cellmath__39_I512 (.CO(N1463), .S(N1462), .A(N1369), .B(N1278), .CI(N1370));
ADDFX1 inst_blk01_cellmath__39_I513 (.CO(N1465), .S(N1464), .A(N1371), .B(N1282), .CI(N1372));
ADDFX1 inst_blk01_cellmath__39_I514 (.CO(N1467), .S(N1466), .A(N1373), .B(N1286), .CI(N1374));
ADDFX1 inst_blk01_cellmath__39_I515 (.CO(N1469), .S(N1468), .A(N1376), .B(N1287), .CI(N1375));
ADDFX1 inst_blk01_cellmath__39_I516 (.CO(N1471), .S(N1470), .A(N1377), .B(inst_blk01_cellmath__39_in0[16]), .CI(N1378));
ADDFX1 inst_blk01_cellmath__39_I517 (.CO(N1473), .S(N1472), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[18]), .CI(N1379));
ADDHX1 inst_blk01_cellmath__39_I518 (.CO(N1475), .S(N1474), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[21]));
ADDHX1 inst_blk01_cellmath__39_I519 (.CO(N1477), .S(N1476), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[22]));
INVXL inst_blk01_cellmath__39_I1588 (.Y(inst_blk01_cellmath__39_out0[1]), .A(N1482));
INVXL inst_blk01_cellmath__39_I522 (.Y(N1483), .A(N354));
NOR2XL inst_blk01_cellmath__39_I524 (.Y(N1485), .A(N1482), .B(N1380));
NAND2XL inst_blk01_cellmath__39_I525 (.Y(N1486), .A(N1482), .B(N1380));
NOR2XL inst_blk01_cellmath__39_I526 (.Y(N1487), .A(N1381), .B(N1384));
NAND2XL inst_blk01_cellmath__39_I527 (.Y(N1488), .A(N1381), .B(N1384));
NOR2XL inst_blk01_cellmath__39_I528 (.Y(N1489), .A(N1385), .B(N1386));
NAND2XL inst_blk01_cellmath__39_I529 (.Y(N1490), .A(N1385), .B(N1386));
NOR2XL inst_blk01_cellmath__39_I530 (.Y(N1491), .A(N1387), .B(N1388));
NAND2XL inst_blk01_cellmath__39_I531 (.Y(N1492), .A(N1387), .B(N1388));
NOR2XL inst_blk01_cellmath__39_I532 (.Y(N1493), .A(N1389), .B(N1390));
NAND2XL inst_blk01_cellmath__39_I533 (.Y(N1494), .A(N1389), .B(N1390));
NOR2XL inst_blk01_cellmath__39_I534 (.Y(N1495), .A(N1391), .B(N1392));
NAND2XL inst_blk01_cellmath__39_I535 (.Y(N1496), .A(N1391), .B(N1392));
NOR2XL inst_blk01_cellmath__39_I536 (.Y(N1497), .A(N1393), .B(N1394));
NAND2XL inst_blk01_cellmath__39_I537 (.Y(N1498), .A(N1393), .B(N1394));
NOR2XL inst_blk01_cellmath__39_I538 (.Y(N1499), .A(N1395), .B(N1396));
NAND2XL inst_blk01_cellmath__39_I539 (.Y(N1500), .A(N1395), .B(N1396));
NOR2XL inst_blk01_cellmath__39_I540 (.Y(N1501), .A(N1397), .B(N1398));
NAND2XL inst_blk01_cellmath__39_I541 (.Y(N1502), .A(N1397), .B(N1398));
NOR2XL inst_blk01_cellmath__39_I542 (.Y(N1503), .A(N1399), .B(N1400));
NAND2X1 inst_blk01_cellmath__39_I543 (.Y(N1504), .A(N1399), .B(N1400));
NOR2XL inst_blk01_cellmath__39_I544 (.Y(N1505), .A(N1401), .B(N1402));
NAND2XL inst_blk01_cellmath__39_I545 (.Y(N1506), .A(N1401), .B(N1402));
NOR2XL inst_blk01_cellmath__39_I546 (.Y(N1507), .A(N1403), .B(N1404));
NAND2XL inst_blk01_cellmath__39_I547 (.Y(N1508), .A(N1403), .B(N1404));
NOR2XL inst_blk01_cellmath__39_I550 (.Y(N1511), .A(N1483), .B(inst_blk01_cellmath__39_out0[1]));
NAND2XL inst_blk01_cellmath__39_I558 (.Y(N1521), .A(N1484), .B(N1511));
AOI21XL inst_blk01_cellmath__39_I566 (.Y(N1531), .A0(N1486), .A1(N1521), .B0(N1485));
AOI21XL inst_blk01_cellmath__39_I570 (.Y(N1535), .A0(N1490), .A1(N1487), .B0(N1489));
NAND2XL inst_blk01_cellmath__39_I571 (.Y(N1536), .A(N1490), .B(N1488));
OAI21XL inst_blk01_cellmath__39_I582 (.Y(N1547), .A0(N1536), .A1(N1531), .B0(N1535));
AOI21XL inst_blk01_cellmath__39_I596 (.Y(N1561), .A0(N1492), .A1(N1547), .B0(N1491));
AOI21XL inst_blk01_cellmath__39_I600 (.Y(N1565), .A0(N1496), .A1(N1493), .B0(N1495));
NAND2XL inst_blk01_cellmath__39_I601 (.Y(N1566), .A(N1496), .B(N1494));
OAI21X1 inst_blk01_cellmath__39_I618 (.Y(N1583), .A0(N1566), .A1(N1561), .B0(N1565));
AO21XL inst_blk01_cellmath__39_I1916 (.Y(N3069), .A0(N1500), .A1(N1497), .B0(N1499));
AND2XL inst_blk01_cellmath__39_I1843 (.Y(N3070), .A(N1500), .B(N1498));
NOR2BX1 andori2bb1_A_I3341 (.Y(N3282), .AN(N1488), .B(N1531));
NOR2XL andori2bb1_A_I1970 (.Y(N3075), .A(N3282), .B(N1487));
NOR2BX1 andori2bb1_A_I3342 (.Y(N3289), .AN(N1494), .B(N1561));
NOR2XL andori2bb1_A_I1972 (.Y(N3078), .A(N3289), .B(N1493));
AOI21XL inst_blk01_cellmath__39_I646 (.Y(N1611), .A0(N1498), .A1(N1583), .B0(N1497));
AOI21X1 inst_blk01_cellmath__39_I648 (.Y(N1613), .A0(N3070), .A1(N1583), .B0(N3069));
AOI21XL inst_blk01_cellmath__39_I652 (.Y(N1617), .A0(N1504), .A1(N1501), .B0(N1503));
NAND2XL inst_blk01_cellmath__39_I653 (.Y(N1618), .A(N1504), .B(N1502));
INVXL inst_blk01_cellmath__39_I1640 (.Y(N3087), .A(N1506));
AOI21XL inst_blk01_cellmath__39_I656 (.Y(N1621), .A0(N1508), .A1(N1505), .B0(N1507));
NAND2XL inst_blk01_cellmath__39_I657 (.Y(N1622), .A(N1508), .B(N1506));
INVXL inst_blk01_cellmath__39_I1645 (.Y(N3092), .A(N1501));
INVXL inst_blk01_cellmath__39_I1646 (.Y(N3093), .A(N1502));
NOR2XL andori2bb1_A_I1973 (.Y(N3296), .A(N3087), .B(N1617));
NOR2XL andori2bb1_A_I1974 (.Y(N3096), .A(N3296), .B(N1505));
OA21X1 inst_blk01_cellmath__39_I1921 (.Y(N3098), .A0(N1622), .A1(N1617), .B0(N1621));
OR2XL inst_blk01_cellmath__39_I1850 (.Y(N3099), .A(N1622), .B(N1618));
OAI21XL inst_blk01_cellmath__39_I696 (.Y(N1661), .A0(N3093), .A1(N1613), .B0(N3092));
OAI21XL inst_blk01_cellmath__39_I698 (.Y(N1663), .A0(N1618), .A1(N1613), .B0(N1617));
OAI31X1 inst_blk01_cellmath__39_I1852 (.Y(N1665), .A0(N3087), .A1(N1618), .A2(N1613), .B0(N3096));
OAI21X1 inst_blk01_cellmath__39_I702 (.Y(N1734), .A0(N3099), .A1(N1613), .B0(N3098));
NAND2BXL inst_blk01_cellmath__39_I715 (.Y(N1684), .AN(N1485), .B(N1486));
NAND2BXL inst_blk01_cellmath__39_I718 (.Y(N1687), .AN(N1487), .B(N1488));
NAND2BXL inst_blk01_cellmath__39_I721 (.Y(N1690), .AN(N1489), .B(N1490));
NAND2BXL inst_blk01_cellmath__39_I724 (.Y(N1693), .AN(N1491), .B(N1492));
NAND2BXL inst_blk01_cellmath__39_I727 (.Y(N1696), .AN(N1493), .B(N1494));
NAND2BXL inst_blk01_cellmath__39_I730 (.Y(N1699), .AN(N1495), .B(N1496));
NAND2BXL inst_blk01_cellmath__39_I733 (.Y(N1702), .AN(N1497), .B(N1498));
NAND2BXL inst_blk01_cellmath__39_I736 (.Y(N1705), .AN(N1499), .B(N1500));
NAND2BXL inst_blk01_cellmath__39_I739 (.Y(N1708), .AN(N1501), .B(N1502));
NAND2BXL inst_blk01_cellmath__39_I742 (.Y(N1711), .AN(N1503), .B(N1504));
NAND2BXL inst_blk01_cellmath__39_I745 (.Y(N1714), .AN(N1505), .B(N1506));
NAND2BXL inst_blk01_cellmath__39_I748 (.Y(N1717), .AN(N1507), .B(N1508));
XOR2XL inst_blk01_cellmath__39_I3345 (.Y(inst_blk01_cellmath__39_out0[2]), .A(inst_blk01_cellmath__39_out0[1]), .B(N1483));
XOR2XL inst_blk01_cellmath__39_I1855 (.Y(inst_blk01_cellmath__39_out0[3]), .A(N1511), .B(N1484));
XOR2XL inst_blk01_cellmath__39_I1856 (.Y(inst_blk01_cellmath__39_out0[4]), .A(N1521), .B(N1684));
XNOR2X1 inst_blk01_cellmath__39_I753 (.Y(inst_blk01_cellmath__39_out0[5]), .A(N1531), .B(N1687));
XNOR2X1 inst_blk01_cellmath__39_I754 (.Y(inst_blk01_cellmath__39_out0[6]), .A(N3075), .B(N1690));
XOR2XL inst_blk01_cellmath__39_I1857 (.Y(inst_blk01_cellmath__39_out0[7]), .A(N1547), .B(N1693));
XNOR2X1 inst_blk01_cellmath__39_I756 (.Y(inst_blk01_cellmath__39_out0[8]), .A(N1561), .B(N1696));
XNOR2X1 inst_blk01_cellmath__39_I757 (.Y(inst_blk01_cellmath__39_out0[9]), .A(N3078), .B(N1699));
XOR2XL inst_blk01_cellmath__39_I1858 (.Y(inst_blk01_cellmath__39_out0[10]), .A(N1583), .B(N1702));
XNOR2X1 inst_blk01_cellmath__39_I759 (.Y(inst_blk01_cellmath__39_out0[11]), .A(N1611), .B(N1705));
XNOR2X1 inst_blk01_cellmath__39_I760 (.Y(inst_blk01_cellmath__39_out0[12]), .A(N1613), .B(N1708));
XOR2XL inst_blk01_cellmath__39_I761 (.Y(inst_blk01_cellmath__39_out0[13]), .A(N1661), .B(N1711));
XOR2XL inst_blk01_cellmath__39_I762 (.Y(inst_blk01_cellmath__39_out0[14]), .A(N1663), .B(N1714));
XOR2XL inst_blk01_cellmath__39_I763 (.Y(inst_blk01_cellmath__39_out0[15]), .A(N1665), .B(N1717));
NOR2XL inst_blk01_cellmath__39_I766 (.Y(N1736), .A(N1405), .B(N1406));
NAND2XL inst_blk01_cellmath__39_I767 (.Y(N1737), .A(N1405), .B(N1406));
NOR2XL inst_blk01_cellmath__39_I768 (.Y(N1738), .A(N1407), .B(N1408));
NAND2XL inst_blk01_cellmath__39_I769 (.Y(N1739), .A(N1407), .B(N1408));
NOR2XL inst_blk01_cellmath__39_I770 (.Y(N1740), .A(N1409), .B(N1410));
NAND2XL inst_blk01_cellmath__39_I771 (.Y(N1741), .A(N1409), .B(N1410));
NOR2XL inst_blk01_cellmath__39_I772 (.Y(N1742), .A(N1411), .B(N1412));
NAND2XL inst_blk01_cellmath__39_I773 (.Y(N1743), .A(N1411), .B(N1412));
NOR2XL inst_blk01_cellmath__39_I774 (.Y(N1744), .A(N1413), .B(N1414));
NAND2X1 inst_blk01_cellmath__39_I775 (.Y(N1745), .A(N1413), .B(N1414));
NOR2X2 inst_blk01_cellmath__39_I776 (.Y(N1746), .A(N1415), .B(N1416));
NAND2X2 inst_blk01_cellmath__39_I777 (.Y(N1747), .A(N1415), .B(N1416));
NOR2X1 inst_blk01_cellmath__39_I778 (.Y(N1748), .A(N1417), .B(N1418));
NAND2X4 inst_blk01_cellmath__39_I779 (.Y(N1749), .A(N1417), .B(N1418));
NOR2X4 inst_blk01_cellmath__39_I780 (.Y(N1750), .A(N1419), .B(N1420));
NAND2X2 inst_blk01_cellmath__39_I781 (.Y(N1751), .A(N1419), .B(N1420));
NOR2X1 inst_blk01_cellmath__39_I782 (.Y(N1752), .A(N1421), .B(N1422));
NAND2X4 inst_blk01_cellmath__39_I783 (.Y(N1753), .A(N1421), .B(N1422));
NOR2X2 inst_blk01_cellmath__39_I784 (.Y(N1754), .A(N1423), .B(N1424));
NAND2X2 inst_blk01_cellmath__39_I785 (.Y(N1755), .A(N1423), .B(N1424));
NOR2X1 inst_blk01_cellmath__39_I1859 (.Y(N1756), .A(N1426), .B(N1425));
NAND2X4 inst_blk01_cellmath__39_I787 (.Y(N1757), .A(N1425), .B(N1426));
NOR2X2 inst_blk01_cellmath__39_I788 (.Y(N1758), .A(N1427), .B(N1428));
NAND2X2 inst_blk01_cellmath__39_I789 (.Y(N1759), .A(N1427), .B(N1428));
NOR2X1 inst_blk01_cellmath__39_I790 (.Y(N1760), .A(N1429), .B(N1430));
NAND2X4 inst_blk01_cellmath__39_I791 (.Y(N1761), .A(N1429), .B(N1430));
NOR2X2 inst_blk01_cellmath__39_I792 (.Y(N1762), .A(N1431), .B(N1432));
NAND2X4 inst_blk01_cellmath__39_I793 (.Y(N1763), .A(N1431), .B(N1432));
NOR2X1 inst_blk01_cellmath__39_I794 (.Y(N1764), .A(N1433), .B(N1434));
NAND2X4 inst_blk01_cellmath__39_I795 (.Y(N1765), .A(N1433), .B(N1434));
NOR2X2 inst_blk01_cellmath__39_I796 (.Y(N1766), .A(N1435), .B(N1436));
NAND2X1 inst_blk01_cellmath__39_I797 (.Y(N1767), .A(N1435), .B(N1436));
NOR2X1 inst_blk01_cellmath__39_I1926 (.Y(N1768), .A(N1438), .B(N1437));
NAND2X4 inst_blk01_cellmath__39_I799 (.Y(N1769), .A(N1437), .B(N1438));
NOR2X2 inst_blk01_cellmath__39_I800 (.Y(N1770), .A(N1439), .B(N1440));
NAND2X2 inst_blk01_cellmath__39_I801 (.Y(N1771), .A(N1439), .B(N1440));
NOR2X1 inst_blk01_cellmath__39_I802 (.Y(N1772), .A(N1441), .B(N1442));
NAND2X4 inst_blk01_cellmath__39_I803 (.Y(N1773), .A(N1441), .B(N1442));
NOR2X2 inst_blk01_cellmath__39_I804 (.Y(N1774), .A(N1443), .B(N1444));
NAND2X1 inst_blk01_cellmath__39_I805 (.Y(N1775), .A(N1443), .B(N1444));
NOR2X1 inst_blk01_cellmath__39_I806 (.Y(N1776), .A(N1445), .B(N1446));
NAND2X4 inst_blk01_cellmath__39_I807 (.Y(N1777), .A(N1445), .B(N1446));
NOR2X2 inst_blk01_cellmath__39_I808 (.Y(N1778), .A(N1447), .B(N1448));
NAND2X4 inst_blk01_cellmath__39_I809 (.Y(N1779), .A(N1447), .B(N1448));
NOR2XL inst_blk01_cellmath__39_I810 (.Y(N1780), .A(N1449), .B(N1450));
NAND2X4 inst_blk01_cellmath__39_I811 (.Y(N1781), .A(N1449), .B(N1450));
NOR2X2 inst_blk01_cellmath__39_I812 (.Y(N1782), .A(N1451), .B(N1452));
NAND2X1 inst_blk01_cellmath__39_I813 (.Y(N1783), .A(N1451), .B(N1452));
NOR2XL inst_blk01_cellmath__39_I814 (.Y(N1784), .A(N1453), .B(N1454));
NAND2X2 inst_blk01_cellmath__39_I815 (.Y(N1785), .A(N1453), .B(N1454));
NOR2XL inst_blk01_cellmath__39_I816 (.Y(N1786), .A(N1455), .B(N1456));
NAND2XL inst_blk01_cellmath__39_I817 (.Y(N1787), .A(N1455), .B(N1456));
NOR2XL inst_blk01_cellmath__39_I818 (.Y(N1788), .A(N1458), .B(N1457));
NAND2XL inst_blk01_cellmath__39_I819 (.Y(N1789), .A(N1458), .B(N1457));
NOR2XL inst_blk01_cellmath__39_I820 (.Y(N1790), .A(N1459), .B(N1460));
NAND2XL inst_blk01_cellmath__39_I821 (.Y(N1791), .A(N1459), .B(N1460));
NOR2XL inst_blk01_cellmath__39_I822 (.Y(N1792), .A(N1461), .B(N1462));
NAND2XL inst_blk01_cellmath__39_I823 (.Y(N1793), .A(N1461), .B(N1462));
NOR2XL inst_blk01_cellmath__39_I824 (.Y(N1794), .A(N1463), .B(N1464));
NAND2XL inst_blk01_cellmath__39_I825 (.Y(N1795), .A(N1463), .B(N1464));
NOR2XL inst_blk01_cellmath__39_I826 (.Y(N1796), .A(N1465), .B(N1466));
NAND2XL inst_blk01_cellmath__39_I827 (.Y(N1797), .A(N1465), .B(N1466));
NOR2XL inst_blk01_cellmath__39_I828 (.Y(N1798), .A(N1467), .B(N1468));
NAND2XL inst_blk01_cellmath__39_I829 (.Y(N1799), .A(N1467), .B(N1468));
NOR2XL inst_blk01_cellmath__39_I830 (.Y(N1800), .A(N1469), .B(N1470));
NAND2XL inst_blk01_cellmath__39_I831 (.Y(N1801), .A(N1469), .B(N1470));
NOR2XL inst_blk01_cellmath__39_I832 (.Y(N1802), .A(N1472), .B(N1471));
NAND2XL inst_blk01_cellmath__39_I833 (.Y(N1803), .A(N1472), .B(N1471));
NOR2XL inst_blk01_cellmath__39_I834 (.Y(N1804), .A(N1474), .B(N1473));
NAND2XL inst_blk01_cellmath__39_I835 (.Y(N1805), .A(N1474), .B(N1473));
NOR2XL inst_blk01_cellmath__39_I836 (.Y(N1806), .A(N1475), .B(N1476));
NAND2XL inst_blk01_cellmath__39_I837 (.Y(N1807), .A(N1475), .B(N1476));
NOR2XL inst_blk01_cellmath__39_I838 (.Y(N1808), .A(N394), .B(N1477));
NAND2XL inst_blk01_cellmath__39_I839 (.Y(N1809), .A(N394), .B(N1477));
NOR2XL inst_blk01_cellmath__39_I840 (.Y(N1810), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[21]));
NAND2XL inst_blk01_cellmath__39_I841 (.Y(N1811), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[21]));
AOI21X2 inst_blk01_cellmath__39_I844 (.Y(N1814), .A0(N1737), .A1(N1734), .B0(N1736));
AOI21XL inst_blk01_cellmath__39_I848 (.Y(N1818), .A0(N1741), .A1(N1738), .B0(N1740));
NAND2XL inst_blk01_cellmath__39_I849 (.Y(N1819), .A(N1741), .B(N1739));
OAI21X2 inst_blk01_cellmath__39_I856 (.Y(N1826), .A0(N1819), .A1(N1814), .B0(N1818));
AOI21X2 inst_blk01_cellmath__39_I860 (.Y(N1830), .A0(N1745), .A1(N1742), .B0(N1744));
NAND2X1 inst_blk01_cellmath__39_I861 (.Y(N1831), .A(N1745), .B(N1743));
INVXL inst_blk01_cellmath__39_I1666 (.Y(N3113), .A(N1747));
AOI21X4 inst_blk01_cellmath__39_I864 (.Y(N1834), .A0(N1749), .A1(N1746), .B0(N1748));
NAND2X4 inst_blk01_cellmath__39_I865 (.Y(N1835), .A(N1749), .B(N1747));
OAI21X4 inst_blk01_cellmath__39_I872 (.Y(N1842), .A0(N1835), .A1(N1830), .B0(N1834));
NOR2X4 inst_blk01_cellmath__39_I873 (.Y(N1843), .A(N1835), .B(N1831));
AOI21X4 inst_blk01_cellmath__39_I876 (.Y(N1846), .A0(N1753), .A1(N1750), .B0(N1752));
NAND2X2 inst_blk01_cellmath__39_I877 (.Y(N1847), .A(N1753), .B(N1751));
INVXL inst_blk01_cellmath__39_I1674 (.Y(N3121), .A(N1755));
AOI21X4 inst_blk01_cellmath__39_I880 (.Y(N1850), .A0(N1757), .A1(N1754), .B0(N1756));
NAND2X4 inst_blk01_cellmath__39_I881 (.Y(N1851), .A(N1757), .B(N1755));
OAI21X4 inst_blk01_cellmath__39_I888 (.Y(N1858), .A0(N1851), .A1(N1846), .B0(N1850));
NOR2X4 inst_blk01_cellmath__39_I889 (.Y(N1859), .A(N1851), .B(N1847));
AOI21X4 inst_blk01_cellmath__39_I892 (.Y(N1862), .A0(N1761), .A1(N1758), .B0(N1760));
NAND2X4 inst_blk01_cellmath__39_I893 (.Y(N1863), .A(N1761), .B(N1759));
INVXL inst_blk01_cellmath__39_I1684 (.Y(N3131), .A(N1763));
AOI21X4 inst_blk01_cellmath__39_I896 (.Y(N1866), .A0(N1765), .A1(N1762), .B0(N1764));
NAND2X4 inst_blk01_cellmath__39_I897 (.Y(N1867), .A(N1765), .B(N1763));
OAI21X4 inst_blk01_cellmath__39_I904 (.Y(N1874), .A0(N1867), .A1(N1862), .B0(N1866));
NOR2X6 inst_blk01_cellmath__39_I905 (.Y(N1875), .A(N1867), .B(N1863));
AOI21X4 inst_blk01_cellmath__39_I908 (.Y(N1878), .A0(N1769), .A1(N1766), .B0(N1768));
NAND2X2 inst_blk01_cellmath__39_I909 (.Y(N1879), .A(N1769), .B(N1767));
INVXL inst_blk01_cellmath__39_I1694 (.Y(N3141), .A(N1771));
AOI21X4 inst_blk01_cellmath__39_I912 (.Y(N1882), .A0(N1773), .A1(N1770), .B0(N1772));
NAND2X4 inst_blk01_cellmath__39_I913 (.Y(N1883), .A(N1773), .B(N1771));
OAI21X4 inst_blk01_cellmath__39_I920 (.Y(N1890), .A0(N1883), .A1(N1878), .B0(N1882));
NOR2X6 inst_blk01_cellmath__39_I921 (.Y(N1891), .A(N1883), .B(N1879));
AOI21X4 inst_blk01_cellmath__39_I924 (.Y(N1894), .A0(N1777), .A1(N1774), .B0(N1776));
NAND2X2 inst_blk01_cellmath__39_I925 (.Y(N1895), .A(N1777), .B(N1775));
INVXL inst_blk01_cellmath__39_I1704 (.Y(N3151), .A(N1779));
AOI21X2 inst_blk01_cellmath__39_I928 (.Y(N1898), .A0(N1781), .A1(N1778), .B0(N1780));
NAND2X6 inst_blk01_cellmath__39_I929 (.Y(N1899), .A(N1781), .B(N1779));
OAI21X4 inst_blk01_cellmath__39_I936 (.Y(N1906), .A0(N1899), .A1(N1894), .B0(N1898));
NOR2X4 inst_blk01_cellmath__39_I937 (.Y(N1907), .A(N1899), .B(N1895));
AOI21X2 inst_blk01_cellmath__39_I940 (.Y(N1910), .A0(N1785), .A1(N1782), .B0(N1784));
NAND2X2 inst_blk01_cellmath__39_I941 (.Y(N1911), .A(N1785), .B(N1783));
INVXL inst_blk01_cellmath__39_I1712 (.Y(N3159), .A(N1787));
AOI21XL inst_blk01_cellmath__39_I944 (.Y(N1914), .A0(N1789), .A1(N1786), .B0(N1788));
NAND2X1 inst_blk01_cellmath__39_I945 (.Y(N1915), .A(N1789), .B(N1787));
OAI21X2 inst_blk01_cellmath__39_I952 (.Y(N1922), .A0(N1915), .A1(N1910), .B0(N1914));
NOR2X4 inst_blk01_cellmath__39_I953 (.Y(N1923), .A(N1915), .B(N1911));
AOI21X1 inst_blk01_cellmath__39_I956 (.Y(N1926), .A0(N1793), .A1(N1790), .B0(N1792));
NAND2XL inst_blk01_cellmath__39_I957 (.Y(N1927), .A(N1793), .B(N1791));
INVXL inst_blk01_cellmath__39_I1720 (.Y(N3167), .A(N1795));
AOI21XL inst_blk01_cellmath__39_I960 (.Y(N1930), .A0(N1797), .A1(N1794), .B0(N1796));
NAND2XL inst_blk01_cellmath__39_I961 (.Y(N1931), .A(N1797), .B(N1795));
OAI21XL inst_blk01_cellmath__39_I968 (.Y(N1938), .A0(N1931), .A1(N1926), .B0(N1930));
NOR2XL inst_blk01_cellmath__39_I969 (.Y(N1939), .A(N1931), .B(N1927));
AOI21XL inst_blk01_cellmath__39_I972 (.Y(N1942), .A0(N1801), .A1(N1798), .B0(N1800));
NAND2XL inst_blk01_cellmath__39_I973 (.Y(N1943), .A(N1801), .B(N1799));
INVXL inst_blk01_cellmath__39_I1727 (.Y(N3174), .A(N1802));
INVXL inst_blk01_cellmath__39_I1728 (.Y(N3175), .A(N1803));
AOI21XL inst_blk01_cellmath__39_I976 (.Y(N1946), .A0(N1805), .A1(N1802), .B0(N1804));
NAND2XL inst_blk01_cellmath__39_I977 (.Y(N1947), .A(N1805), .B(N1803));
INVXL inst_blk01_cellmath__39_I1731 (.Y(N3178), .A(N1942));
INVXL inst_blk01_cellmath__39_I1732 (.Y(N3179), .A(N1943));
OAI21XL inst_blk01_cellmath__39_I982 (.Y(N1952), .A0(N3175), .A1(N1942), .B0(N3174));
NOR2XL inst_blk01_cellmath__39_I983 (.Y(N1953), .A(N3175), .B(N1943));
OAI21XL inst_blk01_cellmath__39_I984 (.Y(N1954), .A0(N1947), .A1(N1942), .B0(N1946));
NOR2XL inst_blk01_cellmath__39_I985 (.Y(N1955), .A(N1947), .B(N1943));
AOI21XL inst_blk01_cellmath__39_I994 (.Y(N1964), .A0(N1799), .A1(N1938), .B0(N1798));
AOI21XL inst_blk01_cellmath__39_I996 (.Y(N1966), .A0(N3179), .A1(N1938), .B0(N3178));
AOI21XL inst_blk01_cellmath__39_I998 (.Y(N1968), .A0(N1953), .A1(N1938), .B0(N1952));
AOI21XL inst_blk01_cellmath__39_I1004 (.Y(N1974), .A0(N1809), .A1(N1806), .B0(N1808));
NAND2XL inst_blk01_cellmath__39_I1005 (.Y(N1975), .A(N1809), .B(N1807));
INVXL inst_blk01_cellmath__39_I1744 (.Y(N3191), .A(N1811));
AO21XL inst_blk01_cellmath__39_I1864 (.Y(N3210), .A0(N1955), .A1(N1938), .B0(N1954));
AND2XL inst_blk01_cellmath__39_I1865 (.Y(N3211), .A(N1955), .B(N1939));
INVX1 inst_blk01_cellmath__39_I1765 (.Y(N3212), .A(N1826));
AOI21X4 inst_blk01_cellmath__39_I1032 (.Y(N2002), .A0(N1843), .A1(N1826), .B0(N1842));
AOI21X4 inst_blk01_cellmath__39_I1034 (.Y(N2004), .A0(N1859), .A1(N1842), .B0(N1858));
NAND2X4 inst_blk01_cellmath__39_I1035 (.Y(N2005), .A(N1859), .B(N1843));
AOI21X4 inst_blk01_cellmath__39_I1036 (.Y(N2006), .A0(N1875), .A1(N1858), .B0(N1874));
NAND2X4 inst_blk01_cellmath__39_I1037 (.Y(N2007), .A(N1875), .B(N1859));
AOI21X4 inst_blk01_cellmath__39_I1038 (.Y(N2008), .A0(N1891), .A1(N1874), .B0(N1890));
NAND2X4 inst_blk01_cellmath__39_I1039 (.Y(N2009), .A(N1891), .B(N1875));
AOI21X4 inst_blk01_cellmath__39_I1040 (.Y(N2010), .A0(N1907), .A1(N1890), .B0(N1906));
NAND2X4 inst_blk01_cellmath__39_I1041 (.Y(N2011), .A(N1907), .B(N1891));
AOI21X2 inst_blk01_cellmath__39_I1042 (.Y(N2012), .A0(N1923), .A1(N1906), .B0(N1922));
NAND2X2 inst_blk01_cellmath__39_I1043 (.Y(N2013), .A(N1923), .B(N1907));
AOI21X1 inst_blk01_cellmath__39_I1044 (.Y(N2014), .A0(N3211), .A1(N1922), .B0(N3210));
NAND2X2 inst_blk01_cellmath__39_I1045 (.Y(N2015), .A(N3211), .B(N1923));
INVXL inst_blk01_cellmath__39_I1766 (.Y(N3213), .A(N3212));
INVXL inst_blk01_cellmath__39_I1767 (.Y(N3214), .A(N2002));
OAI21X4 inst_blk01_cellmath__39_I1050 (.Y(N2020), .A0(N2005), .A1(N3212), .B0(N2004));
OAI21X4 inst_blk01_cellmath__39_I1052 (.Y(N2022), .A0(N2007), .A1(N2002), .B0(N2006));
OAI21X2 inst_blk01_cellmath__39_I1054 (.Y(N2024), .A0(N2009), .A1(N2004), .B0(N2008));
NOR2X2 inst_blk01_cellmath__39_I1055 (.Y(N2025), .A(N2009), .B(N2005));
OAI21X2 inst_blk01_cellmath__39_I1056 (.Y(N2026), .A0(N2011), .A1(N2006), .B0(N2010));
NOR2X1 inst_blk01_cellmath__39_I1057 (.Y(N2027), .A(N2011), .B(N2007));
OAI21X2 inst_blk01_cellmath__39_I1058 (.Y(N2028), .A0(N2013), .A1(N2008), .B0(N2012));
NOR2X2 inst_blk01_cellmath__39_I1059 (.Y(N2029), .A(N2013), .B(N2009));
OAI21X2 inst_blk01_cellmath__39_I1060 (.Y(N2030), .A0(N2015), .A1(N2010), .B0(N2014));
NOR2X2 inst_blk01_cellmath__39_I1061 (.Y(N2031), .A(N2015), .B(N2011));
INVXL inst_blk01_cellmath__39_I1768 (.Y(N3215), .A(N3213));
INVXL inst_blk01_cellmath__39_I1769 (.Y(N3216), .A(N3214));
INVXL inst_blk01_cellmath__39_I1770 (.Y(N3217), .A(N2020));
INVXL inst_blk01_cellmath__39_I1771 (.Y(N3218), .A(N2022));
AOI21X2 inst_blk01_cellmath__39_I1070 (.Y(N2040), .A0(N2025), .A1(N3213), .B0(N2024));
AOI21X2 inst_blk01_cellmath__39_I1072 (.Y(N2042), .A0(N2027), .A1(N3214), .B0(N2026));
AOI21X4 inst_blk01_cellmath__39_I1074 (.Y(N2044), .A0(N2029), .A1(N2020), .B0(N2028));
AOI21X4 inst_blk01_cellmath__39_I1076 (.Y(N2046), .A0(N2031), .A1(N2022), .B0(N2030));
NOR2BX1 andori2bb1_A_I3346 (.Y(N3303), .AN(N1739), .B(N1814));
NOR2XL andori2bb1_A_I1976 (.Y(N3223), .A(N3303), .B(N1738));
NOR2XL andori2bb1_A_I1977 (.Y(N3310), .A(N3113), .B(N1830));
NOR2XL andori2bb1_A_I1978 (.Y(N3228), .A(N3310), .B(N1746));
NOR2XL andori2bb1_A_I1979 (.Y(N3317), .A(N3121), .B(N1846));
NOR2XL andori2bb1_A_I1980 (.Y(N3234), .A(N3317), .B(N1754));
NOR2XL andori2bb1_A_I1981 (.Y(N3324), .A(N3131), .B(N1862));
NOR2XL andori2bb1_A_I1982 (.Y(N3240), .A(N3324), .B(N1762));
NOR2XL andori2bb1_A_I3358 (.Y(N5103), .A(N3141), .B(N1878));
NOR2XL andori2bb1_A_I3359 (.Y(N3246), .A(N5103), .B(N1770));
NOR2XL andori2bb1_A_I1983 (.Y(N3331), .A(N3151), .B(N1894));
NOR2XL andori2bb1_A_I1984 (.Y(N3252), .A(N3331), .B(N1778));
NOR2XL andori2bb1_A_I1985 (.Y(N3338), .A(N3159), .B(N1910));
NOR2XL andori2bb1_A_I1986 (.Y(N3258), .A(N3338), .B(N1786));
NOR2XL andori2bb1_A_I1987 (.Y(N3345), .A(N3167), .B(N1926));
NOR2XL andori2bb1_A_I1988 (.Y(N3264), .A(N3345), .B(N1794));
INVXL inst_blk01_cellmath__39_I1819 (.Y(N3266), .A(N1938));
NOR2XL andori2bb1_A_I1989 (.Y(N3352), .A(N3191), .B(N1974));
NOR2XL andori2bb1_A_I1990 (.Y(N3278), .A(N3352), .B(N1810));
OR2XL inst_blk01_cellmath__39_I1883 (.Y(N3279), .A(N3191), .B(N1975));
NAND2BXL inst_blk01_cellmath__39_I1184 (.Y(N2154), .AN(N1736), .B(N1737));
NAND2BXL inst_blk01_cellmath__39_I1187 (.Y(N2157), .AN(N1738), .B(N1739));
NAND2BXL inst_blk01_cellmath__39_I1190 (.Y(N2160), .AN(N1740), .B(N1741));
NAND2BXL inst_blk01_cellmath__39_I1193 (.Y(N2163), .AN(N1742), .B(N1743));
NAND2BXL inst_blk01_cellmath__39_I1196 (.Y(N2166), .AN(N1744), .B(N1745));
NAND2BXL inst_blk01_cellmath__39_I1199 (.Y(N2601), .AN(N1746), .B(N1747));
NAND2BXL inst_blk01_cellmath__39_I1202 (.Y(N2612), .AN(N1748), .B(N1749));
NAND2BXL inst_blk01_cellmath__39_I1205 (.Y(N2175), .AN(N1750), .B(N1751));
NAND2BXL inst_blk01_cellmath__39_I1208 (.Y(N2178), .AN(N1752), .B(N1753));
NAND2BXL inst_blk01_cellmath__39_I1211 (.Y(N2630), .AN(N1754), .B(N1755));
NAND2BXL inst_blk01_cellmath__39_I1214 (.Y(N2641), .AN(N1756), .B(N1757));
NAND2BXL inst_blk01_cellmath__39_I1217 (.Y(N2187), .AN(N1758), .B(N1759));
NAND2BXL inst_blk01_cellmath__39_I1220 (.Y(N2190), .AN(N1760), .B(N1761));
NAND2BXL inst_blk01_cellmath__39_I1223 (.Y(N2659), .AN(N1762), .B(N1763));
NAND2BXL inst_blk01_cellmath__39_I1226 (.Y(N2670), .AN(N1764), .B(N1765));
NAND2BXL inst_blk01_cellmath__39_I1229 (.Y(N2199), .AN(N1766), .B(N1767));
NAND2BXL inst_blk01_cellmath__39_I1232 (.Y(N2202), .AN(N1768), .B(N1769));
NAND2BXL inst_blk01_cellmath__39_I1235 (.Y(N2688), .AN(N1770), .B(N1771));
NAND2BXL inst_blk01_cellmath__39_I1238 (.Y(N2699), .AN(N1772), .B(N1773));
NAND2BXL inst_blk01_cellmath__39_I1241 (.Y(N2211), .AN(N1774), .B(N1775));
NAND2BXL inst_blk01_cellmath__39_I1244 (.Y(N2214), .AN(N1776), .B(N1777));
NAND2BXL inst_blk01_cellmath__39_I1247 (.Y(N2717), .AN(N1778), .B(N1779));
NAND2BXL inst_blk01_cellmath__39_I1250 (.Y(N2728), .AN(N1780), .B(N1781));
NAND2BXL inst_blk01_cellmath__39_I1253 (.Y(N2223), .AN(N1782), .B(N1783));
NAND2BXL inst_blk01_cellmath__39_I1256 (.Y(N2226), .AN(N1784), .B(N1785));
NAND2BXL inst_blk01_cellmath__39_I1259 (.Y(N2746), .AN(N1786), .B(N1787));
NAND2BXL inst_blk01_cellmath__39_I1262 (.Y(N2757), .AN(N1788), .B(N1789));
NAND2BXL inst_blk01_cellmath__39_I1265 (.Y(N2235), .AN(N1790), .B(N1791));
NAND2BXL inst_blk01_cellmath__39_I1268 (.Y(N2238), .AN(N1792), .B(N1793));
NAND2BXL inst_blk01_cellmath__39_I1271 (.Y(N2775), .AN(N1794), .B(N1795));
NAND2BXL inst_blk01_cellmath__39_I1274 (.Y(N2786), .AN(N1796), .B(N1797));
NAND2BXL inst_blk01_cellmath__39_I1277 (.Y(N2797), .AN(N1798), .B(N1799));
NAND2BXL inst_blk01_cellmath__39_I1280 (.Y(N2808), .AN(N1800), .B(N1801));
NAND2BXL inst_blk01_cellmath__39_I1283 (.Y(N2819), .AN(N1802), .B(N1803));
NAND2BXL inst_blk01_cellmath__39_I1286 (.Y(N2830), .AN(N1804), .B(N1805));
NAND2BXL inst_blk01_cellmath__39_I1289 (.Y(N2259), .AN(N1806), .B(N1807));
NAND2BXL inst_blk01_cellmath__39_I1292 (.Y(N2262), .AN(N1808), .B(N1809));
NAND2BXL inst_blk01_cellmath__39_I1295 (.Y(N2848), .AN(N1810), .B(N1811));
XOR2XL inst_blk01_cellmath__39_I1884 (.Y(inst_blk01_cellmath__39_out0[16]), .A(N1734), .B(N2154));
XNOR2X1 inst_blk01_cellmath__39_I1298 (.Y(inst_blk01_cellmath__39_out0[17]), .A(N1814), .B(N2157));
XNOR2X1 inst_blk01_cellmath__39_I1299 (.Y(inst_blk01_cellmath__39_out0[18]), .A(N3223), .B(N2160));
XNOR2X1 inst_blk01_cellmath__39_I1300 (.Y(inst_blk01_cellmath__39_out0[19]), .A(N3215), .B(N2163));
XNOR2X1 inst_blk01_cellmath__39_I1301 (.Y(inst_blk01_cellmath__39_out0[23]), .A(N3216), .B(N2175));
XNOR2X1 inst_blk01_cellmath__39_I1302 (.Y(inst_blk01_cellmath__39_out0[27]), .A(N3217), .B(N2187));
XNOR2X1 inst_blk01_cellmath__39_I1303 (.Y(inst_blk01_cellmath__39_out0[31]), .A(N3218), .B(N2199));
XNOR2X1 inst_blk01_cellmath__39_I3348 (.Y(inst_blk01_cellmath__39_out0[35]), .A(N2040), .B(N2211));
XNOR2X1 inst_blk01_cellmath__39_I3349 (.Y(inst_blk01_cellmath__39_out0[39]), .A(N2042), .B(N2223));
INVX1 xnor2_A_I1444 (.Y(N2583), .A(N2044));
MXI2XL xnor2_A_I1445 (.Y(inst_blk01_cellmath__39_out0[43]), .A(N2044), .B(N2583), .S0(N2235));
XNOR2XL inst_blk01_cellmath__39_I1307 (.Y(inst_blk01_cellmath__39_out0[51]), .A(N2046), .B(N2259));
XOR2XL node_cs_reduced_ii_local_A_I1888 (.Y(N2279), .A(N2166), .B(N1743));
XOR2XL node_cs_reduced_ii_local_A_I1889 (.Y(N2278), .A(N2166), .B(N1742));
MX2XL inst_blk01_cellmath__39_I1309 (.Y(inst_blk01_cellmath__39_out0[20]), .A(N2279), .B(N2278), .S0(N3215));
XOR2XL node_cs_ii_local_alt_A_I1449 (.Y(N2281), .A(N2601), .B(N1830));
NAND2XL node_cs_ii_local_alt_A_I1450 (.Y(N2599), .A(N1831), .B(N1830));
XNOR2X1 node_cs_ii_local_alt_A_I1451 (.Y(N2282), .A(N2601), .B(N2599));
MXI2XL inst_blk01_cellmath__39_I1311 (.Y(inst_blk01_cellmath__39_out0[21]), .A(N2282), .B(N2281), .S0(N3215));
XOR2XL node_cs_ii_local_alt_A_I1453 (.Y(N2284), .A(N2612), .B(N3228));
OAI21XL node_cs_ii_local_alt_A_I1890 (.Y(N2610), .A0(N3113), .A1(N1831), .B0(N3228));
XNOR2X1 node_cs_ii_local_alt_A_I1455 (.Y(N2285), .A(N2612), .B(N2610));
MXI2XL inst_blk01_cellmath__39_I1313 (.Y(inst_blk01_cellmath__39_out0[22]), .A(N2285), .B(N2284), .S0(N3215));
XOR2XL node_cs_reduced_ii_local_A_I1891 (.Y(N2288), .A(N2178), .B(N1751));
XOR2XL node_cs_reduced_ii_local_A_I1892 (.Y(N2287), .A(N2178), .B(N1750));
MX2XL inst_blk01_cellmath__39_I1315 (.Y(inst_blk01_cellmath__39_out0[24]), .A(N2288), .B(N2287), .S0(N3216));
XOR2XL node_cs_ii_local_alt_A_I1459 (.Y(N2290), .A(N2630), .B(N1846));
NAND2XL node_cs_ii_local_alt_A_I1460 (.Y(N2628), .A(N1847), .B(N1846));
XNOR2X1 node_cs_ii_local_alt_A_I1461 (.Y(N2291), .A(N2630), .B(N2628));
MXI2XL inst_blk01_cellmath__39_I1317 (.Y(inst_blk01_cellmath__39_out0[25]), .A(N2291), .B(N2290), .S0(N3216));
XOR2XL node_cs_ii_local_alt_A_I1463 (.Y(N2293), .A(N2641), .B(N3234));
OAI21XL node_cs_ii_local_alt_A_I1893 (.Y(N2639), .A0(N3121), .A1(N1847), .B0(N3234));
XNOR2X1 node_cs_ii_local_alt_A_I1465 (.Y(N2294), .A(N2641), .B(N2639));
MXI2XL inst_blk01_cellmath__39_I1319 (.Y(inst_blk01_cellmath__39_out0[26]), .A(N2294), .B(N2293), .S0(N3216));
XOR2XL node_cs_reduced_ii_local_A_I1894 (.Y(N2297), .A(N2190), .B(N1759));
XOR2XL node_cs_reduced_ii_local_A_I1895 (.Y(N2296), .A(N2190), .B(N1758));
MX2XL inst_blk01_cellmath__39_I1321 (.Y(inst_blk01_cellmath__39_out0[28]), .A(N2297), .B(N2296), .S0(N3217));
XOR2XL node_cs_ii_local_alt_A_I1469 (.Y(N2299), .A(N2659), .B(N1862));
NAND2XL node_cs_ii_local_alt_A_I1470 (.Y(N2657), .A(N1863), .B(N1862));
XNOR2X1 node_cs_ii_local_alt_A_I1471 (.Y(N2300), .A(N2659), .B(N2657));
MXI2XL inst_blk01_cellmath__39_I1323 (.Y(inst_blk01_cellmath__39_out0[29]), .A(N2300), .B(N2299), .S0(N3217));
XOR2XL node_cs_ii_local_alt_A_I1473 (.Y(N2302), .A(N2670), .B(N3240));
OAI21XL node_cs_ii_local_alt_A_I1896 (.Y(N2668), .A0(N3131), .A1(N1863), .B0(N3240));
XNOR2X1 node_cs_ii_local_alt_A_I1475 (.Y(N2303), .A(N2670), .B(N2668));
MXI2XL inst_blk01_cellmath__39_I1325 (.Y(inst_blk01_cellmath__39_out0[30]), .A(N2303), .B(N2302), .S0(N3217));
XOR2XL node_cs_reduced_ii_local_A_I1897 (.Y(N2306), .A(N2202), .B(N1767));
XOR2XL node_cs_reduced_ii_local_A_I1898 (.Y(N2305), .A(N2202), .B(N1766));
MX2XL inst_blk01_cellmath__39_I1327 (.Y(inst_blk01_cellmath__39_out0[32]), .A(N2306), .B(N2305), .S0(N3218));
XOR2XL node_cs_ii_local_alt_A_I1479 (.Y(N2308), .A(N2688), .B(N1878));
NAND2XL node_cs_ii_local_alt_A_I1480 (.Y(N2686), .A(N1879), .B(N1878));
XNOR2X1 node_cs_ii_local_alt_A_I1481 (.Y(N2309), .A(N2688), .B(N2686));
MXI2XL inst_blk01_cellmath__39_I1329 (.Y(inst_blk01_cellmath__39_out0[33]), .A(N2309), .B(N2308), .S0(N3218));
XOR2XL node_cs_ii_local_alt_A_I1483 (.Y(N2311), .A(N2699), .B(N3246));
OAI21XL node_cs_ii_local_alt_A_I1959 (.Y(N2697), .A0(N3141), .A1(N1879), .B0(N3246));
XNOR2X1 node_cs_ii_local_alt_A_I1485 (.Y(N2312), .A(N2699), .B(N2697));
MXI2XL inst_blk01_cellmath__39_I1331 (.Y(inst_blk01_cellmath__39_out0[34]), .A(N2312), .B(N2311), .S0(N3218));
XOR2XL node_cs_reduced_ii_local_A_I1900 (.Y(N2315), .A(N2214), .B(N1775));
XOR2XL node_cs_reduced_ii_local_A_I1901 (.Y(N2314), .A(N2214), .B(N1774));
MX2XL inst_blk01_cellmath__39_I1333 (.Y(inst_blk01_cellmath__39_out0[36]), .A(N2315), .B(N2314), .S0(N2040));
XOR2XL node_cs_ii_local_alt_A_I1489 (.Y(N2317), .A(N2717), .B(N1894));
NAND2XL node_cs_ii_local_alt_A_I1490 (.Y(N2715), .A(N1895), .B(N1894));
XNOR2X1 node_cs_ii_local_alt_A_I1491 (.Y(N2318), .A(N2717), .B(N2715));
MXI2XL inst_blk01_cellmath__39_I1335 (.Y(inst_blk01_cellmath__39_out0[37]), .A(N2318), .B(N2317), .S0(N2040));
XOR2XL node_cs_ii_local_alt_A_I1493 (.Y(N2320), .A(N2728), .B(N3252));
OAI21XL node_cs_ii_local_alt_A_I1902 (.Y(N2726), .A0(N3151), .A1(N1895), .B0(N3252));
XNOR2X1 node_cs_ii_local_alt_A_I1495 (.Y(N2321), .A(N2728), .B(N2726));
MXI2XL inst_blk01_cellmath__39_I1337 (.Y(inst_blk01_cellmath__39_out0[38]), .A(N2321), .B(N2320), .S0(N2040));
XOR2XL node_cs_reduced_ii_local_A_I1903 (.Y(N2324), .A(N2226), .B(N1783));
XOR2XL node_cs_reduced_ii_local_A_I1904 (.Y(N2323), .A(N2226), .B(N1782));
MX2XL inst_blk01_cellmath__39_I1339 (.Y(inst_blk01_cellmath__39_out0[40]), .A(N2324), .B(N2323), .S0(N2042));
XOR2XL node_cs_ii_local_alt_A_I1499 (.Y(N2326), .A(N2746), .B(N1910));
NAND2XL node_cs_ii_local_alt_A_I1500 (.Y(N2744), .A(N1911), .B(N1910));
XNOR2X1 node_cs_ii_local_alt_A_I1501 (.Y(N2327), .A(N2746), .B(N2744));
MXI2XL inst_blk01_cellmath__39_I1341 (.Y(inst_blk01_cellmath__39_out0[41]), .A(N2327), .B(N2326), .S0(N2042));
XOR2XL node_cs_ii_local_alt_A_I1503 (.Y(N2329), .A(N2757), .B(N3258));
OAI21XL node_cs_ii_local_alt_A_I1905 (.Y(N2755), .A0(N3159), .A1(N1911), .B0(N3258));
XNOR2X1 node_cs_ii_local_alt_A_I1505 (.Y(N2330), .A(N2757), .B(N2755));
MXI2XL inst_blk01_cellmath__39_I1343 (.Y(inst_blk01_cellmath__39_out0[42]), .A(N2330), .B(N2329), .S0(N2042));
XOR2XL node_cs_reduced_ii_local_A_I1906 (.Y(N2333), .A(N2238), .B(N1791));
XOR2XL node_cs_reduced_ii_local_A_I1907 (.Y(N2332), .A(N2238), .B(N1790));
MX2XL inst_blk01_cellmath__39_I1345 (.Y(inst_blk01_cellmath__39_out0[44]), .A(N2333), .B(N2332), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1509 (.Y(N2335), .A(N2775), .B(N1926));
NAND2XL node_cs_ii_local_alt_A_I1510 (.Y(N2773), .A(N1927), .B(N1926));
XNOR2X1 node_cs_ii_local_alt_A_I1511 (.Y(N2336), .A(N2775), .B(N2773));
MXI2XL inst_blk01_cellmath__39_I1347 (.Y(inst_blk01_cellmath__39_out0[45]), .A(N2336), .B(N2335), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1513 (.Y(N2338), .A(N2786), .B(N3264));
OAI21XL node_cs_ii_local_alt_A_I1908 (.Y(N2784), .A0(N3167), .A1(N1927), .B0(N3264));
XNOR2X1 node_cs_ii_local_alt_A_I1515 (.Y(N2339), .A(N2786), .B(N2784));
MXI2XL inst_blk01_cellmath__39_I1349 (.Y(inst_blk01_cellmath__39_out0[46]), .A(N2339), .B(N2338), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1517 (.Y(N2341), .A(N2797), .B(N3266));
NAND2BXL node_cs_ii_local_alt_A_I1909 (.Y(N2795), .AN(N1939), .B(N3266));
XNOR2X1 node_cs_ii_local_alt_A_I1519 (.Y(N2342), .A(N2797), .B(N2795));
MXI2XL inst_blk01_cellmath__39_I1351 (.Y(inst_blk01_cellmath__39_out0[47]), .A(N2342), .B(N2341), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1521 (.Y(N2344), .A(N2808), .B(N1964));
OAI2BB1X1 node_cs_ii_local_alt_A_I1910 (.Y(N2806), .A0N(N1799), .A1N(N1939), .B0(N1964));
XNOR2X1 node_cs_ii_local_alt_A_I1523 (.Y(N2345), .A(N2808), .B(N2806));
MXI2XL inst_blk01_cellmath__39_I1353 (.Y(inst_blk01_cellmath__39_out0[48]), .A(N2345), .B(N2344), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1525 (.Y(N2347), .A(N2819), .B(N1966));
OAI2BB1X1 node_cs_ii_local_alt_A_I1911 (.Y(N2817), .A0N(N3179), .A1N(N1939), .B0(N1966));
XNOR2X1 node_cs_ii_local_alt_A_I1527 (.Y(N2348), .A(N2819), .B(N2817));
MXI2XL inst_blk01_cellmath__39_I1355 (.Y(inst_blk01_cellmath__39_out0[49]), .A(N2348), .B(N2347), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1529 (.Y(N2350), .A(N2830), .B(N1968));
OAI2BB1X1 node_cs_ii_local_alt_A_I1912 (.Y(N2828), .A0N(N1953), .A1N(N1939), .B0(N1968));
XNOR2X1 node_cs_ii_local_alt_A_I1531 (.Y(N2351), .A(N2830), .B(N2828));
MXI2XL inst_blk01_cellmath__39_I1357 (.Y(inst_blk01_cellmath__39_out0[50]), .A(N2351), .B(N2350), .S0(N2044));
XOR2XL node_cs_reduced_ii_local_A_I1913 (.Y(N2354), .A(N2262), .B(N1807));
XOR2XL node_cs_reduced_ii_local_A_I1914 (.Y(N2353), .A(N2262), .B(N1806));
MX2XL inst_blk01_cellmath__39_I1359 (.Y(inst_blk01_cellmath__39_out0[52]), .A(N2354), .B(N2353), .S0(N2046));
XOR2XL node_cs_ii_local_alt_A_I1535 (.Y(N2356), .A(N2848), .B(N1974));
NAND2XL node_cs_ii_local_alt_A_I1536 (.Y(N2846), .A(N1975), .B(N1974));
XNOR2X1 node_cs_ii_local_alt_A_I1537 (.Y(N2357), .A(N2848), .B(N2846));
MXI2XL inst_blk01_cellmath__39_I1361 (.Y(inst_blk01_cellmath__39_out0[53]), .A(N2357), .B(N2356), .S0(N2046));
OA21X1 inst_blk01_cellmath__39_I1560 (.Y(inst_blk01_cellmath__39_out0[55]), .A0(N3279), .A1(N2046), .B0(N3278));
INVXL inst_blk01_cellmath__39_I1833 (.Y(inst_blk01_cellmath__39_out0[54]), .A(inst_blk01_cellmath__39_out0[55]));
assign inst_blk01_cellmath__39_out0[0] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__42_0_bdw1157874770_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0
	); /* architecture "gate_level" */ 
output [8:0] inst_cellmath__42_0_out0;
input [7:0] inst_cellmath__42_0_in0;
wire N32,N36,N38,N63,N72,N84,N200 
	,N201,N202,N203,N217,N224,N231,N238,N245 
	;
INVX2 inst_cellmath__42_0_I5 (.Y(inst_cellmath__42_0_out0[0]), .A(inst_cellmath__42_0_in0[0]));
INVXL inst_cellmath__42_0_I107 (.Y(N200), .A(inst_cellmath__42_0_in0[1]));
INVXL inst_cellmath__42_0_I108 (.Y(N201), .A(inst_cellmath__42_0_in0[2]));
INVXL inst_cellmath__42_0_I8 (.Y(N32), .A(inst_cellmath__42_0_in0[3]));
INVXL inst_cellmath__42_0_I109 (.Y(N202), .A(inst_cellmath__42_0_in0[4]));
INVXL inst_cellmath__42_0_I10 (.Y(N36), .A(inst_cellmath__42_0_in0[5]));
INVXL inst_cellmath__42_0_I11 (.Y(N38), .A(inst_cellmath__42_0_in0[6]));
OAI21XL inst_cellmath__42_0_I31 (.Y(N63), .A0(N201), .A1(N200), .B0(N32));
NAND3XL inst_cellmath__42_0_I38 (.Y(N72), .A(N38), .B(N36), .C(N202));
INVXL inst_cellmath__42_0_I129 (.Y(N203), .A(inst_cellmath__42_0_in0[7]));
NAND2XL hyperpropagate_3_1_A_I132 (.Y(N217), .A(N36), .B(N202));
NOR2XL hyperpropagate_3_1_A_I133 (.Y(N84), .A(N63), .B(N217));
INVXL inst_cellmath__42_0_I117 (.Y(inst_cellmath__42_0_out0[1]), .A(N200));
MXI2XL inst_cellmath__42_0_I91 (.Y(inst_cellmath__42_0_out0[2]), .A(N200), .B(inst_cellmath__42_0_out0[1]), .S0(N201));
NOR2XL node_cs_const1_cs_A_I134 (.Y(N224), .A(N201), .B(N200));
XNOR2X1 node_cs_const1_cs_A_I135 (.Y(inst_cellmath__42_0_out0[3]), .A(N32), .B(N224));
XNOR2X1 inst_cellmath__42_0_I105 (.Y(inst_cellmath__42_0_out0[4]), .A(N63), .B(N202));
NOR2XL node_cs_const1_cs_A_I136 (.Y(N231), .A(inst_cellmath__42_0_in0[4]), .B(N63));
XOR2XL node_cs_const1_cs_A_I194 (.Y(inst_cellmath__42_0_out0[5]), .A(N36), .B(N231));
XOR2XL inst_cellmath__42_0_I126 (.Y(inst_cellmath__42_0_out0[6]), .A(N84), .B(N38));
NOR2XL node_cs_const1_cs_A_I138 (.Y(N238), .A(N72), .B(N63));
XNOR2X1 node_cs_const1_cs_A_I139 (.Y(inst_cellmath__42_0_out0[7]), .A(N203), .B(N238));
NOR2XL andori2bb1_A_I140 (.Y(N245), .A(N72), .B(N63));
NOR2XL andori2bb1_A_I141 (.Y(inst_cellmath__42_0_out0[8]), .A(N245), .B(N203));
endmodule

module cynw_cm_float_cos_inst_cellmath__48_bdw1157874770_bdw (
	inst_cellmath__48_out0,
	inst_cellmath__48_in0,
	inst_cellmath__48_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__48_out0;
input [5:0] inst_cellmath__48_in0;
input [55:26] inst_cellmath__48_in1;
wire N65,N66,N67,N68,N69,N70,N71 
	,N72,N73,N74,N75,N76,N77,N78,N79 
	,N80,N81,N82,N83,N84,N85,N86,N87 
	,N88,N89,N90,N91,N92,N93,N94,N130 
	,N131,N132,N133,N134,N135,N136,N137,N138 
	,N139,N140,N141,N142,N143,N144,N145,N146 
	,N147,N148,N149,N150,N151,N152,N153,N154 
	,N155,N156,N157,N158,N160,N196,N197,N198 
	,N199,N200,N201,N202,N203,N204,N205,N206 
	,N207,N208,N209,N210,N211,N212,N213,N214 
	,N215,N216,N217,N218,N219,N220,N221,N222 
	,N224,N226,N228,N264,N265,N266,N267,N268 
	,N269,N270,N271,N272,N273,N274,N275,N276 
	,N277,N278,N279,N280,N281,N282,N283,N284 
	,N285,N286,N288,N290,N292,N294,N296,N298 
	,N300,N336,N337,N338,N339,N340,N341,N342 
	,N343,N344,N345,N346,N347,N348,N349,N350 
	,N352,N354,N356,N358,N360,N362,N364,N366 
	,N368,N370,N508,N509,N510,N511,N512,N513 
	,N514,N515,N516,N517,N518,N519,N520,N521 
	,N522,N523,N524,N525,N526,N527,N528,N529 
	,N530,N531,N532,N533,N534,N535,N536,N537 
	,N538,N539,N540,N541,N542,N543,N544,N545 
	,N546,N547,N549,N550,N551,N552,N553,N554 
	,N555,N556;
INVXL inst_cellmath__48_I384 (.Y(N508), .A(inst_cellmath__48_in0[0]));
INVXL inst_cellmath__48_I385 (.Y(N509), .A(N508));
INVXL inst_cellmath__48_I391 (.Y(N515), .A(N509));
INVXL inst_cellmath__48_I390 (.Y(N514), .A(N509));
INVXL inst_cellmath__48_I389 (.Y(N513), .A(N509));
INVXL inst_cellmath__48_I388 (.Y(N512), .A(N509));
INVXL inst_cellmath__48_I387 (.Y(N511), .A(N509));
INVXL inst_cellmath__48_I386 (.Y(N510), .A(N509));
MXI2XL inst_cellmath__48_I2 (.Y(N65), .A(inst_cellmath__48_in1[27]), .B(inst_cellmath__48_in1[26]), .S0(N515));
MXI2XL inst_cellmath__48_I3 (.Y(N66), .A(inst_cellmath__48_in1[28]), .B(inst_cellmath__48_in1[27]), .S0(N515));
MXI2XL inst_cellmath__48_I4 (.Y(N67), .A(inst_cellmath__48_in1[29]), .B(inst_cellmath__48_in1[28]), .S0(N515));
MXI2XL inst_cellmath__48_I5 (.Y(N68), .A(inst_cellmath__48_in1[30]), .B(inst_cellmath__48_in1[29]), .S0(N515));
MXI2XL inst_cellmath__48_I6 (.Y(N69), .A(inst_cellmath__48_in1[31]), .B(inst_cellmath__48_in1[30]), .S0(N515));
MXI2XL inst_cellmath__48_I7 (.Y(N70), .A(inst_cellmath__48_in1[32]), .B(inst_cellmath__48_in1[31]), .S0(N514));
MXI2XL inst_cellmath__48_I8 (.Y(N71), .A(inst_cellmath__48_in1[33]), .B(inst_cellmath__48_in1[32]), .S0(N514));
MXI2XL inst_cellmath__48_I9 (.Y(N72), .A(inst_cellmath__48_in1[34]), .B(inst_cellmath__48_in1[33]), .S0(N514));
MXI2XL inst_cellmath__48_I10 (.Y(N73), .A(inst_cellmath__48_in1[35]), .B(inst_cellmath__48_in1[34]), .S0(N514));
MXI2XL inst_cellmath__48_I11 (.Y(N74), .A(inst_cellmath__48_in1[36]), .B(inst_cellmath__48_in1[35]), .S0(N514));
MXI2XL inst_cellmath__48_I12 (.Y(N75), .A(inst_cellmath__48_in1[37]), .B(inst_cellmath__48_in1[36]), .S0(N513));
MXI2XL inst_cellmath__48_I13 (.Y(N76), .A(inst_cellmath__48_in1[38]), .B(inst_cellmath__48_in1[37]), .S0(N513));
MXI2XL inst_cellmath__48_I14 (.Y(N77), .A(inst_cellmath__48_in1[39]), .B(inst_cellmath__48_in1[38]), .S0(N513));
MXI2XL inst_cellmath__48_I15 (.Y(N78), .A(inst_cellmath__48_in1[40]), .B(inst_cellmath__48_in1[39]), .S0(N513));
MXI2XL inst_cellmath__48_I16 (.Y(N79), .A(inst_cellmath__48_in1[41]), .B(inst_cellmath__48_in1[40]), .S0(N513));
MXI2XL inst_cellmath__48_I17 (.Y(N80), .A(inst_cellmath__48_in1[42]), .B(inst_cellmath__48_in1[41]), .S0(N512));
MXI2XL inst_cellmath__48_I18 (.Y(N81), .A(inst_cellmath__48_in1[43]), .B(inst_cellmath__48_in1[42]), .S0(N512));
MXI2XL inst_cellmath__48_I19 (.Y(N82), .A(inst_cellmath__48_in1[44]), .B(inst_cellmath__48_in1[43]), .S0(N512));
MXI2XL inst_cellmath__48_I20 (.Y(N83), .A(inst_cellmath__48_in1[45]), .B(inst_cellmath__48_in1[44]), .S0(N512));
MXI2XL inst_cellmath__48_I21 (.Y(N84), .A(inst_cellmath__48_in1[46]), .B(inst_cellmath__48_in1[45]), .S0(N512));
MXI2XL inst_cellmath__48_I22 (.Y(N85), .A(inst_cellmath__48_in1[47]), .B(inst_cellmath__48_in1[46]), .S0(N511));
MXI2XL inst_cellmath__48_I23 (.Y(N86), .A(inst_cellmath__48_in1[48]), .B(inst_cellmath__48_in1[47]), .S0(N511));
MXI2X1 inst_cellmath__48_I24 (.Y(N87), .A(inst_cellmath__48_in1[49]), .B(inst_cellmath__48_in1[48]), .S0(N511));
MXI2X1 inst_cellmath__48_I25 (.Y(N88), .A(inst_cellmath__48_in1[50]), .B(inst_cellmath__48_in1[49]), .S0(N511));
MXI2X1 inst_cellmath__48_I26 (.Y(N89), .A(inst_cellmath__48_in1[51]), .B(inst_cellmath__48_in1[50]), .S0(N511));
MXI2X1 inst_cellmath__48_I27 (.Y(N90), .A(inst_cellmath__48_in1[52]), .B(inst_cellmath__48_in1[51]), .S0(N510));
MXI2X1 inst_cellmath__48_I28 (.Y(N91), .A(inst_cellmath__48_in1[53]), .B(inst_cellmath__48_in1[52]), .S0(N510));
MXI2X1 inst_cellmath__48_I29 (.Y(N92), .A(inst_cellmath__48_in1[54]), .B(inst_cellmath__48_in1[53]), .S0(N510));
MXI2X1 inst_cellmath__48_I30 (.Y(N93), .A(inst_cellmath__48_in1[55]), .B(inst_cellmath__48_in1[54]), .S0(N510));
NAND2XL inst_cellmath__48_I31 (.Y(N94), .A(inst_cellmath__48_in1[55]), .B(N510));
INVXL inst_cellmath__48_I392 (.Y(N516), .A(inst_cellmath__48_in0[1]));
INVXL inst_cellmath__48_I398 (.Y(N522), .A(N516));
INVXL inst_cellmath__48_I397 (.Y(N521), .A(N516));
INVXL inst_cellmath__48_I396 (.Y(N520), .A(N516));
INVXL inst_cellmath__48_I395 (.Y(N519), .A(N516));
INVXL inst_cellmath__48_I394 (.Y(N518), .A(N516));
INVXL inst_cellmath__48_I393 (.Y(N517), .A(N516));
MXI2XL inst_cellmath__48_I66 (.Y(N130), .A(N65), .B(N67), .S0(N522));
MXI2XL inst_cellmath__48_I67 (.Y(N131), .A(N66), .B(N68), .S0(N522));
MXI2XL inst_cellmath__48_I68 (.Y(N132), .A(N67), .B(N69), .S0(N522));
MXI2XL inst_cellmath__48_I69 (.Y(N133), .A(N68), .B(N70), .S0(N522));
MXI2XL inst_cellmath__48_I70 (.Y(N134), .A(N69), .B(N71), .S0(N522));
MXI2XL inst_cellmath__48_I71 (.Y(N135), .A(N70), .B(N72), .S0(N521));
MXI2XL inst_cellmath__48_I72 (.Y(N136), .A(N71), .B(N73), .S0(N521));
MXI2XL inst_cellmath__48_I73 (.Y(N137), .A(N72), .B(N74), .S0(N521));
MXI2XL inst_cellmath__48_I74 (.Y(N138), .A(N73), .B(N75), .S0(N521));
MXI2XL inst_cellmath__48_I75 (.Y(N139), .A(N74), .B(N76), .S0(N521));
MXI2XL inst_cellmath__48_I76 (.Y(N140), .A(N75), .B(N77), .S0(N520));
MXI2XL inst_cellmath__48_I77 (.Y(N141), .A(N76), .B(N78), .S0(N520));
MXI2XL inst_cellmath__48_I78 (.Y(N142), .A(N77), .B(N79), .S0(N520));
MXI2XL inst_cellmath__48_I79 (.Y(N143), .A(N78), .B(N80), .S0(N520));
MXI2XL inst_cellmath__48_I80 (.Y(N144), .A(N79), .B(N81), .S0(N520));
MXI2XL inst_cellmath__48_I81 (.Y(N145), .A(N80), .B(N82), .S0(N519));
MXI2XL inst_cellmath__48_I82 (.Y(N146), .A(N81), .B(N83), .S0(N519));
MXI2XL inst_cellmath__48_I83 (.Y(N147), .A(N82), .B(N84), .S0(N519));
MXI2XL inst_cellmath__48_I84 (.Y(N148), .A(N83), .B(N85), .S0(N519));
MXI2X1 inst_cellmath__48_I85 (.Y(N149), .A(N84), .B(N86), .S0(N519));
MXI2X1 inst_cellmath__48_I86 (.Y(N150), .A(N85), .B(N87), .S0(N518));
MXI2XL inst_cellmath__48_I87 (.Y(N151), .A(N86), .B(N88), .S0(N518));
MXI2XL inst_cellmath__48_I88 (.Y(N152), .A(N87), .B(N89), .S0(N518));
MXI2X1 inst_cellmath__48_I89 (.Y(N153), .A(N88), .B(N90), .S0(N518));
MXI2XL inst_cellmath__48_I90 (.Y(N154), .A(N89), .B(N91), .S0(N518));
MXI2XL inst_cellmath__48_I91 (.Y(N155), .A(N90), .B(N92), .S0(N517));
MXI2XL inst_cellmath__48_I92 (.Y(N156), .A(N91), .B(N93), .S0(N517));
MXI2X1 inst_cellmath__48_I93 (.Y(N157), .A(N92), .B(N94), .S0(N517));
NOR2XL inst_cellmath__48_I94 (.Y(N158), .A(N93), .B(N517));
NOR2XL inst_cellmath__48_I95 (.Y(N160), .A(N94), .B(N517));
INVXL inst_cellmath__48_I399 (.Y(N523), .A(inst_cellmath__48_in0[2]));
INVXL inst_cellmath__48_I400 (.Y(N524), .A(N523));
INVXL inst_cellmath__48_I406 (.Y(N530), .A(N524));
INVXL inst_cellmath__48_I405 (.Y(N529), .A(N524));
INVXL inst_cellmath__48_I404 (.Y(N528), .A(N524));
INVXL inst_cellmath__48_I403 (.Y(N527), .A(N524));
INVXL inst_cellmath__48_I402 (.Y(N526), .A(N524));
INVXL inst_cellmath__48_I401 (.Y(N525), .A(N524));
MXI2XL inst_cellmath__48_I130 (.Y(N196), .A(N134), .B(N130), .S0(N530));
MXI2XL inst_cellmath__48_I131 (.Y(N197), .A(N135), .B(N131), .S0(N530));
MXI2XL inst_cellmath__48_I132 (.Y(N198), .A(N136), .B(N132), .S0(N530));
MXI2XL inst_cellmath__48_I133 (.Y(N199), .A(N137), .B(N133), .S0(N530));
MXI2XL inst_cellmath__48_I134 (.Y(N200), .A(N138), .B(N134), .S0(N530));
MXI2XL inst_cellmath__48_I135 (.Y(N201), .A(N139), .B(N135), .S0(N529));
MXI2XL inst_cellmath__48_I136 (.Y(N202), .A(N140), .B(N136), .S0(N529));
MXI2XL inst_cellmath__48_I137 (.Y(N203), .A(N141), .B(N137), .S0(N529));
MXI2XL inst_cellmath__48_I138 (.Y(N204), .A(N142), .B(N138), .S0(N529));
MXI2XL inst_cellmath__48_I139 (.Y(N205), .A(N143), .B(N139), .S0(N529));
MXI2XL inst_cellmath__48_I140 (.Y(N206), .A(N144), .B(N140), .S0(N528));
MXI2XL inst_cellmath__48_I141 (.Y(N207), .A(N145), .B(N141), .S0(N528));
MXI2XL inst_cellmath__48_I142 (.Y(N208), .A(N146), .B(N142), .S0(N528));
MXI2XL inst_cellmath__48_I143 (.Y(N209), .A(N147), .B(N143), .S0(N528));
MXI2XL inst_cellmath__48_I144 (.Y(N210), .A(N148), .B(N144), .S0(N528));
MXI2X1 inst_cellmath__48_I145 (.Y(N211), .A(N149), .B(N145), .S0(N527));
MXI2X1 inst_cellmath__48_I146 (.Y(N212), .A(N150), .B(N146), .S0(N527));
MXI2X1 inst_cellmath__48_I147 (.Y(N213), .A(N151), .B(N147), .S0(N527));
MXI2X1 inst_cellmath__48_I148 (.Y(N214), .A(N152), .B(N148), .S0(N527));
MXI2XL inst_cellmath__48_I149 (.Y(N215), .A(N153), .B(N149), .S0(N527));
MXI2XL inst_cellmath__48_I150 (.Y(N216), .A(N154), .B(N150), .S0(N526));
MXI2XL inst_cellmath__48_I151 (.Y(N217), .A(N155), .B(N151), .S0(N526));
MXI2XL inst_cellmath__48_I152 (.Y(N218), .A(N156), .B(N152), .S0(N526));
MXI2X1 inst_cellmath__48_I153 (.Y(N219), .A(N157), .B(N153), .S0(N526));
MXI2XL inst_cellmath__48_I154 (.Y(N220), .A(N158), .B(N154), .S0(N526));
MXI2XL inst_cellmath__48_I155 (.Y(N221), .A(N160), .B(N155), .S0(N525));
NAND2XL inst_cellmath__48_I156 (.Y(N222), .A(N156), .B(N525));
NAND2XL inst_cellmath__48_I157 (.Y(N224), .A(N157), .B(N525));
NAND2XL inst_cellmath__48_I158 (.Y(N226), .A(N158), .B(N525));
NAND2XL inst_cellmath__48_I159 (.Y(N228), .A(N160), .B(N525));
INVXL inst_cellmath__48_I407 (.Y(N531), .A(inst_cellmath__48_in0[3]));
INVXL inst_cellmath__48_I408 (.Y(N532), .A(N531));
INVXL inst_cellmath__48_I415 (.Y(N539), .A(N532));
INVXL inst_cellmath__48_I409 (.Y(N533), .A(N532));
INVXL inst_cellmath__48_I416 (.Y(N540), .A(N539));
INVXL inst_cellmath__48_I414 (.Y(N538), .A(N533));
INVXL inst_cellmath__48_I413 (.Y(N537), .A(N533));
INVXL inst_cellmath__48_I412 (.Y(N536), .A(N533));
INVXL inst_cellmath__48_I411 (.Y(N535), .A(N533));
INVXL inst_cellmath__48_I410 (.Y(N534), .A(N533));
MXI2XL inst_cellmath__48_I194 (.Y(N264), .A(N196), .B(N204), .S0(N540));
MXI2XL inst_cellmath__48_I195 (.Y(N265), .A(N197), .B(N205), .S0(N540));
MXI2XL inst_cellmath__48_I196 (.Y(N266), .A(N198), .B(N206), .S0(N540));
MXI2XL inst_cellmath__48_I197 (.Y(N267), .A(N199), .B(N207), .S0(N540));
MXI2XL inst_cellmath__48_I198 (.Y(N268), .A(N200), .B(N208), .S0(N540));
MXI2XL inst_cellmath__48_I199 (.Y(N269), .A(N201), .B(N209), .S0(N538));
MXI2XL inst_cellmath__48_I200 (.Y(N270), .A(N202), .B(N210), .S0(N538));
MXI2XL inst_cellmath__48_I201 (.Y(N271), .A(N203), .B(N211), .S0(N538));
MXI2X1 inst_cellmath__48_I202 (.Y(N272), .A(N204), .B(N212), .S0(N538));
MXI2X1 inst_cellmath__48_I203 (.Y(N273), .A(N205), .B(N213), .S0(N538));
MXI2X1 inst_cellmath__48_I204 (.Y(N274), .A(N206), .B(N214), .S0(N537));
MXI2XL inst_cellmath__48_I205 (.Y(N275), .A(N207), .B(N215), .S0(N537));
MXI2XL inst_cellmath__48_I206 (.Y(N276), .A(N208), .B(N216), .S0(N537));
MXI2XL inst_cellmath__48_I207 (.Y(N277), .A(N209), .B(N217), .S0(N537));
MXI2XL inst_cellmath__48_I208 (.Y(N278), .A(N210), .B(N218), .S0(N537));
MXI2XL inst_cellmath__48_I209 (.Y(N279), .A(N211), .B(N219), .S0(N536));
MXI2XL inst_cellmath__48_I210 (.Y(N280), .A(N212), .B(N220), .S0(N536));
MXI2XL inst_cellmath__48_I211 (.Y(N281), .A(N213), .B(N221), .S0(N536));
MXI2X1 inst_cellmath__48_I212 (.Y(N282), .A(N214), .B(N222), .S0(N536));
MXI2XL inst_cellmath__48_I213 (.Y(N283), .A(N215), .B(N224), .S0(N536));
MXI2XL inst_cellmath__48_I214 (.Y(N284), .A(N216), .B(N226), .S0(N535));
MXI2XL inst_cellmath__48_I215 (.Y(N285), .A(N217), .B(N228), .S0(N535));
NOR2XL inst_cellmath__48_I216 (.Y(N286), .A(N218), .B(N535));
NOR2X1 inst_cellmath__48_I217 (.Y(N288), .A(N219), .B(N535));
NOR2XL inst_cellmath__48_I218 (.Y(N290), .A(N220), .B(N535));
NOR2XL inst_cellmath__48_I219 (.Y(N292), .A(N221), .B(N534));
NOR2XL inst_cellmath__48_I220 (.Y(N294), .A(N222), .B(N534));
NOR2XL inst_cellmath__48_I221 (.Y(N296), .A(N224), .B(N534));
NOR2XL inst_cellmath__48_I222 (.Y(N298), .A(N226), .B(N534));
NOR2XL inst_cellmath__48_I223 (.Y(N300), .A(N228), .B(N534));
INVXL inst_cellmath__48_I417 (.Y(N541), .A(inst_cellmath__48_in0[4]));
INVXL inst_cellmath__48_I418 (.Y(N542), .A(N541));
INVXL inst_cellmath__48_I423 (.Y(N547), .A(N542));
INVXL inst_cellmath__48_I422 (.Y(N546), .A(N542));
INVXL inst_cellmath__48_I421 (.Y(N545), .A(N542));
INVXL inst_cellmath__48_I420 (.Y(N544), .A(N542));
INVXL inst_cellmath__48_I419 (.Y(N543), .A(N542));
MXI2XL inst_cellmath__48_I258 (.Y(N336), .A(N280), .B(N264), .S0(N547));
MXI2XL inst_cellmath__48_I259 (.Y(N337), .A(N281), .B(N265), .S0(N547));
MXI2X1 inst_cellmath__48_I260 (.Y(N338), .A(N282), .B(N266), .S0(N547));
MXI2XL inst_cellmath__48_I261 (.Y(N339), .A(N283), .B(N267), .S0(N547));
MXI2XL inst_cellmath__48_I262 (.Y(N340), .A(N284), .B(N268), .S0(N547));
MXI2X1 inst_cellmath__48_I263 (.Y(N341), .A(N285), .B(N269), .S0(N546));
MXI2XL inst_cellmath__48_I264 (.Y(N342), .A(N286), .B(N270), .S0(N546));
MXI2X2 inst_cellmath__48_I265 (.Y(N343), .A(N288), .B(N271), .S0(N546));
MXI2X1 inst_cellmath__48_I266 (.Y(N344), .A(N290), .B(N272), .S0(N546));
MXI2X1 inst_cellmath__48_I267 (.Y(N345), .A(N292), .B(N273), .S0(N546));
MXI2X1 inst_cellmath__48_I268 (.Y(N346), .A(N294), .B(N274), .S0(N545));
MXI2XL inst_cellmath__48_I269 (.Y(N347), .A(N296), .B(N275), .S0(N545));
MXI2X1 inst_cellmath__48_I270 (.Y(N348), .A(N298), .B(N276), .S0(N545));
MXI2X1 inst_cellmath__48_I271 (.Y(N349), .A(N300), .B(N277), .S0(N545));
NAND2XL inst_cellmath__48_I272 (.Y(N350), .A(N278), .B(N545));
NAND2XL inst_cellmath__48_I273 (.Y(N352), .A(N279), .B(N544));
NAND2XL inst_cellmath__48_I274 (.Y(N354), .A(N280), .B(N544));
NAND2XL inst_cellmath__48_I275 (.Y(N356), .A(N281), .B(N544));
NAND2XL inst_cellmath__48_I276 (.Y(N358), .A(N282), .B(N544));
NAND2XL inst_cellmath__48_I277 (.Y(N360), .A(N283), .B(N544));
NAND2XL inst_cellmath__48_I278 (.Y(N362), .A(N284), .B(N543));
NAND2XL inst_cellmath__48_I279 (.Y(N364), .A(N285), .B(N543));
NAND2XL inst_cellmath__48_I280 (.Y(N366), .A(N286), .B(N543));
NAND2X2 inst_cellmath__48_I281 (.Y(N368), .A(N288), .B(N543));
NAND2XL inst_cellmath__48_I282 (.Y(N370), .A(N290), .B(N543));
INVXL inst_cellmath__48_I425 (.Y(N549), .A(inst_cellmath__48_in0[5]));
INVXL inst_cellmath__48_I426 (.Y(N550), .A(N549));
INVXL inst_cellmath__48_I427 (.Y(N551), .A(N550));
INVXL inst_cellmath__48_I432 (.Y(N556), .A(N551));
INVXL inst_cellmath__48_I431 (.Y(N555), .A(N551));
INVXL inst_cellmath__48_I430 (.Y(N554), .A(N551));
INVXL inst_cellmath__48_I429 (.Y(N553), .A(N551));
INVXL inst_cellmath__48_I428 (.Y(N552), .A(N551));
NOR2XL inst_cellmath__48_I322 (.Y(inst_cellmath__48_out0[0]), .A(N336), .B(N556));
NOR2XL inst_cellmath__48_I323 (.Y(inst_cellmath__48_out0[1]), .A(N337), .B(N556));
NOR2X1 inst_cellmath__48_I324 (.Y(inst_cellmath__48_out0[2]), .A(N338), .B(N556));
NOR2XL inst_cellmath__48_I325 (.Y(inst_cellmath__48_out0[3]), .A(N339), .B(N556));
NOR2XL inst_cellmath__48_I326 (.Y(inst_cellmath__48_out0[4]), .A(N340), .B(N556));
NOR2X1 inst_cellmath__48_I327 (.Y(inst_cellmath__48_out0[5]), .A(N341), .B(N555));
NOR2XL inst_cellmath__48_I328 (.Y(inst_cellmath__48_out0[6]), .A(N342), .B(N555));
NOR2X2 inst_cellmath__48_I329 (.Y(inst_cellmath__48_out0[7]), .A(N343), .B(N555));
NOR2X1 inst_cellmath__48_I330 (.Y(inst_cellmath__48_out0[8]), .A(N344), .B(N555));
NOR2X2 inst_cellmath__48_I331 (.Y(inst_cellmath__48_out0[9]), .A(N345), .B(N555));
NOR2X1 inst_cellmath__48_I332 (.Y(inst_cellmath__48_out0[10]), .A(N346), .B(N554));
NOR2XL inst_cellmath__48_I333 (.Y(inst_cellmath__48_out0[11]), .A(N347), .B(N554));
NOR2X1 inst_cellmath__48_I334 (.Y(inst_cellmath__48_out0[12]), .A(N348), .B(N554));
NOR2XL inst_cellmath__48_I335 (.Y(inst_cellmath__48_out0[13]), .A(N349), .B(N554));
NOR2XL inst_cellmath__48_I336 (.Y(inst_cellmath__48_out0[14]), .A(N350), .B(N554));
NOR2XL inst_cellmath__48_I337 (.Y(inst_cellmath__48_out0[15]), .A(N352), .B(N553));
NOR2XL inst_cellmath__48_I338 (.Y(inst_cellmath__48_out0[16]), .A(N354), .B(N553));
NOR2XL inst_cellmath__48_I339 (.Y(inst_cellmath__48_out0[17]), .A(N356), .B(N553));
NOR2XL inst_cellmath__48_I340 (.Y(inst_cellmath__48_out0[18]), .A(N358), .B(N553));
NOR2XL inst_cellmath__48_I341 (.Y(inst_cellmath__48_out0[19]), .A(N360), .B(N553));
NOR2XL inst_cellmath__48_I342 (.Y(inst_cellmath__48_out0[20]), .A(N362), .B(N552));
NOR2XL inst_cellmath__48_I343 (.Y(inst_cellmath__48_out0[21]), .A(N364), .B(N552));
NOR2XL inst_cellmath__48_I344 (.Y(inst_cellmath__48_out0[22]), .A(N366), .B(N552));
NOR2X4 inst_cellmath__48_I345 (.Y(inst_cellmath__48_out0[23]), .A(N368), .B(N552));
NOR2XL inst_cellmath__48_I346 (.Y(inst_cellmath__48_out0[24]), .A(N370), .B(N552));
endmodule

module cynw_cm_float_cos_inst_cellmath__58__24__bdw1157874770_bdw (
	inst_cellmath__58__24__out0,
	inst_cellmath__58__24__in0
	); /* architecture "gate_level" */ 
output [1:0] inst_cellmath__58__24__out0;
input [24:23] inst_cellmath__58__24__in0;
INVX3 inst_cellmath__58__24__I15 (.Y(inst_cellmath__58__24__out0[0]), .A(inst_cellmath__58__24__in0[23]));
XOR2XL inst_cellmath__58__24__I16 (.Y(inst_cellmath__58__24__out0[1]), .A(inst_cellmath__58__24__in0[24]), .B(inst_cellmath__58__24__in0[23]));
endmodule

module cynw_cm_float_cos_inst_cellmath__61_0_bdw1157874770_bdw (
	inst_cellmath__61_0_out0,
	inst_cellmath__61_0_in0,
	inst_cellmath__61_0_in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__61_0_out0;
input [0:0] inst_cellmath__61_0_in0;
input [22:0] inst_cellmath__61_0_in1;
wire N95,N102,N104,N143,N145,N146,N147 
	,N148;
INVXL inst_cellmath__61_0_I46 (.Y(N95), .A(inst_cellmath__61_0_in1[0]));
INVX1 inst_cellmath__61_0_I53 (.Y(N102), .A(inst_cellmath__61_0_in1[7]));
INVXL inst_cellmath__61_0_I55 (.Y(N104), .A(inst_cellmath__61_0_in1[9]));
CLKINVX4 inst_cellmath__61_0_I93 (.Y(N143), .A(inst_cellmath__61_0_in0[0]));
INVX1 inst_cellmath__61_0_I98 (.Y(N148), .A(N143));
INVX2 inst_cellmath__61_0_I97 (.Y(N147), .A(N143));
CLKINVX4 inst_cellmath__61_0_I96 (.Y(N146), .A(N143));
INVX2 inst_cellmath__61_0_I95 (.Y(N145), .A(N143));
MXI2XL inst_cellmath__61_0_I69 (.Y(inst_cellmath__61_0_out0[0]), .A(N95), .B(inst_cellmath__61_0_in1[0]), .S0(N148));
XOR2XL inst_cellmath__61_0_I412 (.Y(inst_cellmath__61_0_out0[1]), .A(inst_cellmath__61_0_in1[1]), .B(N148));
CLKXOR2X1 inst_cellmath__61_0_I413 (.Y(inst_cellmath__61_0_out0[2]), .A(inst_cellmath__61_0_in1[2]), .B(N148));
XOR2XL inst_cellmath__61_0_I414 (.Y(inst_cellmath__61_0_out0[3]), .A(inst_cellmath__61_0_in1[3]), .B(N147));
XOR2XL inst_cellmath__61_0_I415 (.Y(inst_cellmath__61_0_out0[4]), .A(inst_cellmath__61_0_in1[4]), .B(N147));
CLKXOR2X1 inst_cellmath__61_0_I416 (.Y(inst_cellmath__61_0_out0[5]), .A(inst_cellmath__61_0_in1[5]), .B(N147));
XOR2XL inst_cellmath__61_0_I417 (.Y(inst_cellmath__61_0_out0[6]), .A(inst_cellmath__61_0_in1[6]), .B(N147));
MXI2X1 inst_cellmath__61_0_I76 (.Y(inst_cellmath__61_0_out0[7]), .A(N102), .B(inst_cellmath__61_0_in1[7]), .S0(N147));
CLKXOR2X1 inst_cellmath__61_0_I419 (.Y(inst_cellmath__61_0_out0[8]), .A(inst_cellmath__61_0_in1[8]), .B(N146));
MXI2X1 inst_cellmath__61_0_I78 (.Y(inst_cellmath__61_0_out0[9]), .A(N104), .B(inst_cellmath__61_0_in1[9]), .S0(N146));
XOR2XL inst_cellmath__61_0_I421 (.Y(inst_cellmath__61_0_out0[10]), .A(inst_cellmath__61_0_in1[10]), .B(N146));
XOR2XL inst_cellmath__61_0_I422 (.Y(inst_cellmath__61_0_out0[11]), .A(inst_cellmath__61_0_in1[11]), .B(N146));
XOR2XL inst_cellmath__61_0_I423 (.Y(inst_cellmath__61_0_out0[12]), .A(inst_cellmath__61_0_in1[12]), .B(N146));
XOR2XL inst_cellmath__61_0_I424 (.Y(inst_cellmath__61_0_out0[13]), .A(inst_cellmath__61_0_in1[13]), .B(N145));
XOR2XL inst_cellmath__61_0_I425 (.Y(inst_cellmath__61_0_out0[14]), .A(inst_cellmath__61_0_in1[14]), .B(N145));
XOR2XL inst_cellmath__61_0_I426 (.Y(inst_cellmath__61_0_out0[15]), .A(inst_cellmath__61_0_in1[15]), .B(N145));
XOR2XL inst_cellmath__61_0_I427 (.Y(inst_cellmath__61_0_out0[16]), .A(inst_cellmath__61_0_in1[16]), .B(N145));
XOR2XL inst_cellmath__61_0_I428 (.Y(inst_cellmath__61_0_out0[17]), .A(inst_cellmath__61_0_in1[17]), .B(N145));
XOR2XL inst_cellmath__61_0_I429 (.Y(inst_cellmath__61_0_out0[18]), .A(inst_cellmath__61_0_in1[18]), .B(N146));
XOR2XL inst_cellmath__61_0_I430 (.Y(inst_cellmath__61_0_out0[19]), .A(inst_cellmath__61_0_in1[19]), .B(N146));
XOR2XL inst_cellmath__61_0_I431 (.Y(inst_cellmath__61_0_out0[20]), .A(inst_cellmath__61_0_in1[20]), .B(N146));
XOR2XL inst_cellmath__61_0_I432 (.Y(inst_cellmath__61_0_out0[21]), .A(inst_cellmath__61_0_in1[21]), .B(N146));
XOR2XL inst_cellmath__61_0_I433 (.Y(inst_cellmath__61_0_out0[22]), .A(inst_cellmath__61_0_in1[22]), .B(N146));
endmodule

module cynw_cm_float_cos_inst_cellmath__195__80__2WWMM_2WWMM_bdw1157874770_bdw (
	inst_cellmath__195__80__2WWMM_2WWMM_out0,
	inst_cellmath__195__80__2WWMM_2WWMM_in0
	); /* architecture "gate_level" */ 
output [72:0] inst_cellmath__195__80__2WWMM_2WWMM_out0;
input [22:17] inst_cellmath__195__80__2WWMM_2WWMM_in0;
wire N82,N85,N88,N89,N92,N93,N95 
	,N96,N98,N102,N104,N107,N108,N110,N111 
	,N112,N113,N114,N115,N117,N118,N119,N121 
	,N122,N123,N126,N128,N129,N131,N132,N134 
	,N135,N136,N137,N138,N140,N141,N142,N143 
	,N144,N145,N146,N147,N149,N150,N151,N152 
	,N153,N154,N155,N156,N159,N160,N161,N162 
	,N163,N164,N165,N167,N168,N170,N173,N174 
	,N4260,N4261,N4263,N4264,N4265,N4272,N4273,N4274 
	,N4275,N4276,N4278,N4279,N4280,N4281,N4282,N4283 
	,N4290,N4291,N4292,N4297,N4299,N4300,N4303,N4304 
	,N4305,N4307,N4309,N4311,N4312,N4323,N4325,N4326 
	,N4327,N4329,N4330,N4332,N4333,N4334,N4335,N4337 
	,N4339,N4340,N4348,N4349,N4350,N4351,N4352,N4353 
	,N4355,N4356,N4357,N4358,N4364,N4365,N4367,N4368 
	,N4369,N4371,N4373,N4374,N4375,N4389,N4397,N4399 
	,N4402,N4403,N4404,N4405,N4418,N4419,N4421,N4424 
	,N4425,N4427,N4429,N4430,N4431,N4432,N4439,N4440 
	,N4441,N4442,N4444,N4445,N4451,N4455,N4456,N4457 
	,N4458,N4459,N4460,N4461,N4465,N4466,N4467,N4479 
	,N4480,N4481,N4482,N4483,N4484,N4490,N4491,N4492 
	,N4493,N4497,N4498,N4499,N4500,N4501,N4508,N4509 
	,N4510,N4511,N4513,N4514,N4515,N4518,N4520,N4522 
	,N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4533 
	,N4534,N4538,N4542,N4545,N4546,N4547,N4549,N4553 
	,N4554,N4555,N4556,N4557,N4559,N4561,N4563,N4566 
	,N4567,N4577,N4579,N4580,N4581,N4582,N4585,N4587 
	,N4588,N4589,N4590,N4592,N4594,N4598,N4599,N4600 
	,N4612,N4613,N4614,N4616,N4617,N4618,N4622,N4625 
	,N4627,N4628,N4630,N4631,N4633,N4635,N4636,N4637 
	,N4638,N4648,N4649,N4655,N4657,N4662,N4663,N4665 
	,N4666,N4667,N4669,N4671,N4672,N4673,N4685,N4692 
	,N4693,N4699,N4700,N4701,N4702,N4704,N4705,N4707 
	,N4709,N4710,N4717,N4718,N4721,N4722,N4723,N4724 
	,N4725,N4726,N4727,N4728,N4732,N4733,N4734,N4735 
	,N4738,N4739,N4742,N4743,N4755,N4758,N4760,N4761 
	,N4763,N4764,N4767,N4769,N4771,N4778,N4780,N4781 
	,N4782,N4783,N4784,N4785,N4786,N4794,N4795,N4796 
	,N4797,N4798,N4799,N4801,N4802,N4803,N4806,N4807 
	,N4808,N4820,N4821,N4823,N4829,N4831,N4832,N4833 
	,N4834,N4836,N4837,N4838,N4839,N4841,N4854,N4855 
	,N4858,N4859,N4861,N4863,N4867,N4868,N4870,N4871 
	,N4872,N4886,N4888,N4891,N4892,N4893,N4894,N4896 
	,N4909,N4910,N4912,N4914,N4916,N4918,N4919,N4921 
	,N4922,N4923,N4934,N4936,N4939,N4942,N4943,N4945 
	,N4947,N4949,N4950,N4976,N4978,N4979,N4982,N4988 
	,N4989,N4991,N4992,N4994,N4995,N4997,N4998,N5007 
	,N5008,N5009,N5010,N5011,N5012,N5013,N5020,N5021 
	,N5023,N5024,N5025,N5026,N5039,N5040,N5042,N5043 
	,N5047,N5048,N5049,N5050,N5051,N5053,N5054,N5055 
	,N5056,N5067,N5071,N5073,N5075,N5076,N5080,N5081 
	,N5084,N5085,N5087,N5098,N5102,N5105,N5106,N5108 
	,N5109,N5115,N5116,N5117,N5120,N5121,N5123,N5126 
	,N5127,N5128,N5135,N5142,N5143,N5148,N5151,N5152 
	,N5153,N5155,N5156,N5157,N5174,N5175,N5181,N5186 
	,N5188,N5189,N5209,N5210,N5213,N5215,N5216,N5219 
	,N5220,N5221,N5222,N5223,N5225,N5226,N5235,N5241 
	,N5247,N5248,N5249,N5250,N5253,N5255,N5257,N5258 
	,N5265,N5268,N5269,N5270,N5272,N5276,N5280,N5281 
	,N5282,N5284,N5287,N5288,N5289,N5290,N5296,N5297 
	,N5298,N5302,N5305,N5308,N5314,N5315,N5316,N5319 
	,N5320,N5321,N5322,N5329,N5331,N5332,N5337,N5340 
	,N5341,N5346,N5349,N5350,N5351,N5353,N5354,N5356 
	,N5357,N5364,N5365,N5366,N5368,N5369,N5371,N5373 
	,N5375,N5376,N5377,N5378,N5379,N5380,N5382,N5383 
	,N5385,N5386,N5387,N5394,N5397,N5398,N5402,N5403 
	,N5408,N5409,N5410,N5412,N5414,N5416,N5417,N5418 
	,N5426,N5427,N5429,N5431,N5437,N5443,N5444,N5447 
	,N5448,N5451,N5452,N5455,N5456,N5466,N5469,N5474 
	,N5477,N5478,N5480,N5482,N5483,N5484,N5486,N5498 
	,N5500,N5501,N5504,N5505,N5506,N5509,N5510,N5512 
	,N5522,N5526,N5529,N5533,N5535,N5536,N5538,N5539 
	,N5540,N5541,N5543,N5544,N5545,N5546,N5555,N5565 
	,N5567,N5569,N5571,N5573,N5574,N5576,N5578,N5589 
	,N5596,N5598,N5599,N5601,N5604,N5605,N5606,N5614 
	,N5620,N5628,N5629,N5632,N5633,N5634,N5636,N5637 
	,N5655,N5658,N5661,N5662,N5663,N5664,N5666,N5668 
	,N5669,N5671,N5672,N5673,N5674,N5687,N5691,N5693 
	,N5698,N5700,N5702,N5707,N5708,N5710,N5711,N5721 
	,N5722,N5732,N5733,N5734,N5735,N5737,N5738,N5740 
	,N5741,N5742,N5744,N5745,N5754,N5759,N5763,N5767 
	,N5769,N5770,N5772,N5774,N5777,N5778,N5788,N5789 
	,N5790,N5792,N5794,N5795,N5798,N5799,N5800,N5801 
	,N5802,N5803,N5804,N5818,N5830,N5832,N5833,N5834 
	,N5836,N5837,N5838,N5839,N5841,N5842,N5843,N5851 
	,N5855,N5861,N5862,N5863,N5864,N5866,N5867,N5868 
	,N5871,N5874,N5875,N5888,N5890,N5895,N5900,N5901 
	,N5902,N5904,N5905,N5908,N5910,N5911,N5921,N5923 
	,N5924,N5925,N5927,N5930,N5933,N5935,N5936,N5937 
	,N5938,N5939,N5941,N5943,N5956,N5959,N5965,N5966 
	,N5967,N5971,N5973,N5974,N5975,N5976,N5986,N5989 
	,N5990,N5994,N5996,N5998,N5999,N6000,N6001,N6002 
	,N6014,N6020,N6027,N6028,N6029,N6030,N6033,N6034 
	,N6037,N6038,N6039,N6040,N6050,N6061,N6064,N6066 
	,N6067,N6073,N6075,N6076,N6077,N6082,N6083,N6089 
	,N6093,N6097,N6098,N6099,N6100,N6101,N6102,N6105 
	,N6108,N6109,N6111,N6117,N6120,N6127,N6129,N6131 
	,N6136,N6138,N6139,N6142,N6144,N6146,N6156,N6159 
	,N6162,N6166,N6171,N6173,N6174,N6175,N6176,N6177 
	,N6178,N6179,N6180,N6196,N6202,N6204,N6205,N6206 
	,N6208,N6209,N6210,N6227,N6231,N6232,N6233,N6237 
	,N6238,N6240,N6243,N6252,N6254,N6257,N6261,N6264 
	,N6266,N6267,N6271,N6272,N6273,N6275,N6276,N6277 
	,N6287,N6293,N6294,N6296,N6299,N6301,N6302,N6303 
	,N6304,N6306,N6307,N6308,N6309,N6310,N6311,N6330 
	,N6336,N6340,N6341,N6344,N6345,N6346,N6349,N6350 
	,N6356,N6360,N6365,N6366,N6367,N6368,N6370,N6373 
	,N6374,N6377,N6378,N6379,N6380,N6381,N6383,N6389 
	,N6391,N6395,N6397,N6400,N6403,N6404,N6406,N6407 
	,N6409,N6411,N6412,N6413,N6414,N6415,N6417,N6418 
	,N6419,N6424,N6442,N6446,N6448,N6449,N6453,N6454 
	,N6455,N6457,N6458,N6459,N6477,N6479,N6480,N6482 
	,N6483,N6484,N6485,N6487,N6488,N6490,N6502,N6511 
	,N6512,N6513,N6516,N6519,N6521,N6522,N6536,N6542 
	,N6543,N6545,N6546,N6547,N6548,N6550,N6553,N6554 
	,N6565,N6567,N6571,N6573,N6578,N6579,N6581,N6583 
	,N6585,N6586,N6587,N6594,N6605,N6606,N6608,N6609 
	,N6611,N6615,N6623,N6627,N6635,N6643,N6647,N6651 
	,N6653,N6655,N6659,N6667,N6671,N6675,N6677,N6679 
	,N6681,N6683,N6685,N6687,N6695,N6697,N6701,N6703 
	,N6705,N6707,N6709,N6711,N6715,N6717,N6721,N6725 
	,N6727,N6729,N6733,N6735,N6737,N6741,N6745,N6747 
	,N6749,N6751,N6753,N6755,N6757,N6759,N6765,N6767 
	,N6769,N6771,N6773,N6775,N6777,N6779,N6781,N6783 
	,N6785,N6787,N6789,N6791,N6793,N6795,N6797,N7996 
	,N7997,N7998,N7999,N8000,N8001,N8004,N8005,N8006 
	,N8007,N8010,N8011,N8012,N8015,N8016,N8017,N8018 
	,N8019,N8020,N8023,N8024,N8025,N8028,N8029,N8030 
	,N8031,N8032,N8033,N8034,N8035,N8036,N8039,N8040 
	,N8041,N8044,N8045,N8046,N8054,N8055,N8056,N8059 
	,N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067 
	,N8070,N8071,N8072,N8075,N8076,N8077,N8080,N8081 
	,N8086,N8087,N8096,N8097,N8098,N8099,N8107,N8109 
	,N8113,N8114,N8115,N8118,N8119,N8120,N8121,N8122 
	,N8123,N8128,N8129,N8130,N8131,N8132,N8133,N8134 
	,N8135,N8136,N8137,N8143,N8144,N8147,N8150,N8151 
	,N8152,N8153,N8156,N8160,N8161,N8162,N8165,N8168 
	,N8171,N8172,N8175,N8176,N8179,N8183,N8184,N8185 
	,N8190,N8193,N8194,N8196,N8197,N8198,N8201,N8202 
	,N8203,N8206,N8207,N8212,N8213,N8215,N8216,N8217 
	,N8220,N8222,N8223,N8224,N8227,N8230,N8231,N8234 
	,N8235,N8236,N8237,N8238,N8243,N8244,N8245,N8248 
	,N8251,N8252,N8253,N8256,N8257,N8258,N8260,N8261 
	,N8262,N8265,N8266,N8270,N8279,N8280,N8287,N8288 
	,N8290,N8313,N8323,N8330,N8337,N8344,N8351,N8358 
	,N8365,N8372,N8379,N8388,N8396,N8404,N8412,N8420 
	,N8428,N8436,N8444,N8452,N8460,N8468,N8476,N8484 
	,N8492,N8500,N8508,N8516,N8524,N8532,N8540,N11162 
	;
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5316 (.Y(N7996), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5317 (.Y(N7997), .A(N7996));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5318 (.Y(N7998), .A(N7997));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1 (.Y(N82), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8609 (.Y(N7999), .A(N7998), .B(N82));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5321 (.Y(N8001), .A(N7999));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5320 (.Y(N8000), .A(N7999));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5324 (.Y(N8004), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4 (.Y(N85), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I8610 (.Y(N8005), .A(N85), .B(N8004));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5327 (.Y(N8007), .A(N8005));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5326 (.Y(N8006), .A(N8005));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I6 (.Y(N6623), .A(N8007), .B(N8001));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I7 (.Y(N88), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8 (.Y(N89), .A(N88), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8611 (.Y(N8010), .A(N8004), .B(N89));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5332 (.Y(N8012), .A(N8010));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5331 (.Y(N8011), .A(N8010));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10 (.Y(N6627), .A(N8012), .B(N8001));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I11 (.Y(N92), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I12 (.Y(N93), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B(N92));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8612 (.Y(N8015), .A(N8004), .B(N93));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5337 (.Y(N8017), .A(N8015));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5336 (.Y(N8016), .A(N8015));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I14 (.Y(N95), .A(N8017), .B(N8000));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I15 (.Y(N96), .A(N88), .B(N92));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8613 (.Y(N8018), .A(N8004), .B(N96));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5340 (.Y(N8020), .A(N8018));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5339 (.Y(N8019), .A(N8018));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I17 (.Y(N98), .A(N8020), .B(N8000));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5871 (.Y(N8023), .A(N85), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5345 (.Y(N8025), .A(N8023));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5344 (.Y(N8024), .A(N8023));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I19 (.Y(N6635), .A(N8025), .B(N8000));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5824 (.Y(N8028), .A(N89), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5350 (.Y(N8030), .A(N8028));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5349 (.Y(N8029), .A(N8028));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I21 (.Y(N102), .A(N8030), .B(N8000));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5825 (.Y(N8031), .A(N93), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5353 (.Y(N8033), .A(N8031));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5352 (.Y(N8032), .A(N8031));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I23 (.Y(N104), .A(N8033), .B(N8000));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8614 (.Y(N8034), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]), .B(N96));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5356 (.Y(N8036), .A(N8034));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5355 (.Y(N8035), .A(N8034));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I25 (.Y(N6643), .A(N8036), .B(N8000));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I26 (.Y(N107), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I27 (.Y(N108), .A(N107), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8615 (.Y(N8039), .A(N7998), .B(N108));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5361 (.Y(N8041), .A(N8039));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5360 (.Y(N8040), .A(N8039));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I29 (.Y(N110), .A(N8007), .B(N8041));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I30 (.Y(N111), .A(N8012), .B(N8041));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I31 (.Y(N112), .A(N8017), .B(N8041));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I32 (.Y(N113), .A(N8020), .B(N8040));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I33 (.Y(N114), .A(N8025), .B(N8040));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I34 (.Y(N115), .A(N8030), .B(N8040));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I35 (.Y(N6647), .A(N8033), .B(N8040));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I36 (.Y(N117), .A(N8036), .B(N8040));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I37 (.Y(N118), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I38 (.Y(N119), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]), .B(N118));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I8616 (.Y(N8044), .A(N119), .B(N7998));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5366 (.Y(N8046), .A(N8044));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5365 (.Y(N8045), .A(N8044));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I40 (.Y(N121), .A(N8007), .B(N8046));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I41 (.Y(N122), .A(N8012), .B(N8046));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I42 (.Y(N123), .A(N8016), .B(N8045));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I43 (.Y(N6651), .A(N8020), .B(N8045));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I44 (.Y(N6653), .A(N8025), .B(N8045));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I45 (.Y(N126), .A(N8030), .B(N8045));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I46 (.Y(N6655), .A(N8033), .B(N8045));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I47 (.Y(N128), .A(N8036), .B(N8045));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I48 (.Y(N129), .A(N107), .B(N118));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8617 (.Y(N8054), .A(N7998), .B(N129));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5376 (.Y(N8056), .A(N8054));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5375 (.Y(N8055), .A(N8054));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I50 (.Y(N131), .A(N8006), .B(N8056));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I51 (.Y(N132), .A(N8011), .B(N8056));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I52 (.Y(N6659), .A(N8016), .B(N8056));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I53 (.Y(N134), .A(N8019), .B(N8055));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I54 (.Y(N135), .A(N8025), .B(N8055));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I55 (.Y(N136), .A(N8029), .B(N8055));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I56 (.Y(N137), .A(N8033), .B(N8055));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I57 (.Y(N138), .A(N8035), .B(N8055));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I8618 (.Y(N8059), .A(N82), .B(N7997));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5381 (.Y(N8061), .A(N8059));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5380 (.Y(N8060), .A(N8059));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I59 (.Y(N140), .A(N8006), .B(N8061));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I60 (.Y(N141), .A(N8011), .B(N8061));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I61 (.Y(N142), .A(N8016), .B(N8061));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I62 (.Y(N143), .A(N8019), .B(N8060));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I63 (.Y(N144), .A(N8024), .B(N8060));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I64 (.Y(N145), .A(N8029), .B(N8060));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I65 (.Y(N146), .A(N8032), .B(N8060));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I66 (.Y(N147), .A(N8035), .B(N8060));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5832 (.Y(N8062), .A(N108), .B(N7997));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5384 (.Y(N8064), .A(N8062));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5383 (.Y(N8063), .A(N8062));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I68 (.Y(N149), .A(N8006), .B(N8064));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I69 (.Y(N150), .A(N8011), .B(N8064));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I70 (.Y(N151), .A(N8016), .B(N8064));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I71 (.Y(N152), .A(N8019), .B(N8063));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I72 (.Y(N153), .A(N8024), .B(N8063));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I73 (.Y(N154), .A(N8029), .B(N8063));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I74 (.Y(N155), .A(N8032), .B(N8063));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I75 (.Y(N156), .A(N8035), .B(N8063));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I8619 (.Y(N8065), .A(N119), .B(N7997));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5387 (.Y(N8067), .A(N8065));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5386 (.Y(N8066), .A(N8065));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I77 (.Y(N6667), .A(N8006), .B(N8067));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I78 (.Y(N159), .A(N8011), .B(N8067));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I79 (.Y(N160), .A(N8016), .B(N8067));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I80 (.Y(N161), .A(N8019), .B(N8066));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I81 (.Y(N162), .A(N8024), .B(N8066));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I82 (.Y(N163), .A(N8029), .B(N8066));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I83 (.Y(N164), .A(N8032), .B(N8066));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I84 (.Y(N165), .A(N8035), .B(N8066));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I8620 (.Y(N8070), .A(N129), .B(N7997));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5392 (.Y(N8072), .A(N8070));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5391 (.Y(N8071), .A(N8070));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I86 (.Y(N167), .A(N8006), .B(N8072));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I87 (.Y(N168), .A(N8011), .B(N8072));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I88 (.Y(N6671), .A(N8016), .B(N8072));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I89 (.Y(N170), .A(N8019), .B(N8071));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I5835 (.Y(N8075), .A(N8024), .B(N8071));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5397 (.Y(N8077), .A(N8075));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5396 (.Y(N8076), .A(N8075));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I91 (.Y(N6675), .A(N8029), .B(N8071));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I92 (.Y(N173), .A(N8032), .B(N8071));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I93 (.Y(N174), .A(N8035), .B(N8071));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5400 (.Y(N8080), .A(N6623));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5401 (.Y(N8081), .A(N6627));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I106 (.Y(N6677), .A(N6627), .B(N6623));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5406 (.Y(N8086), .A(N95));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5407 (.Y(N8087), .A(N98));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I190 (.Y(N6679), .A(N98), .B(N95));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I249 (.Y(N6681), .A(N102), .B(N6635));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5416 (.Y(N8096), .A(N102));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5417 (.Y(N8097), .A(N6635));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5418 (.Y(N8098), .A(N104));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5419 (.Y(N8099), .A(N6643));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I329 (.Y(N6683), .A(N6643), .B(N104));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I401 (.Y(N6685), .A(N111), .B(N110));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5427 (.Y(N8107), .A(N110));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5429 (.Y(N8109), .A(N111));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I477 (.Y(N6687), .A(N113), .B(N112));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5433 (.Y(N8113), .A(N113));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5434 (.Y(N8114), .A(N112));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5435 (.Y(N8115), .A(N115));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5439 (.Y(N8119), .A(N114));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5438 (.Y(N8118), .A(N114));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8621 (.Y(N8120), .A(N115), .B(N114));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5443 (.Y(N8123), .A(N8120));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5442 (.Y(N8122), .A(N8120));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5441 (.Y(N8121), .A(N8120));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5448 (.Y(N8128), .A(N6647));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8622 (.Y(N8129), .A(N117), .B(N6647));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5452 (.Y(N8132), .A(N8129));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5451 (.Y(N8131), .A(N8129));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5450 (.Y(N8130), .A(N8129));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5453 (.Y(N8133), .A(N117));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5454 (.Y(N8134), .A(N121));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8623 (.Y(N8135), .A(N122), .B(N121));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5457 (.Y(N8137), .A(N8135));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5456 (.Y(N8136), .A(N8135));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5463 (.Y(N8143), .A(N122));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5464 (.Y(N8144), .A(N6651));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I783 (.Y(N6695), .A(N6651), .B(N123));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5467 (.Y(N8147), .A(N123));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I857 (.Y(N6697), .A(N126), .B(N6653));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5470 (.Y(N8150), .A(N6653));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5471 (.Y(N8151), .A(N126));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5472 (.Y(N8152), .A(N128));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5473 (.Y(N8153), .A(N6655));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8624 (.Y(N8156), .A(N128), .B(N6655));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5481 (.Y(N8161), .A(N132));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5480 (.Y(N8160), .A(N132));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5482 (.Y(N8162), .A(N131));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1011 (.Y(N6701), .A(N132), .B(N131));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5485 (.Y(N8165), .A(N134));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1087 (.Y(N6703), .A(N134), .B(N6659));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5488 (.Y(N8168), .A(N6659));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1162 (.Y(N6705), .A(N136), .B(N135));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5491 (.Y(N8171), .A(N136));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5492 (.Y(N8172), .A(N135));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1237 (.Y(N6707), .A(N138), .B(N137));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5495 (.Y(N8175), .A(N137));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5496 (.Y(N8176), .A(N138));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1313 (.Y(N6709), .A(N141), .B(N140));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5499 (.Y(N8179), .A(N140));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5504 (.Y(N8184), .A(N141));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5503 (.Y(N8183), .A(N141));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5505 (.Y(N8185), .A(N143));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5510 (.Y(N8190), .A(N142));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1396 (.Y(N6711), .A(N143), .B(N142));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5513 (.Y(N8193), .A(N144));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8625 (.Y(N8194), .A(N145), .B(N144));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5517 (.Y(N8197), .A(N8194));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5516 (.Y(N8196), .A(N8194));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5518 (.Y(N8198), .A(N145));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1542 (.Y(N6715), .A(N147), .B(N146));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5521 (.Y(N8201), .A(N147));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5522 (.Y(N8202), .A(N146));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5523 (.Y(N8203), .A(N149));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1618 (.Y(N6717), .A(N150), .B(N149));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5526 (.Y(N8206), .A(N150));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5527 (.Y(N8207), .A(N152));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5533 (.Y(N8213), .A(N151));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5532 (.Y(N8212), .A(N151));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I5843 (.Y(N8215), .A(N152), .B(N151));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5536 (.Y(N8216), .A(N153));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5537 (.Y(N8217), .A(N154));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1771 (.Y(N6721), .A(N154), .B(N153));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5540 (.Y(N8220), .A(N156));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I5739 (.Y(N8222), .A(N156), .B(N155));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5543 (.Y(N8223), .A(N155));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5544 (.Y(N8224), .A(N159));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1922 (.Y(N6725), .A(N159), .B(N6667));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5547 (.Y(N8227), .A(N6667));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1997 (.Y(N6727), .A(N161), .B(N160));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5550 (.Y(N8230), .A(N161));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5551 (.Y(N8231), .A(N160));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2074 (.Y(N6729), .A(N163), .B(N162));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5554 (.Y(N8234), .A(N162));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5555 (.Y(N8235), .A(N163));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I8626 (.Y(N8236), .A(N165), .B(N164));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5558 (.Y(N8238), .A(N8236));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5557 (.Y(N8237), .A(N8236));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5563 (.Y(N8243), .A(N165));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5564 (.Y(N8244), .A(N164));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5565 (.Y(N8245), .A(N167));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2227 (.Y(N6733), .A(N168), .B(N167));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5568 (.Y(N8248), .A(N168));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2301 (.Y(N6735), .A(N170), .B(N6671));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5571 (.Y(N8251), .A(N6671));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5572 (.Y(N8252), .A(N170));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5573 (.Y(N8253), .A(N6675));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2379 (.Y(N6737), .A(N6675), .B(N8077));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5576 (.Y(N8256), .A(N8077));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5577 (.Y(N8257), .A(N174));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I5845 (.Y(N8258), .A(N174), .B(N173));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5581 (.Y(N8261), .A(N8258));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5580 (.Y(N8260), .A(N8258));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5582 (.Y(N8262), .A(N173));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2531 (.Y(N4976), .A(N8193), .B(N8134));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2533 (.Y(N4260), .A(N8203), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2534 (.Y(N4261), .A(N8161), .B(N6697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2535 (.Y(N6741), .A(N6681), .B(N6709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2536 (.Y(N4263), .A(N8185), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2537 (.Y(N4264), .A(N8152), .B(N8086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2538 (.Y(N4265), .A(N6685), .B(N8128));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2540 (.Y(N4278), .A(N8080), .B(N8165));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2541 (.Y(N5668), .A(N6687), .B(N8237));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2542 (.Y(N4276), .A(N6707), .B(N6735));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2544 (.Y(N4281), .A(N6727), .B(N4976));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5217 (.Y(N4272), .A(N8253), .B(N8216), .C(N4260));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2546 (.Y(N4273), .A(N4261), .B(N4263));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2547 (.Y(N4274), .A(N4264), .B(N6741));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2548 (.Y(N4275), .A(N4265), .B(N5668));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2552 (.Y(N4279), .A(N4278), .B(N4273));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2553 (.Y(N4280), .A(N4274), .B(N4275));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2555 (.Y(N4282), .A(N4281), .B(N4280));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4960 (.Y(N4283), .A(N4276), .B(N4272), .C(N4279));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2557 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[0]), .A(N4282), .B(N4283));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2563 (.Y(N4290), .A(N8179), .B(N8134));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2564 (.Y(N4291), .A(N8162), .B(N8245));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2565 (.Y(N4292), .A(N8150), .B(N8253));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5683 (.Y(N8265), .A(N6705), .B(N6729));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5586 (.Y(N8266), .A(N8265));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2569 (.Y(N6745), .A(N8152), .B(N6725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2570 (.Y(N4297), .A(N8087), .B(N6717));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2571 (.Y(N5383), .A(N8144), .B(N8165));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2572 (.Y(N4299), .A(N8132));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2573 (.Y(N4300), .A(N4299), .B(N4291));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5590 (.Y(N8270), .A(N6715));
NAND2XL hyperpropagate_3_1_A_I5947 (.Y(N8323), .A(N8107), .B(N8217));
NOR2XL hyperpropagate_3_1_A_I5948 (.Y(N4303), .A(N8270), .B(N8323));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2577 (.Y(N4304), .A(N4290), .B(N4292));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2578 (.Y(N4305), .A(N4297), .B(N8266));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2580 (.Y(N4307), .A(N5383), .B(N4276));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2582 (.Y(N4309), .A(N4300), .B(N4303));
NAND3XL hyperpropagate_4_1_A_I8635 (.Y(N11162), .A(N8207), .B(N4307), .C(N8098));
NOR2XL hyperpropagate_4_1_A_I8636 (.Y(N4312), .A(N6745), .B(N11162));
NAND2XL hyperpropagate_3_1_A_I5949 (.Y(N8330), .A(N4304), .B(N4305));
NOR2XL hyperpropagate_3_1_A_I5950 (.Y(N4311), .A(N4309), .B(N8330));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2586 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[1]), .A(N4312), .B(N4311));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2593 (.Y(N6747), .A(N6705), .B(N6697));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5854 (.Y(N6749), .AN(N8135), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2595 (.Y(N4323), .A(N8185), .B(N8113));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2596 (.Y(N6751), .A(N6721), .B(N8197));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2597 (.Y(N4325), .A(N8243), .B(N8087));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2598 (.Y(N4326), .A(N6685), .B(N6701));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2599 (.Y(N4327), .A(N6717), .B(N8175));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2600 (.Y(N6101), .A(N8213), .B(N8099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2601 (.Y(N4329), .A(N8201), .B(N6735));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2602 (.Y(N4330), .A(N6695), .B(N6703));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2604 (.Y(N4332), .A(N6749), .B(N6751));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2605 (.Y(N4333), .A(N4325), .B(N4323));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2606 (.Y(N4334), .A(N6747), .B(N4326));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2607 (.Y(N4335), .A(N4327), .B(N4330));
NAND2XL hyperpropagate_3_1_A_I5951 (.Y(N8337), .A(N6737), .B(N6101));
NOR2XL hyperpropagate_3_1_A_I5952 (.Y(N4337), .A(N4329), .B(N8337));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2611 (.Y(N4339), .A(N4334), .B(N4335));
NAND2XL hyperpropagate_3_1_A_I5953 (.Y(N8344), .A(N4332), .B(N4333));
NOR2XL hyperpropagate_3_1_A_I5954 (.Y(N4340), .A(N4339), .B(N8344));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2613 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[2]), .A(N4337), .B(N4340));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2619 (.Y(N4348), .A(N8253), .B(N8171));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2620 (.Y(N4349), .A(N8151), .B(N8143));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2621 (.Y(N4350), .A(N8096), .B(N8184));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2622 (.Y(N4351), .A(N8217), .B(N8198));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2623 (.Y(N4352), .A(N8224), .B(N8161));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2624 (.Y(N4353), .A(N6729), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2625 (.Y(N6753), .A(N8152), .B(N8243));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2626 (.Y(N4355), .A(N8190), .B(N8257));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2627 (.Y(N4356), .A(N8220), .B(N8201));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2628 (.Y(N4357), .A(N8128), .B(N6687));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2629 (.Y(N4358), .A(N4349), .B(N4350));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5599 (.Y(N8279), .A(N6703));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4952 (.Y(N4367), .A(N6753), .B(N4351));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4950 (.Y(N4371), .A(N4367), .B(N4358));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2634 (.Y(N4368), .A(N4352), .B(N4355));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2635 (.Y(N4364), .A(N4348), .B(N4356));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2636 (.Y(N4365), .A(N4353), .B(N4357));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I4973 (.Y(N4369), .A(N8245), .B(N6735), .C(N4368));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2641 (.Y(N4373), .A(N4364), .B(N4365));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2643 (.Y(N4375), .A(N4371), .B(N8279));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2645 (.Y(N4374), .A(N4373), .B(N4369));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2647 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[3]), .A(N4375), .B(N4374));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2659 (.Y(N4389), .A(N8115), .B(N8151));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2664 (.Y(N4399), .A(N6701), .B(N8244));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5600 (.Y(N8280), .A(N6683));
NAND2XL hyperpropagate_3_1_A_I5955 (.Y(N8351), .A(N8172), .B(N8107));
NOR2XL hyperpropagate_3_1_A_I5956 (.Y(N4397), .A(N8280), .B(N8351));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4976 (.Y(N4405), .A(N6659), .B(N6635), .C(N4399));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5233 (.Y(N4403), .A(N8207), .B(N8251), .C(N6707), .D(N6721));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I4978 (.Y(N4402), .A(N4389), .B(N4260), .C(N4397));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2674 (.Y(N4404), .A(N4403), .B(N4402));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2676 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[4]), .A(N4405), .B(N4404));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5700 (.Y(N6755), .AN(N110), .B(N8119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2685 (.Y(N6232), .A(N8248), .B(N8234));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2686 (.Y(N6757), .A(N8096), .B(N8217));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2688 (.Y(N4418), .A(N8137), .B(N8185));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2689 (.Y(N4419), .A(N8244), .B(N8213));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2690 (.Y(N5053), .A(N8230), .B(N8251));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2691 (.Y(N4421), .A(N8128), .B(N8261));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2692 (.Y(N4427), .A(N6715), .B(N6695));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2694 (.Y(N4424), .A(N6757), .B(N5053));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2695 (.Y(N4425), .A(N4419), .B(N4418));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I4979 (.Y(N4430), .AN(N4421), .B(N8160), .C(N6705));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4980 (.Y(N4432), .A(N6232), .B(N6755), .C(N4427));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2699 (.Y(N4429), .A(N4424), .B(N4425));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2701 (.Y(N4431), .A(N4430), .B(N4429));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2703 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[5]), .A(N4432), .B(N4431));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2708 (.Y(N4439), .A(N8097), .B(N8245));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2709 (.Y(N4440), .A(N8172), .B(N8151));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2710 (.Y(N4441), .A(N8234), .B(N8184));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2711 (.Y(N4442), .A(N8217), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2712 (.Y(N6304), .A(N8206), .B(N8123));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2713 (.Y(N4444), .A(N8137), .B(N8114));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2714 (.Y(N4445), .A(N8202), .B(N8087));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2716 (.Y(N4799), .A(N8220), .B(N8212));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2717 (.Y(N6759), .A(N8176), .B(N8252));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2720 (.Y(N4451), .A(N8132), .B(N6683));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5607 (.Y(N8287), .A(N6695));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2723 (.Y(N4459), .A(N4441), .B(N4439));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2724 (.Y(N4455), .A(N6759), .B(N4440));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2725 (.Y(N4456), .A(N4355), .B(N4445));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2726 (.Y(N4457), .A(N4799), .B(N4442));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2727 (.Y(N4458), .A(N4444), .B(N4451));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2729 (.Y(N4460), .A(N4459), .B(N4278));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2730 (.Y(N4461), .A(N4455), .B(N4456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2731 (.Y(N4465), .A(N4457), .B(N4458));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4981 (.Y(N4467), .A(N6304), .B(N8287), .C(N4461));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2735 (.Y(N4466), .A(N4465), .B(N4460));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2737 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[6]), .A(N4467), .B(N4466));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2747 (.Y(N4479), .A(N8137), .B(N6709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2748 (.Y(N4480), .A(N8207), .B(N8196));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2749 (.Y(N4481), .A(N8086), .B(N6685));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2750 (.Y(N4482), .A(N6701), .B(N8133));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2751 (.Y(N4483), .A(N8251), .B(N6711));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2752 (.Y(N4484), .A(N6687), .B(N8261));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2758 (.Y(N4490), .A(N4481), .B(N4483));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2759 (.Y(N4491), .A(N6757), .B(N4482));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5234 (.Y(N4498), .A(N8168), .B(N8121), .C(N4490), .D(N4491));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2760 (.Y(N4492), .A(N8266), .B(N4479));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2761 (.Y(N4493), .A(N4484), .B(N4480));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5235 (.Y(N4500), .AN(N6623), .B(N6715), .C(N8222), .D(N6707));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2765 (.Y(N4497), .A(N4492), .B(N4493));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2767 (.Y(N4499), .A(N4498), .B(N8287));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2769 (.Y(N4501), .A(N4500), .B(N4497));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2770 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[7]), .A(N4499), .B(N4501));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5701 (.Y(N8288), .A(N8081), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2776 (.Y(N4508), .A(N8115), .B(N8203));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2777 (.Y(N4509), .A(N8184), .B(N8217));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2778 (.Y(N4510), .A(N8198), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2779 (.Y(N4511), .A(N8109), .B(N8153));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2781 (.Y(N4513), .A(N6697), .B(N8086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2782 (.Y(N4514), .A(N8190), .B(N8220));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2783 (.Y(N4515), .A(N8212), .B(N8251));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5703 (.Y(N8290), .A(N8237), .B(N8260));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2786 (.Y(N4518), .A(N4299), .B(N4511));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2788 (.Y(N4520), .A(N8288), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2790 (.Y(N4522), .A(N8270), .B(N4508));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2793 (.Y(N4525), .A(N4514), .B(N4513));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2794 (.Y(N4526), .A(N4510), .B(N4515));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2795 (.Y(N4527), .A(N8290), .B(N4509));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2796 (.Y(N4528), .A(N8266), .B(N4520));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2797 (.Y(N4529), .A(N4525), .B(N4526));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2798 (.Y(N4530), .A(N4518), .B(N4527));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2799 (.Y(N4531), .A(N4522), .B(N4528));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I4987 (.Y(N4533), .AN(N8245), .BN(N8253), .C(N8287), .D(N4529));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2802 (.Y(N4534), .A(N4530), .B(N4531));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2803 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[8]), .A(N4534), .B(N4533));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2806 (.Y(N4538), .A(N8179), .B(N8162));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2809 (.Y(N6131), .A(N8109), .B(N8206));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2810 (.Y(N4542), .A(N6677), .B(N8123));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2811 (.Y(N6581), .A(N6729), .B(N8137));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2813 (.Y(N4545), .A(N8223), .B(N6725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2814 (.Y(N4546), .A(N8086), .B(N8190));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2815 (.Y(N4547), .A(N8175), .B(N8133));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2817 (.Y(N4549), .A(N8201), .B(N8165));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2818 (.Y(N6765), .A(N6687), .B(N8156));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2819 (.Y(N4557), .A(N4538), .B(N6131));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2820 (.Y(N4561), .A(N6735), .B(N6727));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2821 (.Y(N4553), .A(N4545), .B(N4547));
NAND2XL hyperpropagate_3_1_A_I5957 (.Y(N8358), .A(N8096), .B(N8198));
NOR2XL hyperpropagate_3_1_A_I5958 (.Y(N4554), .A(N4542), .B(N8358));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5236 (.Y(N4555), .A(N8171), .B(N8147), .C(N6721), .D(N8245));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2824 (.Y(N4556), .A(N4546), .B(N4549));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2827 (.Y(N4559), .A(N6581), .B(N6765));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2831 (.Y(N4563), .A(N4556), .B(N4559));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5237 (.Y(N4567), .A(N4553), .B(N4557), .C(N6101), .D(N4554));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4992 (.Y(N4566), .A(N4555), .B(N4561), .C(N4563));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2836 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[9]), .A(N4567), .B(N4566));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2843 (.Y(N6767), .A(N8183), .B(N8198));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2844 (.Y(N4577), .A(N8161), .B(N8206));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2846 (.Y(N4579), .A(N6681), .B(N8185));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2847 (.Y(N4580), .A(N8113), .B(N8087));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2848 (.Y(N4581), .A(N6685), .B(N8244));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2849 (.Y(N4582), .A(N8257), .B(N8201));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2850 (.Y(N6769), .A(N8230), .B(N8128));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2852 (.Y(N4585), .A(N8215), .B(N8222));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I4994 (.Y(N4592), .A(N8248), .B(N8216), .C(N4389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2854 (.Y(N4587), .A(N6767), .B(N6675));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2855 (.Y(N4588), .A(N4577), .B(N4585));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2856 (.Y(N4589), .A(N4579), .B(N4580));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2857 (.Y(N4590), .A(N4582), .B(N6769));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2861 (.Y(N4594), .A(N4587), .B(N4588));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2862 (.Y(N4598), .A(N4589), .B(N4590));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4996 (.Y(N4600), .A(N4581), .B(N5383), .C(N4594));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4997 (.Y(N4599), .A(N4592), .B(N8266), .C(N4598));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2868 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[10]), .A(N4600), .B(N4599));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2877 (.Y(N4625), .A(N8160), .B(N8153));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2878 (.Y(N4612), .A(N6729), .B(N6697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2879 (.Y(N4613), .A(N8114), .B(N8196));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2880 (.Y(N4614), .A(N8086), .B(N6717));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2882 (.Y(N4616), .A(N8099), .B(N8201));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2883 (.Y(N4617), .A(N8165), .B(N6711));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2884 (.Y(N4618), .A(N8215), .B(N8237));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2885 (.Y(N6771), .A(N8260), .B(N8222));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I4998 (.Y(N4622), .A(N8179), .B(N8081), .C(N6695));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I4999 (.Y(N4635), .A(N168), .B(N6667), .C(N4625));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2893 (.Y(N4627), .A(N4616), .B(N4614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2894 (.Y(N4628), .A(N6757), .B(N6771));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I5238 (.Y(N4630), .AN(N6755), .BN(N6759), .C(N8130), .D(N6727));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2897 (.Y(N4631), .A(N4617));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5001 (.Y(N4638), .AN(N4631), .B(N4613), .C(N4618));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2899 (.Y(N4633), .A(N4612), .B(N4622));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2902 (.Y(N4636), .A(N4635), .B(N4633));
NAND2XL hyperpropagate_3_1_A_I5959 (.Y(N8365), .A(N4627), .B(N4628));
NOR2XL hyperpropagate_3_1_A_I5960 (.Y(N4637), .A(N4630), .B(N8365));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5004 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[11]), .AN(N4636), .B(N4638), .C(N4637));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2914 (.Y(N4648), .A(N8172), .B(N8234));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2915 (.Y(N4649), .A(N8206), .B(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2917 (.Y(N6773), .A(N6733), .B(N6709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2920 (.Y(N6030), .A(N8087), .B(N6701));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2921 (.Y(N4655), .A(N8244), .B(N8128));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2923 (.Y(N4657), .A(N6651), .B(N4648));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2926 (.Y(N4669), .A(N6707), .B(N8288));
NAND2XL hyperpropagate_3_1_A_I5961 (.Y(N8372), .A(N8114), .B(N8202));
NOR2XL hyperpropagate_3_1_A_I5962 (.Y(N4666), .A(N6773), .B(N8372));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2928 (.Y(N4662), .A(N4649), .B(N4655));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2929 (.Y(N4663), .A(N6030), .B(N4263));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5006 (.Y(N4665), .A(N8231), .B(N8136), .C(N4657));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5008 (.Y(N4667), .A(N8165), .B(N8261), .C(N4666));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2934 (.Y(N4671), .A(N4662), .B(N4663));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2936 (.Y(N4673), .A(N4669), .B(N4665));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2938 (.Y(N4672), .A(N4671), .B(N4667));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2940 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[12]), .A(N4673), .B(N4672));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2946 (.Y(N6775), .A(N8119), .B(N8151));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2950 (.Y(N4685), .A(N8227), .B(N6705));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2953 (.Y(N4693), .A(N8147), .B(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2957 (.Y(N4692), .A(N8176), .B(N8230));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2963 (.Y(N4705), .A(N4441), .B(N6753));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2960 (.Y(N6206), .A(N6683), .B(N6715));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5241 (.Y(N4700), .A(N8216), .B(N8203), .C(N8288));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2964 (.Y(N4699), .A(N4482), .B(N4481));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2966 (.Y(N4701), .A(N4700), .B(N6206));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2967 (.Y(N4702), .A(N4685), .B(N4480));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5010 (.Y(N4704), .A(N6775), .B(N6749), .C(N4692));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5011 (.Y(N4709), .AN(N4693), .B(N4705), .C(N8165));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2972 (.Y(N4707), .A(N4699), .B(N4702));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2975 (.Y(N4710), .A(N4709), .B(N4707));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5014 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[13]), .A(N4701), .B(N4704), .C(N4710));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2982 (.Y(N4717), .A(N8080), .B(N8256));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2983 (.Y(N4718), .A(N8162), .B(N8172));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2986 (.Y(N4721), .A(N8231), .B(N8153));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2987 (.Y(N4722), .A(N6729), .B(N6681));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2988 (.Y(N4723), .A(N8113), .B(N8262));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2989 (.Y(N4724), .A(N8196), .B(N8243));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2990 (.Y(N4725), .A(N6717), .B(N8212));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2991 (.Y(N4726), .A(N8099), .B(N8251));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2992 (.Y(N4727), .A(N6711), .B(N8222));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2993 (.Y(N4728), .A(N4717), .B(N4718));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5016 (.Y(N4732), .AN(N8270), .B(N8109), .C(N8248));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2998 (.Y(N4733), .A(N4723), .B(N6775));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2999 (.Y(N4734), .A(N4726), .B(N4727));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3000 (.Y(N4735), .A(N4724), .B(N4725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3001 (.Y(N4739), .A(N4728), .B(N4733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3003 (.Y(N4738), .A(N4734), .B(N4735));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3005 (.Y(N4743), .A(N4739), .B(N4732));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I8629 (.Y(N4742), .AN(N6707), .B(N4722), .C(N4738), .D(N4721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3009 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[14]), .A(N4743), .B(N4742));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3017 (.Y(N6777), .A(N8143), .B(N8248));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3018 (.Y(N6779), .A(N8109), .B(N8160));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3019 (.Y(N4755), .A(N8122), .B(N8153));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3022 (.Y(N4758), .A(N6681), .B(N8098));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3023 (.Y(N5376), .A(N8114), .B(N6725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3024 (.Y(N4760), .A(N8244), .B(N8133));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3025 (.Y(N4761), .A(N8144), .B(N8260));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3026 (.Y(N6781), .A(N8222), .B(N6707));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3027 (.Y(N4763), .A(N6735));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3028 (.Y(N4764), .A(N4763), .B(N6777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3031 (.Y(N4767), .A(N4760), .B(N4761));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5243 (.Y(N4771), .A(N4758), .B(N5376), .C(N6779), .D(N4755));
NAND2XL hyperpropagate_3_1_A_I5963 (.Y(N8379), .A(N8171), .B(N6729));
NOR2XL hyperpropagate_3_1_A_I5964 (.Y(N4769), .A(N6781), .B(N8379));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5244 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[15]), .A(N4767), .B(N4769), .C(N4771), .D(N4764));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3041 (.Y(N6783), .A(N8179), .B(N8193));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3042 (.Y(N4778), .A(N8162), .B(N8253));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3044 (.Y(N4780), .A(N8151), .B(N8216));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3045 (.Y(N4781), .A(N8203), .B(N8143));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3046 (.Y(N4782), .A(N8234), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3047 (.Y(N4783), .A(N8122), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3048 (.Y(N4784), .A(N6681), .B(N8262));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3049 (.Y(N4785), .A(N8147), .B(N8202));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3050 (.Y(N4786), .A(N8244), .B(N8190));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3057 (.Y(N4802), .A(N8280), .B(N4785));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5024 (.Y(N4794), .AN(N4781), .B(N8107), .C(N8171));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3059 (.Y(N4795), .A(N4778), .B(N6759));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3060 (.Y(N4796), .A(N4782), .B(N4783));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3061 (.Y(N4797), .A(N4784), .B(N4780));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3062 (.Y(N4798), .A(N6769), .B(N4786));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3065 (.Y(N4801), .A(N4795), .B(N4796));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5025 (.Y(N4803), .AN(N6783), .B(N8165), .C(N4802));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3068 (.Y(N4806), .A(N4797), .B(N4798));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5026 (.Y(N4808), .A(N4799), .B(N4794), .C(N4801));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3071 (.Y(N4807), .A(N4806), .B(N4803));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3073 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[16]), .A(N4808), .B(N4807));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3083 (.Y(N4820), .A(N8248), .B(N6677));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3084 (.Y(N4821), .A(N8122), .B(N6709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3086 (.Y(N4823), .A(N6717), .B(N8220));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5027 (.Y(N4838), .A(N8134), .B(N8172), .C(N8165));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3092 (.Y(N4829), .A(N8156), .B(N8238));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3093 (.Y(N6785), .A(N6679), .B(N8132));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3094 (.Y(N4831), .A(N4820), .B(N4829));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3095 (.Y(N4832), .A(N4692), .B(N4823));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3096 (.Y(N4833), .A(N6751), .B(N4821));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5028 (.Y(N4834), .AN(N6785), .B(N8227), .C(N8251));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5029 (.Y(N4836), .A(N8253), .B(N8151), .C(N4831));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3100 (.Y(N4837), .A(N4832), .B(N4833));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3102 (.Y(N4839), .A(N4838), .B(N4834));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3103 (.Y(N4841), .A(N4836), .B(N4837));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3105 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[17]), .A(N4841), .B(N4839));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3116 (.Y(N4854), .A(N6653), .B(N8077));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3117 (.Y(N4855), .A(N8248), .B(N8122));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3120 (.Y(N4858), .A(N8196), .B(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3121 (.Y(N4859), .A(N8175), .B(N8230));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3122 (.Y(N4868), .A(N4854), .B(N8165));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3123 (.Y(N4861), .A(N8131), .B(N6735));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3125 (.Y(N4863), .A(N4859), .B(N4855));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5030 (.Y(N4870), .AN(N4427), .B(N8136), .C(N6721));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5633 (.Y(N8313), .A(N8266));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3129 (.Y(N4867), .A(N8313), .B(N4863));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5031 (.Y(N4872), .A(N4868), .B(N4861), .C(N4858));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3133 (.Y(N4871), .A(N4870), .B(N4867));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3135 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[18]), .A(N4872), .B(N4871));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3146 (.Y(N5222), .A(N6697), .B(N8137));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3148 (.Y(N4886), .A(N6717), .B(N8230));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3149 (.Y(N6787), .A(N8215), .B(N8156));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3150 (.Y(N4888), .A(N8238), .B(N8131));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5245 (.Y(N4892), .A(N8168), .B(N8245), .C(N6701), .D(N8197));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3153 (.Y(N4891), .A(N4886), .B(N4888));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3155 (.Y(N4893), .A(N4892), .B(N6787));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3156 (.Y(N4894), .A(N5222), .B(N4427));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5033 (.Y(N4896), .A(N8121), .B(N6729), .C(N4891));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5035 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[19]), .AN(N4896), .B(N4894), .C(N4893));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3171 (.Y(N4909), .A(N6677), .B(N8231));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3172 (.Y(N4910), .A(N6681), .B(N6721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3174 (.Y(N4912), .A(N6685), .B(N6717));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3175 (.Y(N6789), .A(N6687), .B(N8215));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3176 (.Y(N4914), .A(N6679), .B(N8222));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3178 (.Y(N4916), .A(N8280), .B(N4909));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3180 (.Y(N4918), .A(N8270), .B(N6789));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3181 (.Y(N4919), .A(N4910), .B(N4912));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5036 (.Y(N4922), .AN(N4914), .B(N8197), .C(N6725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3183 (.Y(N4921), .A(N4916), .B(N4919));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3185 (.Y(N4923), .A(N4922), .B(N4921));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3186 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[20]), .A(N4918), .B(N4923));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3196 (.Y(N4934), .A(N8136), .B(N6681));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3198 (.Y(N4936), .A(N6701), .B(N6711));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3201 (.Y(N4939), .A(N6707), .B(N6683));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3204 (.Y(N4942), .A(N4936), .B(N4542));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3205 (.Y(N4943), .A(N6785), .B(N6747));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3207 (.Y(N4945), .A(N4330));
NAND3XL hyperpropagate_4_1_A_I5965 (.Y(N8388), .A(N6709), .B(N6685), .C(N4945));
NOR2XL hyperpropagate_4_1_A_I5966 (.Y(N4950), .A(N6765), .B(N8388));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3209 (.Y(N4947), .A(N4942), .B(N4943));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5038 (.Y(N4949), .A(N4939), .B(N4934), .C(N4947));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3213 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[21]), .A(N4950), .B(N4949));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3240 (.Y(N4978), .A(N6729), .B(N8098));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3241 (.Y(N4979), .A(N6721), .B(N8190));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3244 (.Y(N4982), .A(N8251), .B(N8128));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3245 (.Y(N5483), .A(N8165), .B(N8156));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5039 (.Y(N4992), .AN(N6779), .B(N8176), .C(N8201));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3250 (.Y(N4988), .A(N6775), .B(N4982));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3251 (.Y(N4989), .A(N4979), .B(N4799));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5040 (.Y(N4991), .AN(N8290), .B(N6727), .C(N4260));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3256 (.Y(N4994), .A(N4988), .B(N4989));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3257 (.Y(N4995), .A(N4978), .B(N5483));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3258 (.Y(N4998), .A(N4991), .B(N4994));
NAND3XL hyperpropagate_4_1_A_I5967 (.Y(N8396), .A(N4976), .B(N6705), .C(N4995));
NOR2XL hyperpropagate_4_1_A_I5968 (.Y(N4997), .A(N4992), .B(N8396));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3261 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[23]), .A(N4998), .B(N4997));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3269 (.Y(N5007), .A(N8245), .B(N8150));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3270 (.Y(N5008), .A(N8107), .B(N8235));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3271 (.Y(N5009), .A(N8216), .B(N8183));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3272 (.Y(N5010), .A(N8198), .B(N8121));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3273 (.Y(N5011), .A(N8223), .B(N8202));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3274 (.Y(N5012), .A(N8243), .B(N6701));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3275 (.Y(N5013), .A(N8175), .B(N8257));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3282 (.Y(N5020), .A(N8287), .B(N5009));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3283 (.Y(N5021), .A(N5008), .B(N5007));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5043 (.Y(N5023), .A(N5013), .B(N5011), .C(N5012));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3286 (.Y(N5024), .A(N4982), .B(N6789));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5044 (.Y(N5025), .A(N8227), .B(N8081), .C(N6679), .D(N5021));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3288 (.Y(N5026), .A(N5010), .B(N5025));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5248 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[24]), .A(N5020), .B(N5023), .C(N5024), .D(N5026));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3300 (.Y(N5039), .A(N8162), .B(N8150));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3301 (.Y(N5040), .A(N8171), .B(N8234));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3303 (.Y(N5042), .A(N8168), .B(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3304 (.Y(N5043), .A(N6721), .B(N8114));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3308 (.Y(N5047), .A(N8144), .B(N8131));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3309 (.Y(N5048), .A(N5042), .B(N5039));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3310 (.Y(N5049), .A(N6635), .B(N5040));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5046 (.Y(N5050), .AN(N6745), .B(N8183), .C(N8206));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3312 (.Y(N5051), .A(N5048), .B(N5049));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3315 (.Y(N5054), .A(N5053), .B(N5050));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3316 (.Y(N5055), .A(N5047), .B(N5051));
NAND3XL hyperpropagate_4_1_A_I5969 (.Y(N8404), .A(N6685), .B(N8201), .C(N5055));
NOR2XL hyperpropagate_4_1_A_I5970 (.Y(N5056), .A(N5043), .B(N8404));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3318 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[25]), .A(N5054), .B(N5056));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3328 (.Y(N5067), .A(N8136), .B(N8262));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3332 (.Y(N5071), .A(N8176), .B(N8099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3334 (.Y(N5073), .A(N6711), .B(N6687));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3335 (.Y(N5081), .A(N6735), .B(N6703));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5250 (.Y(N5075), .A(N8147), .B(N8152), .C(N8202), .D(N8243));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5251 (.Y(N5076), .A(N8234), .B(N8172), .C(N8248), .D(N8096));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3339 (.Y(N5085), .A(N5073), .B(N6030));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3341 (.Y(N5080), .A(N6769), .B(N5075));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3343 (.Y(N5087), .A(N5081), .B(N5076));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5050 (.Y(N5084), .A(N5071), .B(N6767), .C(N5067));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5252 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[26]), .A(N5085), .B(N5084), .C(N5080), .D(N5087));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3358 (.Y(N5098), .A(N8171), .B(N8143));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3362 (.Y(N5102), .A(N8224), .B(N8206));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3364 (.Y(N5573), .A(N6729), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3365 (.Y(N5105), .A(N6685), .B(N8133));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3366 (.Y(N5106), .A(N8212), .B(N8176));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3367 (.Y(N5117), .A(N8201), .B(N8251));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3368 (.Y(N5108), .A(N6711), .B(N6679));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3369 (.Y(N5109), .A(N8260), .B(N6727));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3373 (.Y(N5121), .A(N5108), .B(N6767));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5052 (.Y(N5115), .A(N102), .B(N8076), .C(N5106));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3376 (.Y(N5116), .A(N5105), .B(N5109));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5054 (.Y(N5120), .A(N5102), .B(N5098), .C(N4755));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3382 (.Y(N5126), .A(N5121), .B(N5573));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3383 (.Y(N5123), .A(N5116), .B(N5115));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I5055 (.Y(N5128), .AN(N5120), .B(N5117), .C(N5039), .D(N8279));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3387 (.Y(N5127), .A(N5126), .B(N5123));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3389 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[27]), .A(N5128), .B(N5127));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3395 (.Y(N5135), .A(N8179), .B(N8150));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3402 (.Y(N5142), .A(N8087), .B(N6685));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3403 (.Y(N5143), .A(N6717), .B(N8128));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5056 (.Y(N5151), .AN(N6651), .B(N8098), .C(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3408 (.Y(N5148), .A(N6711), .B(N6707));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5058 (.Y(N5156), .AN(N4352), .B(N8118), .C(N8248));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3412 (.Y(N5152), .A(N5151), .B(N5143));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3413 (.Y(N5153), .A(N5142), .B(N4858));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5059 (.Y(N5155), .A(N5148), .B(N6753), .C(N6757));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5060 (.Y(N5157), .AN(N8165), .B(N5135), .C(N5156));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5253 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[28]), .A(N5153), .B(N5157), .C(N5155), .D(N5152));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3433 (.Y(N5174), .A(N8193), .B(N6705));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3434 (.Y(N5175), .A(N6729), .B(N8113));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3440 (.Y(N5181), .A(N8287), .B(N4760));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3444 (.Y(N5189), .A(N5174), .B(N6781));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5254 (.Y(N5186), .A(N4577), .B(N4350), .C(N6777), .D(N6775));
NAND3XL hyperpropagate_4_1_A_I5971 (.Y(N8412), .A(N6721), .B(N8202), .C(N5175));
NOR2XL hyperpropagate_4_1_A_I5972 (.Y(N5188), .A(N4561), .B(N8412));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5256 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[29]), .A(N5181), .B(N5186), .C(N5189), .D(N5188));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3467 (.Y(N5209), .A(N8147), .B(N6701));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3468 (.Y(N5210), .A(N8244), .B(N8257));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3470 (.Y(N5220), .A(N8222), .B(N8130));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5065 (.Y(N5213), .AN(N6683), .B(N163), .C(N8076));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3473 (.Y(N5215), .A(N4263), .B(N5210));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3474 (.Y(N5216), .A(N6741), .B(N5222));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5066 (.Y(N5219), .A(N5209), .B(N6755), .C(N4721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3479 (.Y(N5221), .A(N5220), .B(N5215));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3481 (.Y(N5223), .A(N5213), .B(N5216));
NAND3XL hyperpropagate_4_1_A_I5973 (.Y(N8420), .A(N8252), .B(N8201), .C(N5219));
NOR2XL hyperpropagate_4_1_A_I5974 (.Y(N5226), .A(N5102), .B(N8420));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3483 (.Y(N5225), .A(N5221), .B(N5223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3485 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[30]), .A(N5226), .B(N5225));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3493 (.Y(N5235), .A(N8160), .B(N6677));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3499 (.Y(N5241), .A(N8099), .B(N8230));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3502 (.Y(N6791), .A(N6679), .B(N8260));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5258 (.Y(N5247), .A(N8147), .B(N8244), .C(N6697), .D(N6681));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3506 (.Y(N5248), .A(N5235), .B(N6777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3507 (.Y(N5249), .A(N4782), .B(N5241));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3508 (.Y(N5250), .A(N6791), .B(N5106));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3511 (.Y(N5253), .A(N5248), .B(N5249));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5070 (.Y(N5255), .A(N8179), .B(N8172), .C(N8165), .D(N5250));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5071 (.Y(N5257), .A(N4299), .B(N4514), .C(N5253));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5072 (.Y(N5258), .A(N6751), .B(N5247), .C(N5255));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3517 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[31]), .A(N5257), .B(N5258));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3523 (.Y(N5265), .A(N8081), .B(N8115));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3524 (.Y(N5282), .A(N8171), .B(N8151));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3526 (.Y(N5268), .A(N8096), .B(N8168));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3527 (.Y(N5269), .A(N6737), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3528 (.Y(N5270), .A(N8262), .B(N8098));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3530 (.Y(N5272), .A(N6725), .B(N8087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3534 (.Y(N5276), .A(N5270), .B(N5265));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3536 (.Y(N5284), .A(N4693), .B(N5272));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5073 (.Y(N5280), .A(N8156), .B(N6727), .C(N5276));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3539 (.Y(N5281), .A(N5269), .B(N5268));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5075 (.Y(N5289), .A(N6711), .B(N8128), .C(N5284));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5076 (.Y(N5287), .A(N6701), .B(N8176), .C(N5281));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5077 (.Y(N5288), .A(N5282), .B(N4781), .C(N6783), .D(N5280));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3548 (.Y(N5290), .A(N5289), .B(N5287));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3549 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[32]), .A(N5288), .B(N5290));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3554 (.Y(N5296), .A(N8134), .B(N8245));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3555 (.Y(N5297), .A(N8253), .B(N8119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3556 (.Y(N5298), .A(N8107), .B(N8216));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3560 (.Y(N5302), .A(N8098), .B(N8114));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3563 (.Y(N5305), .A(N8230), .B(N8144));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3566 (.Y(N5308), .A(N5302), .B(N5296));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3567 (.Y(N5314), .A(N5298), .B(N5297));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5078 (.Y(N5316), .AN(N6745), .B(N6697), .C(N6709));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5079 (.Y(N5320), .A(N8198), .B(N8160), .C(N5308));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3573 (.Y(N5315), .A(N5314), .B(N5305));
NAND3XL hyperpropagate_4_1_A_I5975 (.Y(N8428), .A(N8201), .B(N8244), .C(N8265));
NOR2XL hyperpropagate_4_1_A_I5976 (.Y(N5319), .A(N4914), .B(N8428));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3579 (.Y(N5321), .A(N5320), .B(N5315));
NAND3XL hyperpropagate_4_1_A_I5977 (.Y(N8436), .A(N8130), .B(N6703), .C(N5319));
NOR2XL hyperpropagate_4_1_A_I5978 (.Y(N5322), .A(N5316), .B(N8436));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3581 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[33]), .A(N5321), .B(N5322));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3587 (.Y(N5329), .A(N8256), .B(N8134));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3589 (.Y(N5331), .A(N8150), .B(N8115));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3590 (.Y(N5332), .A(N8216), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3595 (.Y(N5337), .A(N6717), .B(N8190));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3598 (.Y(N5340), .A(N6671), .B(N5329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3599 (.Y(N5341), .A(N8128), .B(N8215));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5083 (.Y(N5350), .AN(N4291), .B(N8147), .C(N8114));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3604 (.Y(N5346), .A(N6753), .B(N5337));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3607 (.Y(N5349), .A(N5332), .B(N4356));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3609 (.Y(N5351), .A(N5350), .B(N5341));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5085 (.Y(N5353), .A(N8231), .B(N8109), .C(N6707), .D(N5346));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3612 (.Y(N5354), .A(N5340), .B(N5349));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I5086 (.Y(N5357), .AN(N5351), .B(N6783), .C(N4758), .D(N5331));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3614 (.Y(N5356), .A(N5354), .B(N5353));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3616 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[34]), .A(N5357), .B(N5356));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3622 (.Y(N5364), .A(N8134), .B(N8150));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3623 (.Y(N5365), .A(N8171), .B(N8235));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3624 (.Y(N5366), .A(N8216), .B(N8160));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3626 (.Y(N5368), .A(N8243), .B(N6685));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3627 (.Y(N5369), .A(N6717), .B(N8133));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3629 (.Y(N5371), .A(N8201), .B(N8230));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3631 (.Y(N5373), .A(N6711), .B(N8215));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3633 (.Y(N5375), .A(N5364), .B(N5365));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3635 (.Y(N5377), .A(N5376), .B(N5371));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3636 (.Y(N5378), .A(N5373), .B(N5369));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3637 (.Y(N5379), .A(N5366), .B(N5368));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5087 (.Y(N5380), .AN(N5071), .B(N8156), .C(N6735));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3639 (.Y(N5385), .A(N5375), .B(N5377));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3640 (.Y(N5382), .A(N5378), .B(N5379));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3642 (.Y(N5387), .A(N5383), .B(N5380));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3644 (.Y(N5386), .A(N5385), .B(N5382));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3646 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[35]), .A(N5387), .B(N5386));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3651 (.Y(N5394), .A(N8150), .B(N8235));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3654 (.Y(N5397), .A(N6677), .B(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3655 (.Y(N5398), .A(N8231), .B(N6705));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3659 (.Y(N5402), .A(N8244), .B(N8220));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3660 (.Y(N5403), .A(N8213), .B(N6679));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3662 (.Y(N5740), .A(N6683), .B(N6695));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5260 (.Y(N5408), .A(N4781), .B(N5394), .C(N5397), .D(N140));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3666 (.Y(N5409), .A(N5402), .B(N5403));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3667 (.Y(N5410), .A(N4579), .B(N5043));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3669 (.Y(N5412), .A(N4326), .B(N5398));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3670 (.Y(N5416), .A(N5740), .B(N5408));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3671 (.Y(N5414), .A(N5409), .B(N5410));
NAND3XL hyperpropagate_4_1_A_I5979 (.Y(N8444), .A(N5412), .B(N8261), .C(N6735));
NOR2XL hyperpropagate_4_1_A_I5980 (.Y(N5418), .A(N4510), .B(N8444));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3674 (.Y(N5417), .A(N5416), .B(N5414));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3676 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[36]), .A(N5418), .B(N5417));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3682 (.Y(N5426), .A(N8097), .B(N8162));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3683 (.Y(N5427), .A(N8107), .B(N8115));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3685 (.Y(N5429), .A(N8143), .B(N8153));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3687 (.Y(N5431), .A(N8185), .B(N8098));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5090 (.Y(N5437), .AN(N6651), .B(N8201), .C(N8133));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3699 (.Y(N5443), .A(N5427), .B(N5365));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3700 (.Y(N5444), .A(N5429), .B(N6773));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5093 (.Y(N5451), .AN(N5431), .B(N8080), .C(N8220));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5094 (.Y(N5447), .AN(N6789), .B(N8175), .C(N8237), .D(N8086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3704 (.Y(N5448), .A(N5443), .B(N5444));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3708 (.Y(N5452), .A(N5451), .B(N5448));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5095 (.Y(N5456), .AN(N8165), .B(N5426), .C(N5447));
NAND3XL hyperpropagate_4_1_A_I5981 (.Y(N8452), .A(N8227), .B(N8193), .C(N5452));
NOR2XL hyperpropagate_4_1_A_I5982 (.Y(N5455), .A(N5437), .B(N8452));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3713 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[37]), .A(N5456), .B(N5455));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3722 (.Y(N5466), .A(N8172), .B(N8115));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3725 (.Y(N5469), .A(N6709), .B(N8147));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3726 (.Y(N5569), .A(N6725), .B(N6685));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3730 (.Y(N5474), .A(N6647), .B(N5466));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5097 (.Y(N5477), .A(N8143), .B(N8234), .C(N6727));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3734 (.Y(N5478), .A(N5469), .B(N5337));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5098 (.Y(N5480), .AN(N5477), .B(N6677), .C(N6681));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3738 (.Y(N5482), .A(N5478), .B(N5474));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5099 (.Y(N5484), .A(N5569), .B(N4356), .C(N5483));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3741 (.Y(N5486), .A(N5480), .B(N5482));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3743 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[38]), .A(N5486), .B(N5484));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3754 (.Y(N5498), .A(N6677), .B(N6705));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3755 (.Y(N5506), .A(N6697), .B(N6721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3756 (.Y(N5500), .A(N8223), .B(N6685));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3757 (.Y(N5501), .A(N6717), .B(N8201));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3758 (.Y(N6180), .A(N8165), .B(N6687));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3760 (.Y(N5504), .A(N6707), .B(N6695));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5263 (.Y(N5505), .A(N8143), .B(N8215), .C(N8118), .D(N6679));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3763 (.Y(N5512), .A(N5506), .B(N5505));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3764 (.Y(N5510), .A(N5498), .B(N5500));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3765 (.Y(N5509), .A(N5504), .B(N5501));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5264 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[39]), .A(N6180), .B(N5510), .C(N5509), .D(N5512));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3777 (.Y(N5522), .A(N6677), .B(N8168));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3779 (.Y(N6272), .A(N6697), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3781 (.Y(N5526), .A(N6725), .B(N6701));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3784 (.Y(N5529), .A(N8238), .B(N6679));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3786 (.Y(N6793), .A(N6735), .B(N6683));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3787 (.Y(N6546), .A(N6727), .B(N6695));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3788 (.Y(N5533), .A(N5522), .B(N122));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3789 (.Y(N5539), .A(N5529), .B(N6272));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3790 (.Y(N5535), .A(N6787), .B(N6771));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3791 (.Y(N5536), .A(N5526));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3792 (.Y(N5543), .A(N5536), .B(N5533));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3793 (.Y(N5538), .A(N4910), .B(N6793));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3795 (.Y(N5540), .A(N5539), .B(N6546));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5102 (.Y(N5541), .AN(N5501), .B(N6737), .C(N6729));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3797 (.Y(N5545), .A(N5535), .B(N5538));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3799 (.Y(N5544), .A(N5543), .B(N5541));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3801 (.Y(N5546), .A(N5545), .B(N5540));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3802 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[40]), .A(N5544), .B(N5546));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3810 (.Y(N5555), .A(N6737), .B(N8121));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5103 (.Y(N5565), .AN(N5555), .B(N8134), .C(N6677));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5104 (.Y(N5571), .AN(N5529), .B(N6727), .C(N6683));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3822 (.Y(N5567), .A(N6789), .B(N6771));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3829 (.Y(N5574), .A(N5573), .B(N5567));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5265 (.Y(N5576), .A(N4910), .B(N5569), .C(N4861), .D(N5565));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5106 (.Y(N5578), .A(N5501), .B(N5571), .C(N5574));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3834 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[41]), .A(N5576), .B(N5578));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3844 (.Y(N5589), .A(N6709), .B(N8196));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3851 (.Y(N5596), .A(N5589), .B(N4542));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3853 (.Y(N5598), .A(N4934), .B(N6747));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3854 (.Y(N5599), .A(N6785), .B(N4939));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5107 (.Y(N5601), .A(N8202), .B(N6685), .C(N5596));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5108 (.Y(N5606), .AN(N4945), .B(N4936), .C(N6765));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3859 (.Y(N5604), .A(N5598), .B(N5599));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3860 (.Y(N5605), .A(N5601), .B(N5604));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3862 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[42]), .A(N5606), .B(N5605));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3868 (.Y(N5614), .A(N8245), .B(N8119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3870 (.Y(N5629), .A(N8096), .B(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3874 (.Y(N5620), .A(N8113), .B(N8207));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3882 (.Y(N5628), .A(N5614), .B(N5620));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5110 (.Y(N5632), .A(N8216), .B(N8143), .C(N5628));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3887 (.Y(N5633), .A(N6793), .B(N6785));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5111 (.Y(N5634), .A(N6655), .B(N6627), .C(N6747), .D(N5629));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5112 (.Y(N5636), .A(N161), .B(N5013), .C(N4581));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3891 (.Y(N5637), .A(N5632), .B(N4617));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5266 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[43]), .A(N5636), .B(N5634), .C(N5637), .D(N5633));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3908 (.Y(N5655), .A(N6685), .B(N8213));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3911 (.Y(N5658), .A(N6679), .B(N6735));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3914 (.Y(N5661), .A(N8279), .B(N4718));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5267 (.Y(N5662), .A(N8234), .B(N8143), .C(N8198), .D(N8253));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5116 (.Y(N5663), .A(N6715), .B(N6727));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5117 (.Y(N5664), .AN(N6627), .B(N6733), .C(N5663));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5118 (.Y(N5666), .A(N6711), .B(N8099), .C(N5661));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5119 (.Y(N5671), .AN(N6304), .B(N8153), .C(N6697));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3922 (.Y(N5669), .A(N5668), .B(N5662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3923 (.Y(N5674), .A(N5658), .B(N6741));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3925 (.Y(N5672), .A(N5671), .B(N5655));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3926 (.Y(N5673), .A(N5664), .B(N5666));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5268 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[44]), .A(N5669), .B(N5674), .C(N5672), .D(N5673));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3939 (.Y(N5687), .A(N8151), .B(N8096));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3943 (.Y(N5691), .A(N8257), .B(N8099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3944 (.Y(N6795), .A(N8128), .B(N8144));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3945 (.Y(N5693), .A(N6627), .B(N5691));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3950 (.Y(N5698), .A(N5296), .B(N5687));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5121 (.Y(N5700), .A(N8183), .B(N8160), .C(N5693));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3954 (.Y(N5702), .A(N5663), .B(N5698));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5122 (.Y(N5708), .AN(N6789), .B(N8237), .C(N6707));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5123 (.Y(N5707), .A(N5702), .B(N4614), .C(N6795));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3961 (.Y(N5711), .A(N5708), .B(N4617));
NAND3XL hyperpropagate_4_1_A_I5983 (.Y(N8460), .A(N6705), .B(N6725), .C(N5707));
NOR2XL hyperpropagate_4_1_A_I5984 (.Y(N5710), .A(N5700), .B(N8460));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3964 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[45]), .A(N5711), .B(N5710));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3972 (.Y(N5721), .A(N8160), .B(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3973 (.Y(N5722), .A(N6709), .B(N8185));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3975 (.Y(N5901), .A(N8202), .B(N8086));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5125 (.Y(N5733), .AN(N6627), .B(N8257), .C(N8252));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5126 (.Y(N5732), .AN(N5901), .B(N8235), .C(N8151));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3985 (.Y(N5734), .A(N5733), .B(N5722));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3986 (.Y(N5735), .A(N5721), .B(N6777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3988 (.Y(N5737), .A(N6787), .B(N5732));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3989 (.Y(N5738), .A(N6751), .B(N4357));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3992 (.Y(N5741), .A(N5740), .B(N5735));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3993 (.Y(N5742), .A(N5734), .B(N5738));
NAND3XL hyperpropagate_4_1_A_I5985 (.Y(N8468), .A(N8244), .B(N6717), .C(N5737));
NOR2XL hyperpropagate_4_1_A_I5986 (.Y(N5744), .A(N6781), .B(N8468));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3996 (.Y(N5745), .A(N5742), .B(N5741));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3997 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[46]), .A(N5745), .B(N5744));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4004 (.Y(N5754), .A(N8256), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4009 (.Y(N5759), .A(N8098), .B(N8243));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4012 (.Y(N5763), .A(N8175), .B(N8252));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4017 (.Y(N5767), .A(N8287), .B(N5039));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5128 (.Y(N5769), .A(N6623), .B(N4648), .C(N5754));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4020 (.Y(N5770), .A(N5759), .B(N4323));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5129 (.Y(N5772), .A(N8183), .B(N8153), .C(N5770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4024 (.Y(N5774), .A(N5663), .B(N5769));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4026 (.Y(N5778), .A(N4912), .B(N5774));
NAND3XL hyperpropagate_4_1_A_I5987 (.Y(N8476), .A(N5763), .B(N8130), .C(N5767));
NOR2XL hyperpropagate_4_1_A_I5988 (.Y(N5777), .A(N5772), .B(N8476));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4029 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[47]), .A(N5778), .B(N5777));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4037 (.Y(N5788), .A(N8256), .B(N8162));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4038 (.Y(N5789), .A(N8198), .B(N8109));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4039 (.Y(N5790), .A(N6705), .B(N8136));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4041 (.Y(N5792), .A(N8113), .B(N6721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4043 (.Y(N5794), .A(N8133), .B(N8099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4044 (.Y(N5795), .A(N8201), .B(N8238));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4047 (.Y(N5798), .A(N6627), .B(N5788));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4048 (.Y(N5799), .A(N5794), .B(N5789));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4049 (.Y(N5800), .A(N5798), .B(N5799));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4050 (.Y(N5801), .A(N6771), .B(N5792));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4051 (.Y(N5802), .A(N5800), .B(N6741));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4052 (.Y(N5803), .A(N5081), .B(N5795));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4053 (.Y(N5804), .A(N5790), .B(N4327));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5272 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[48]), .A(N5804), .B(N5803), .C(N5802), .D(N5801));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4067 (.Y(N5818), .A(N8262), .B(N6721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4068 (.Y(N5830), .A(N8197), .B(N8152));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4069 (.Y(N6797), .A(N8202), .B(N6725));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4078 (.Y(N5834), .A(N6797), .B(N4577));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5133 (.Y(N5838), .A(N4546), .B(N5830), .C(N5042));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4081 (.Y(N5832), .A(N4783), .B(N4618));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4082 (.Y(N5833), .A(N6769), .B(N5818));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5134 (.Y(N5842), .A(N8235), .B(N8109), .C(N6681), .D(N5834));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4085 (.Y(N5836), .A(N6781), .B(N6793));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4086 (.Y(N5837), .A(N5832), .B(N5833));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4088 (.Y(N5839), .A(N5838), .B(N5836));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5135 (.Y(N5841), .A(N5364), .B(N8287), .C(N5837));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4092 (.Y(N5843), .A(N5842), .B(N5839));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4093 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[49]), .A(N5841), .B(N5843));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4099 (.Y(N5851), .A(N8234), .B(N8217));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4103 (.Y(N5855), .A(N8262), .B(N8147));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4106 (.Y(N6028), .A(N8190), .B(N8213));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4109 (.Y(N5861), .A(N8222), .B(N6735));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4110 (.Y(N5862), .A(N5855), .B(N114));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4111 (.Y(N5863), .A(N5851), .B(N5789));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4112 (.Y(N5864), .A(N5397), .B(N6028));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5136 (.Y(N5866), .A(N8086), .B(N8244), .C(N5862));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5137 (.Y(N5867), .AN(N6797), .B(N8231), .C(N6709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4116 (.Y(N5868), .A(N5863), .B(N5864));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4119 (.Y(N5871), .A(N5861), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4120 (.Y(N5875), .A(N5866), .B(N5483));
NAND3XL hyperpropagate_4_1_A_I5989 (.Y(N8484), .A(N8099), .B(N8128), .C(N5871));
NOR2XL hyperpropagate_4_1_A_I5990 (.Y(N5874), .A(N5867), .B(N8484));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4124 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[50]), .A(N5875), .B(N5874));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4135 (.Y(N5888), .A(N6659), .B(N8076));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4137 (.Y(N5890), .A(N6697), .B(N8262));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4142 (.Y(N5895), .A(N8230), .B(N8131));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5140 (.Y(N5900), .A(N8245), .B(N8203), .C(N5888));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5141 (.Y(N5902), .AN(N5901), .B(N8109), .C(N5763), .D(N8217));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4151 (.Y(N5904), .A(N5890), .B(N5900));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4152 (.Y(N5905), .A(N5895), .B(N5902));
NAND3XL hyperpropagate_4_1_A_I5991 (.Y(N8492), .A(N8313), .B(N8098), .C(N8197));
NOR2XL hyperpropagate_4_1_A_I5992 (.Y(N5911), .A(N4786), .B(N8492));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4155 (.Y(N5908), .A(N5904), .B(N5905));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5143 (.Y(N5910), .A(N5426), .B(N8287), .C(N5908));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4159 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[51]), .A(N5911), .B(N5910));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4167 (.Y(N5921), .A(N8134), .B(N8253));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4169 (.Y(N5923), .A(N8183), .B(N8109));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4170 (.Y(N5924), .A(N8206), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4171 (.Y(N5925), .A(N8098), .B(N8152));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4173 (.Y(N5927), .A(N8080), .B(N6701));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5144 (.Y(N5935), .AN(N5921), .B(N8115), .C(N8216));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4176 (.Y(N5930), .A(N8165), .B(N8222));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4179 (.Y(N5933), .A(N8270), .B(N5924));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4180 (.Y(N5937), .A(N5925), .B(N5923));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4182 (.Y(N5936), .A(N5935), .B(N5927));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4184 (.Y(N5938), .A(N5937), .B(N5305));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4185 (.Y(N5939), .A(N5933), .B(N5936));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4187 (.Y(N5941), .A(N4276), .B(N5938));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4188 (.Y(N5943), .A(N5939), .B(N5930));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4190 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[52]), .A(N5943), .B(N5941));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4201 (.Y(N5956), .A(N6677), .B(N8113));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4204 (.Y(N5959), .A(N8175), .B(N8213));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5145 (.Y(N5965), .A(N8171), .B(N8216), .C(N6727));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4211 (.Y(N5966), .A(N5011), .B(N6767));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4212 (.Y(N5967), .A(N5956), .B(N5959));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5147 (.Y(N5974), .AN(N6791), .B(N6725), .C(N8244));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4216 (.Y(N5971), .A(N5966), .B(N5967));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4218 (.Y(N5973), .A(N6795), .B(N5965));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4220 (.Y(N5975), .A(N5974), .B(N5971));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I5148 (.Y(N5976), .AN(N5973), .B(N6643), .C(N6779), .D(N8076));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4222 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[53]), .A(N5975), .B(N5976));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4230 (.Y(N6306), .A(N8096), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4231 (.Y(N5986), .A(N6677), .B(N6697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4234 (.Y(N5989), .A(N8197), .B(N8147));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4235 (.Y(N5990), .A(N8223), .B(N8152));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4237 (.Y(N5996), .A(N8190), .B(N8252));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5275 (.Y(N5994), .A(N8172), .B(N8114), .C(N8207), .D(N8253));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4240 (.Y(N5999), .A(N5990), .B(N6306));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4242 (.Y(N6002), .A(N5996), .B(N5994));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4243 (.Y(N5998), .A(N4479), .B(N5986));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4245 (.Y(N6000), .A(N5999), .B(N5989));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4246 (.Y(N6001), .A(N4614), .B(N4451));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5276 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[54]), .A(N6000), .B(N6001), .C(N5998), .D(N6002));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4258 (.Y(N6014), .A(N8224), .B(N6729));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4264 (.Y(N6020), .A(N8256), .B(N6717));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5151 (.Y(N6027), .AN(N5302), .B(N8216), .C(N8096));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5152 (.Y(N6029), .A(N6028), .B(N8279), .C(N6755));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4277 (.Y(N6033), .A(N6014), .B(N5117));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4278 (.Y(N6034), .A(N6795), .B(N6020));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5153 (.Y(N6039), .A(N6707), .B(N6727), .C(N6029));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5277 (.Y(N6037), .A(N6030), .B(N5830), .C(N6027), .D(N6272));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4282 (.Y(N6038), .A(N6033), .B(N6034));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4284 (.Y(N6040), .A(N6039), .B(N6038));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4285 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[55]), .A(N6037), .B(N6040));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4293 (.Y(N6050), .A(N8151), .B(N8203));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4299 (.Y(N6067), .A(N8244), .B(N8230));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4304 (.Y(N6061), .A(N8279), .B(N5921));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4307 (.Y(N6064), .A(N4351), .B(N6050));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5278 (.Y(N6066), .A(N8114), .B(N6701), .C(N6679), .D(N8144));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5157 (.Y(N6073), .A(N115), .B(N6667), .C(N6067), .D(N4511));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5158 (.Y(N6075), .A(N8130), .B(N6707), .C(N5573));
NAND3XL hyperpropagate_4_1_A_I5993 (.Y(N8500), .A(N6073), .B(N6064), .C(N6061));
NOR2XL hyperpropagate_4_1_A_I5994 (.Y(N6077), .A(N4784), .B(N8500));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5160 (.Y(N6076), .A(N6066), .B(N6793), .C(N6075));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4321 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[56]), .A(N6077), .B(N6076));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4325 (.Y(N6082), .A(N8162), .B(N8107));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4326 (.Y(N6083), .A(N8115), .B(N8235));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4332 (.Y(N6089), .A(N8113), .B(N8243));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4333 (.Y(N6482), .A(N8190), .B(N8175));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4336 (.Y(N6093), .A(N6671), .B(N6083));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4340 (.Y(N6097), .A(N8287), .B(N6089));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4341 (.Y(N6098), .A(N6082), .B(N6050));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4342 (.Y(N6099), .A(N4509), .B(N4510));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4343 (.Y(N6100), .A(N6777), .B(N6482));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4345 (.Y(N6102), .A(N6101), .B(N6093));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5161 (.Y(N6105), .A(N8222), .B(N6727), .C(N6100));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5162 (.Y(N6108), .AN(N4421), .B(N8153), .C(N6681));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4352 (.Y(N6109), .A(N6108), .B(N6105));
NAND3XL hyperpropagate_4_1_A_I5995 (.Y(N8508), .A(N6098), .B(N6099), .C(N6097));
NOR2XL hyperpropagate_4_1_A_I5996 (.Y(N6111), .A(N6102), .B(N8508));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4355 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[57]), .A(N6111), .B(N6109));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4360 (.Y(N6117), .A(N8248), .B(N8217));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4363 (.Y(N6120), .A(N6709), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4370 (.Y(N6127), .A(N8222), .B(N6683));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4371 (.Y(N6138), .A(N6727), .B(N6703));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5164 (.Y(N6129), .AN(N5466), .B(N8227), .C(N8256));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5165 (.Y(N6136), .A(N4547), .B(N6117), .C(N4613));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5166 (.Y(N6139), .A(N4483), .B(N4829), .C(N6138));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5167 (.Y(N6144), .A(N6131), .B(N6129), .C(N6127));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5168 (.Y(N6142), .A(N4349), .B(N6120), .C(N4722));
NAND3XL hyperpropagate_4_1_A_I5997 (.Y(N8516), .A(N8202), .B(N6701), .C(N6136));
NOR2XL hyperpropagate_4_1_A_I5998 (.Y(N6146), .A(N6791), .B(N8516));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5282 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[58]), .A(N6139), .B(N6142), .C(N6144), .D(N6146));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4399 (.Y(N6156), .A(N8097), .B(N8115));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4402 (.Y(N6159), .A(N8183), .B(N8224));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4404 (.Y(N6480), .A(N6737), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4405 (.Y(N6162), .A(N6721), .B(N8223));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4409 (.Y(N6166), .A(N6651), .B(N6156));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4412 (.Y(N6176), .A(N8215), .B(N4976));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5171 (.Y(N6173), .AN(N6480), .B(N8203), .C(N8234));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4414 (.Y(N6171), .A(N5282), .B(N6159));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5172 (.Y(N6178), .AN(N5235), .B(N8190), .C(N8133));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4417 (.Y(N6174), .A(N6173), .B(N6162));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4418 (.Y(N6175), .A(N6166), .B(N6171));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4420 (.Y(N6177), .A(N6176), .B(N5142));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4422 (.Y(N6179), .A(N6178), .B(N6175));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5283 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[59]), .A(N6180), .B(N6177), .C(N6174), .D(N6179));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4439 (.Y(N6196), .A(N8133), .B(N8213));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5284 (.Y(N6202), .A(N8257), .B(N8147), .C(N8081), .D(N8256));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4447 (.Y(N6204), .A(N6773), .B(N5053));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4448 (.Y(N6205), .A(N6765), .B(N6751));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4451 (.Y(N6208), .A(N6781), .B(N6581));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4452 (.Y(N6209), .A(N6204), .B(N6205));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5176 (.Y(N6210), .A(N6196), .B(N6202), .C(N6206), .D(N6209));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4454 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[60]), .A(N6208), .B(N6210));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4467 (.Y(N6406), .A(N8252), .B(N8099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4470 (.Y(N6227), .A(N8165), .B(N8238));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4474 (.Y(N6231), .A(N5990), .B(N6406));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4476 (.Y(N6233), .A(N6232), .B(N6231));
NAND3XL hyperpropagate_4_1_A_I5999 (.Y(N8524), .A(N8118), .B(N8216), .C(N6233));
NOR2XL hyperpropagate_4_1_A_I6000 (.Y(N6237), .A(N8270), .B(N8524));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4481 (.Y(N6238), .A(N4327), .B(N4934));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5178 (.Y(N6240), .A(N6227), .B(N6791), .C(N5526));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5286 (.Y(N6243), .A(N6647), .B(N4613), .C(N5398), .D(N5135));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5287 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[61]), .A(N6238), .B(N6240), .C(N6243), .D(N6237));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4494 (.Y(N6252), .A(N8216), .B(N8198));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4496 (.Y(N6254), .A(N8206), .B(N6677));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4499 (.Y(N6257), .A(N8179), .B(N6681));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4503 (.Y(N6261), .A(N8243), .B(N8175));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4506 (.Y(N6264), .A(N8165), .B(N6679));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4508 (.Y(N6266), .A(N4763), .B(N5431));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4509 (.Y(N6267), .A(N6261), .B(N6252));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5182 (.Y(N6271), .A(N8257), .B(N8213), .C(N6267));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5183 (.Y(N6273), .AN(N6272), .B(N8114), .C(N6254), .D(N8223));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5184 (.Y(N6275), .A(N6779), .B(N6797), .C(N6795));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4518 (.Y(N6276), .A(N6257), .B(N6271));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4519 (.Y(N6277), .A(N6273), .B(N6264));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5288 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[62]), .A(N6266), .B(N6276), .C(N6277), .D(N6275));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4528 (.Y(N6287), .A(N8081), .B(N8134));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4534 (.Y(N6293), .A(N6697), .B(N8113));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4535 (.Y(N6294), .A(N8207), .B(N8202));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4537 (.Y(N6296), .A(N6701), .B(N8220));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4540 (.Y(N6299), .A(N6643), .B(N6287));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4542 (.Y(N6301), .A(N8261), .B(N6695));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4543 (.Y(N6302), .A(N6759), .B(N4325));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4544 (.Y(N6303), .A(N4648), .B(N6294));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4548 (.Y(N6307), .A(N6306), .B(N6302));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4549 (.Y(N6308), .A(N6303), .B(N6299));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4550 (.Y(N6309), .A(N6293), .B(N6296));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5187 (.Y(N6310), .A(N144), .B(N6655), .C(N6304), .D(N6308));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4552 (.Y(N6311), .A(N6301), .B(N6307));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5289 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[63]), .A(N4631), .B(N6309), .C(N6310), .D(N6311));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4570 (.Y(N6330), .A(N8176), .B(N8251));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4576 (.Y(N6336), .A(N8280), .B(N6330));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5189 (.Y(N6341), .AN(N6745), .B(N8183), .C(N8151));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5190 (.Y(N6345), .A(N6675), .B(N6651), .C(N6749));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4580 (.Y(N6340), .A(N4858), .B(N6791));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4584 (.Y(N6344), .A(N8313), .B(N6336));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4586 (.Y(N6346), .A(N6345), .B(N6340));
NAND3XL hyperpropagate_4_1_A_I6001 (.Y(N8532), .A(N6701), .B(N6717), .C(N4631));
NOR2XL hyperpropagate_4_1_A_I6002 (.Y(N6350), .A(N6341), .B(N8532));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4589 (.Y(N6349), .A(N6344), .B(N6346));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4591 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[64]), .A(N6350), .B(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4595 (.Y(N6356), .A(N8150), .B(N8171));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4599 (.Y(N6360), .A(N6729), .B(N6709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4604 (.Y(N6365), .A(N8144), .B(N6711));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4605 (.Y(N6366), .A(N6687), .B(N6679));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4606 (.Y(N6367), .A(N8261), .B(N8131));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4607 (.Y(N6368), .A(N6715), .B(N6703));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4608 (.Y(N6370), .A(N167), .B(N6356));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4610 (.Y(N6377), .A(N6370), .B(N6254));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4612 (.Y(N6373), .A(N6368), .B(N5402));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4613 (.Y(N6374), .A(N6365), .B(N4515));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5192 (.Y(N6383), .A(N5555), .B(N5366), .C(N5569));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4617 (.Y(N6378), .A(N6377), .B(N6367));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4618 (.Y(N6379), .A(N6366), .B(N5830));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4619 (.Y(N6380), .A(N6373), .B(N6374));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4620 (.Y(N6381), .A(N6360), .B(N6380));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5291 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[65]), .A(N6379), .B(N6383), .C(N6378), .D(N6381));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4628 (.Y(N6389), .A(N8080), .B(N8245));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4630 (.Y(N6391), .A(N8235), .B(N8203));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4634 (.Y(N6395), .A(N6709), .B(N8113));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4636 (.Y(N6397), .A(N8243), .B(N8086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4639 (.Y(N6400), .A(N6711), .B(N8156));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4642 (.Y(N6403), .A(N6391), .B(N6389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4643 (.Y(N6404), .A(N5331), .B(N6397));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5292 (.Y(N6411), .A(N8231), .B(N8133), .C(N8220), .D(N6737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4646 (.Y(N6407), .A(N6406), .B(N6403));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5195 (.Y(N6409), .A(N8143), .B(N8096), .C(N6404));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5196 (.Y(N6414), .AN(N6368), .B(N8109), .C(N8224));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4651 (.Y(N6412), .A(N6411), .B(N6395));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4652 (.Y(N6413), .A(N6400), .B(N6407));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4654 (.Y(N6415), .A(N6414), .B(N6751));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5197 (.Y(N6418), .AN(N6409), .B(N8261), .C(N6707));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4656 (.Y(N6417), .A(N6412), .B(N6413));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4658 (.Y(N6419), .A(N6418), .B(N6417));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4659 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[66]), .A(N6415), .B(N6419));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4663 (.Y(N6424), .A(N8134), .B(N8097));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5198 (.Y(N6449), .AN(N6651), .B(N8107), .C(N8203));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5199 (.Y(N6455), .A(N8172), .B(N8118), .C(N8165));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4681 (.Y(N6442), .A(N4763), .B(N6424));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4685 (.Y(N6446), .A(N5721), .B(N6196));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5201 (.Y(N6448), .A(N6482), .B(N6117), .C(N6797));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I5202 (.Y(N6453), .AN(N6446), .B(N6655), .C(N6783), .D(N5241));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4691 (.Y(N6457), .A(N5175), .B(N6448));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4693 (.Y(N6454), .A(N6453), .B(N6442));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5203 (.Y(N6459), .A(N6455), .B(N6791), .C(N6449));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4697 (.Y(N6458), .A(N6457), .B(N6454));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4699 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[67]), .A(N6459), .B(N6458));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4715 (.Y(N6485), .A(N6683), .B(N6703));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5204 (.Y(N6477), .A(N8118), .B(N8150), .C(N8288));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5205 (.Y(N6479), .AN(N5098), .B(N8152), .C(N8202));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5206 (.Y(N6483), .A(N6482), .B(N6767), .C(N6131));
NAND3XL hyperpropagate_4_1_A_I6003 (.Y(N8540), .A(N6725), .B(N8213), .C(N8086));
NOR2XL hyperpropagate_4_1_A_I6004 (.Y(N6484), .A(N8236), .B(N8540));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4725 (.Y(N6490), .A(N6485), .B(N6479));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4726 (.Y(N6487), .A(N4861), .B(N6771));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5207 (.Y(N6488), .AN(N6483), .B(N6480), .C(N6477));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5293 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[68]), .A(N6484), .B(N6490), .C(N6488), .D(N6487));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4741 (.Y(N6502), .A(N6709), .B(N8087));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5294 (.Y(N6512), .A(N8115), .B(N8150), .C(N8097), .D(N6737));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4750 (.Y(N6511), .A(N5795), .B(N6502));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4752 (.Y(N6513), .A(N6512), .B(N5106));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4755 (.Y(N6516), .A(N4945), .B(N6511));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4758 (.Y(N6519), .A(N5573), .B(N6513));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5295 (.Y(N6522), .A(N5337), .B(N4561), .C(N4326), .D(N6367));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4760 (.Y(N6521), .A(N6516), .B(N6519));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4762 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[69]), .A(N6522), .B(N6521));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4773 (.Y(N6543), .A(N6721), .B(N6725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4774 (.Y(N6536), .A(N6685), .B(N8190));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4780 (.Y(N6542), .A(N6749), .B(N6120));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4783 (.Y(N6545), .A(N6536), .B(N6781));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4785 (.Y(N6547), .A(N6546), .B(N6542));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4786 (.Y(N6548), .A(N8290), .B(N6793));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4788 (.Y(N6550), .A(N8313), .B(N6545));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I5212 (.Y(N6554), .AN(N6548), .B(N6653), .C(N6543), .D(N5629));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4791 (.Y(N6553), .A(N6547), .B(N6550));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4793 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[70]), .A(N6554), .B(N6553));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4802 (.Y(N6565), .A(N6733), .B(N8185));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4804 (.Y(N6567), .A(N6725), .B(N6717));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4808 (.Y(N6571), .A(N6735), .B(N6715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4810 (.Y(N6573), .A(N6653), .B(N5555));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4811 (.Y(N6578), .A(N6789), .B(N6565));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4814 (.Y(N6583), .A(N5220), .B(N6573));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4816 (.Y(N6579), .A(N6578), .B(N6546));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4817 (.Y(N6585), .A(N8290), .B(N6571));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4821 (.Y(N6587), .A(N6583), .B(N6579));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I5214 (.Y(N6586), .AN(N6585), .B(N6581), .C(N6567), .D(N6751));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4825 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[71]), .A(N6587), .B(N6586));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4831 (.Y(N6594), .A(N8151), .B(N6737));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4842 (.Y(N6605), .A(N6787), .B(N6594));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4843 (.Y(N6606), .A(N6773), .B(N6138));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4845 (.Y(N6608), .A(N5536), .B(N6605));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4846 (.Y(N6609), .A(N6751), .B(N6781));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5215 (.Y(N6611), .A(N6711), .B(N6717), .C(N6606));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4852 (.Y(N6615), .A(N6608), .B(N6611));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5296 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[72]), .A(N6585), .B(N6609), .C(N8313), .D(N6615));
assign inst_cellmath__195__80__2WWMM_2WWMM_out0[22] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__198_0_bdw1157874770_bdw (
	inst_cellmath__198_0_out0,
	inst_cellmath__198_0_in0,
	inst_cellmath__198_0_in1
	); /* architecture "gate_level" */ 
output [32:0] inst_cellmath__198_0_out0;
input [15:0] inst_cellmath__198_0_in0;
input [0:0] inst_cellmath__198_0_in1;
wire N102,N106,N108,N110,N112,N114,N116 
	,N118,N120,N122,N124,N126,N128,N130,N148 
	,N150,N152,N154,N156,N158,N160,N162,N164 
	,N166,N168,N170,N172,N174,N192,N194,N196 
	,N198,N200,N202,N204,N206,N208,N210,N212 
	,N214,N216,N230,N234,N236,N238,N240,N242 
	,N244,N246,N248,N250,N252,N254,N256,N270 
	,N274,N276,N278,N280,N282,N284,N286,N288 
	,N290,N292,N294,N308,N312,N314,N316,N318 
	,N320,N322,N324,N326,N328,N330,N344,N348 
	,N350,N352,N354,N356,N358,N360,N362,N364 
	,N378,N382,N384,N386,N388,N390,N392,N394 
	,N396,N410,N414,N416,N418,N420,N422,N424 
	,N426,N440,N444,N446,N448,N450,N452,N454 
	,N468,N472,N474,N476,N478,N480,N494,N498 
	,N500,N502,N504,N518,N522,N524,N526,N540 
	,N544,N546,N560,N564,N578,N598,N599,N600 
	,N601,N602,N603,N604,N605,N606,N607,N608 
	,N609,N610,N611,N612,N613,N614,N615,N616 
	,N617,N618,N619,N620,N621,N622,N623,N624 
	,N625,N626,N627,N628,N629,N630,N631,N632 
	,N633,N634,N635,N636,N637,N638,N639,N640 
	,N641,N642,N643,N644,N645,N646,N647,N648 
	,N649,N650,N651,N652,N653,N654,N655,N656 
	,N657,N658,N659,N660,N661,N662,N663,N664 
	,N665,N666,N667,N668,N669,N670,N671,N672 
	,N673,N674,N675,N676,N677,N678,N679,N680 
	,N681,N682,N683,N684,N685,N686,N687,N688 
	,N689,N690,N691,N692,N693,N694,N695,N696 
	,N697,N698,N699,N700,N701,N702,N703,N704 
	,N705,N706,N707,N708,N709,N710,N711,N712 
	,N715,N716,N717,N718,N719,N720,N721,N722 
	,N723,N724,N725,N726,N727,N728,N729,N730 
	,N731,N732,N733,N734,N735,N736,N737,N738 
	,N739,N740,N741,N742,N743,N744,N745,N746 
	,N747,N748,N749,N750,N751,N752,N753,N754 
	,N755,N756,N757,N758,N759,N760,N761,N762 
	,N763,N764,N765,N766,N767,N768,N769,N770 
	,N771,N772,N773,N774,N775,N776,N777,N778 
	,N779,N780,N781,N782,N783,N784,N785,N786 
	,N787,N788,N789,N790,N791,N792,N793,N794 
	,N795,N796,N797,N798,N799,N800,N801,N802 
	,N803,N804,N805,N806,N807,N808,N809,N810 
	,N811,N812,N813,N814,N815,N816,N817,N818 
	,N819,N820,N821,N822,N823,N824,N825,N826 
	,N829,N830,N831,N832,N833,N834,N835,N836 
	,N837,N838,N839,N840,N841,N842,N843,N844 
	,N847,N857,N865,N877,N889,N905,N921,N925 
	,N926,N945,N967,N989,N992,N995,N998,N1001 
	,N1004,N1007,N1010,N1013,N1025,N1027,N1028,N1029 
	,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037 
	,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045 
	,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053 
	,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061 
	,N1062,N1063,N1064,N1069,N1073,N1074,N1077,N1078 
	,N1081,N1082,N1085,N1086,N1089,N1090,N1093,N1094 
	,N1097,N1098,N1103,N1109,N1110,N1113,N1114,N1119 
	,N1143,N1145,N1146,N1147,N1148,N1149,N1150,N1151 
	,N1152,N1153,N1154,N1155,N1156,N1161,N1163,N1165 
	,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1181 
	,N1183,N1185,N1187,N1220,N1223,N1226,N1229,N1232 
	,N1235,N1238,N1241,N1244,N1247,N1250,N1253,N1256 
	,N1259,N1262,N1265,N1268,N1271,N1274,N1277,N1288 
	,N1289,N1291,N1292,N1294,N1295,N1297,N1298,N1300 
	,N1301,N1303,N1304,N1306,N1307,N1309,N1310,N1312 
	,N1313,N1315,N1316,N1318,N1319,N1546,N1555,N1571 
	,N1580,N1633,N1635,N1636,N1637,N1642,N1643,N1649 
	,N1654,N1658,N1659,N1660,N1661,N1662,N1664,N1665 
	,N1666,N1668,N1669,N1670,N1671,N1672,N1676,N1678 
	,N1684,N1689,N1690,N1695,N1696,N1702,N1708,N1713 
	,N1714,N1719,N1720,N1725,N1728,N1729,N1730,N1731 
	,N1732,N1733,N1734,N1735,N1736,N1737,N1743,N1744 
	,N1754,N1755,N1789,N1807,N1808,N1815,N1816,N1827 
	,N1828,N1835,N1836,N1837,N1838,N1839,N1856,N1862 
	,N1867,N1874,N1881;
BUFX2 inst_cellmath__198_0_I2436 (.Y(N1633), .A(inst_cellmath__198_0_in0[1]));
INVXL inst_cellmath__198_0_I958 (.Y(N1637), .A(N1633));
INVX2 inst_cellmath__198_0_I957 (.Y(N1636), .A(N1633));
INVX1 inst_cellmath__198_0_I956 (.Y(N1635), .A(N1633));
INVXL inst_cellmath__198_0_I964 (.Y(N1643), .A(inst_cellmath__198_0_in0[2]));
INVX1 inst_cellmath__198_0_I963 (.Y(N1642), .A(inst_cellmath__198_0_in0[2]));
INVX2 inst_cellmath__198_0_I970 (.Y(N1649), .A(inst_cellmath__198_0_in0[3]));
INVX2 inst_cellmath__198_0_I975 (.Y(N1654), .A(inst_cellmath__198_0_in0[4]));
INVXL inst_cellmath__198_0_I981 (.Y(N1660), .A(inst_cellmath__198_0_in0[5]));
INVX2 inst_cellmath__198_0_I980 (.Y(N1659), .A(inst_cellmath__198_0_in0[5]));
INVX2 inst_cellmath__198_0_I979 (.Y(N1658), .A(inst_cellmath__198_0_in0[5]));
INVX1 inst_cellmath__198_0_I982 (.Y(N1661), .A(inst_cellmath__198_0_in0[6]));
INVX2 inst_cellmath__198_0_I983 (.Y(N1662), .A(N1661));
INVXL inst_cellmath__198_0_I987 (.Y(N1666), .A(N1662));
INVX2 inst_cellmath__198_0_I986 (.Y(N1665), .A(N1662));
INVX2 inst_cellmath__198_0_I985 (.Y(N1664), .A(N1662));
BUFX3 inst_cellmath__198_0_I1289 (.Y(N1668), .A(inst_cellmath__198_0_in0[7]));
INVXL inst_cellmath__198_0_I993 (.Y(N1672), .A(N1668));
INVX1 inst_cellmath__198_0_I992 (.Y(N1671), .A(N1668));
INVX1 inst_cellmath__198_0_I991 (.Y(N1670), .A(N1668));
INVX1 inst_cellmath__198_0_I990 (.Y(N1669), .A(N1668));
INVXL inst_cellmath__198_0_I999 (.Y(N1678), .A(inst_cellmath__198_0_in0[8]));
INVX1 inst_cellmath__198_0_I997 (.Y(N1676), .A(inst_cellmath__198_0_in0[8]));
INVX1 inst_cellmath__198_0_I1005 (.Y(N1684), .A(inst_cellmath__198_0_in0[9]));
INVXL inst_cellmath__198_0_I1011 (.Y(N1690), .A(inst_cellmath__198_0_in0[10]));
INVX1 inst_cellmath__198_0_I1010 (.Y(N1689), .A(inst_cellmath__198_0_in0[10]));
INVXL inst_cellmath__198_0_I1017 (.Y(N1696), .A(inst_cellmath__198_0_in0[11]));
INVX2 inst_cellmath__198_0_I1016 (.Y(N1695), .A(inst_cellmath__198_0_in0[11]));
INVX1 inst_cellmath__198_0_I1023 (.Y(N1702), .A(inst_cellmath__198_0_in0[12]));
INVX1 inst_cellmath__198_0_I1029 (.Y(N1708), .A(inst_cellmath__198_0_in0[13]));
INVXL inst_cellmath__198_0_I1035 (.Y(N1714), .A(inst_cellmath__198_0_in0[14]));
INVX1 inst_cellmath__198_0_I1034 (.Y(N1713), .A(inst_cellmath__198_0_in0[14]));
INVXL inst_cellmath__198_0_I1041 (.Y(N1720), .A(inst_cellmath__198_0_in0[15]));
INVX1 inst_cellmath__198_0_I1040 (.Y(N1719), .A(inst_cellmath__198_0_in0[15]));
INVX1 inst_cellmath__198_0_I1046 (.Y(N1725), .A(inst_cellmath__198_0_in1[0]));
BUFX3 inst_cellmath__198_0_I1204 (.Y(N1728), .A(inst_cellmath__198_0_in0[0]));
INVXL inst_cellmath__198_0_I1053 (.Y(N1732), .A(N1728));
INVX1 inst_cellmath__198_0_I1052 (.Y(N1731), .A(N1728));
INVX1 inst_cellmath__198_0_I1051 (.Y(N1730), .A(N1728));
INVX1 inst_cellmath__198_0_I1050 (.Y(N1729), .A(N1728));
INVXL inst_cellmath__198_0_I21 (.Y(inst_cellmath__198_0_out0[0]), .A(N1732));
OR2XL inst_cellmath__198_0_I23 (.Y(N102), .A(N1729), .B(N1637));
NOR2XL inst_cellmath__198_0_I24 (.Y(N826), .A(N1732), .B(N1642));
NOR2XL inst_cellmath__198_0_I25 (.Y(N106), .A(N1731), .B(N1649));
NOR2XL inst_cellmath__198_0_I26 (.Y(N108), .A(N1731), .B(N1654));
NOR2XL inst_cellmath__198_0_I27 (.Y(N110), .A(N1731), .B(N1660));
NOR2XL inst_cellmath__198_0_I28 (.Y(N112), .A(N1731), .B(N1666));
NOR2XL inst_cellmath__198_0_I29 (.Y(N114), .A(N1731), .B(N1672));
NOR2XL inst_cellmath__198_0_I30 (.Y(N116), .A(N1730), .B(N1678));
NOR2XL inst_cellmath__198_0_I31 (.Y(N118), .A(N1730), .B(N1684));
NOR2XL inst_cellmath__198_0_I32 (.Y(N120), .A(N1730), .B(N1690));
NOR2XL inst_cellmath__198_0_I33 (.Y(N122), .A(N1730), .B(N1696));
NOR2XL inst_cellmath__198_0_I34 (.Y(N124), .A(N1730), .B(N1702));
NOR2X1 inst_cellmath__198_0_I35 (.Y(N126), .A(N1729), .B(N1708));
NOR2XL inst_cellmath__198_0_I36 (.Y(N128), .A(N1729), .B(N1714));
NOR2X1 inst_cellmath__198_0_I37 (.Y(N130), .A(N1729), .B(N1720));
OR2XL inst_cellmath__198_0_I38 (.Y(N598), .A(N1729), .B(N1725));
NOR2XL inst_cellmath__198_0_I45 (.Y(N148), .A(N1637), .B(N1642));
NOR2XL inst_cellmath__198_0_I46 (.Y(N150), .A(N1636), .B(N1649));
NOR2XL inst_cellmath__198_0_I47 (.Y(N152), .A(N1636), .B(N1654));
NOR2XL inst_cellmath__198_0_I48 (.Y(N154), .A(N1636), .B(N1660));
NOR2XL inst_cellmath__198_0_I49 (.Y(N156), .A(N1636), .B(N1666));
NOR2XL inst_cellmath__198_0_I50 (.Y(N158), .A(N1636), .B(N1672));
NOR2XL inst_cellmath__198_0_I51 (.Y(N160), .A(N1635), .B(N1678));
NOR2XL inst_cellmath__198_0_I52 (.Y(N162), .A(N1635), .B(N1684));
NOR2XL inst_cellmath__198_0_I53 (.Y(N164), .A(N1635), .B(N1690));
NOR2XL inst_cellmath__198_0_I54 (.Y(N166), .A(N1635), .B(N1696));
NOR2XL inst_cellmath__198_0_I55 (.Y(N168), .A(N1635), .B(N1702));
NOR2XL inst_cellmath__198_0_I56 (.Y(N170), .A(N1636), .B(N1708));
NOR2XL inst_cellmath__198_0_I57 (.Y(N172), .A(N1636), .B(N1714));
NOR2XL inst_cellmath__198_0_I58 (.Y(N174), .A(N1636), .B(N1720));
OR2XL inst_cellmath__198_0_I2438 (.Y(N599), .A(N1636), .B(N1725));
NOR2XL inst_cellmath__198_0_I66 (.Y(N192), .A(N1643), .B(N1649));
NOR2XL inst_cellmath__198_0_I67 (.Y(N194), .A(N1643), .B(N1654));
NOR2XL inst_cellmath__198_0_I68 (.Y(N196), .A(N1642), .B(N1659));
NOR2XL inst_cellmath__198_0_I69 (.Y(N198), .A(N1642), .B(N1665));
NOR2XL inst_cellmath__198_0_I70 (.Y(N200), .A(N1642), .B(N1671));
NOR2XL inst_cellmath__198_0_I71 (.Y(N202), .A(N1642), .B(N1678));
NOR2XL inst_cellmath__198_0_I72 (.Y(N204), .A(N1642), .B(N1684));
NOR2XL inst_cellmath__198_0_I73 (.Y(N206), .A(N1642), .B(N1689));
NOR2XL inst_cellmath__198_0_I74 (.Y(N208), .A(N1642), .B(N1695));
NOR2XL inst_cellmath__198_0_I75 (.Y(N210), .A(N1642), .B(N1702));
NOR2XL inst_cellmath__198_0_I76 (.Y(N212), .A(N1642), .B(N1708));
NOR2XL inst_cellmath__198_0_I77 (.Y(N214), .A(N1642), .B(N1713));
NOR2XL inst_cellmath__198_0_I78 (.Y(N216), .A(N1642), .B(N1719));
OR2XL inst_cellmath__198_0_I79 (.Y(N600), .A(N1643), .B(N1725));
INVXL inst_cellmath__198_0_I84 (.Y(N230), .A(N1649));
NOR2XL inst_cellmath__198_0_I86 (.Y(N234), .A(N1649), .B(N1654));
NOR2XL inst_cellmath__198_0_I87 (.Y(N236), .A(N1649), .B(N1659));
NOR2XL inst_cellmath__198_0_I88 (.Y(N238), .A(N1649), .B(N1665));
NOR2XL inst_cellmath__198_0_I89 (.Y(N240), .A(N1649), .B(N1671));
NOR2XL inst_cellmath__198_0_I90 (.Y(N242), .A(N1649), .B(N1678));
NOR2XL inst_cellmath__198_0_I91 (.Y(N244), .A(N1649), .B(N1684));
NOR2XL inst_cellmath__198_0_I92 (.Y(N246), .A(N1649), .B(N1689));
NOR2XL inst_cellmath__198_0_I93 (.Y(N248), .A(N1649), .B(N1695));
NOR2XL inst_cellmath__198_0_I94 (.Y(N250), .A(N1649), .B(N1702));
NOR2XL inst_cellmath__198_0_I95 (.Y(N252), .A(N1649), .B(N1708));
NOR2XL inst_cellmath__198_0_I96 (.Y(N254), .A(N1649), .B(N1713));
NOR2XL inst_cellmath__198_0_I97 (.Y(N256), .A(N1649), .B(N1719));
OR2XL inst_cellmath__198_0_I98 (.Y(N601), .A(N1649), .B(N1725));
INVXL inst_cellmath__198_0_I103 (.Y(N270), .A(N1654));
NOR2XL inst_cellmath__198_0_I105 (.Y(N274), .A(N1654), .B(N1659));
NOR2XL inst_cellmath__198_0_I106 (.Y(N276), .A(N1654), .B(N1665));
NOR2XL inst_cellmath__198_0_I107 (.Y(N278), .A(N1654), .B(N1671));
NOR2XL inst_cellmath__198_0_I108 (.Y(N280), .A(N1654), .B(N1678));
NOR2XL inst_cellmath__198_0_I109 (.Y(N282), .A(N1654), .B(N1684));
NOR2XL inst_cellmath__198_0_I110 (.Y(N284), .A(N1654), .B(N1689));
NOR2XL inst_cellmath__198_0_I111 (.Y(N286), .A(N1654), .B(N1695));
NOR2XL inst_cellmath__198_0_I112 (.Y(N288), .A(N1654), .B(N1702));
NOR2XL inst_cellmath__198_0_I113 (.Y(N290), .A(N1654), .B(N1708));
NOR2XL inst_cellmath__198_0_I114 (.Y(N292), .A(N1654), .B(N1713));
NOR2XL inst_cellmath__198_0_I115 (.Y(N294), .A(N1654), .B(N1719));
OR2XL inst_cellmath__198_0_I116 (.Y(N602), .A(N1654), .B(N1725));
INVXL inst_cellmath__198_0_I121 (.Y(N308), .A(N1659));
NOR2XL inst_cellmath__198_0_I123 (.Y(N312), .A(N1659), .B(N1665));
NOR2XL inst_cellmath__198_0_I124 (.Y(N314), .A(N1659), .B(N1671));
NOR2XL inst_cellmath__198_0_I125 (.Y(N316), .A(N1659), .B(N1678));
NOR2XL inst_cellmath__198_0_I126 (.Y(N318), .A(N1658), .B(N1684));
NOR2X2 inst_cellmath__198_0_I127 (.Y(N320), .A(N1658), .B(N1689));
NOR2XL inst_cellmath__198_0_I128 (.Y(N322), .A(N1658), .B(N1695));
NOR2XL inst_cellmath__198_0_I129 (.Y(N324), .A(N1658), .B(N1702));
NOR2XL inst_cellmath__198_0_I130 (.Y(N326), .A(N1658), .B(N1708));
NOR2XL inst_cellmath__198_0_I131 (.Y(N328), .A(N1659), .B(N1713));
NOR2XL inst_cellmath__198_0_I132 (.Y(N330), .A(N1659), .B(N1719));
OR2XL inst_cellmath__198_0_I133 (.Y(N603), .A(N1659), .B(N1725));
INVXL inst_cellmath__198_0_I138 (.Y(N344), .A(N1665));
NOR2XL inst_cellmath__198_0_I140 (.Y(N348), .A(N1665), .B(N1671));
NOR2XL inst_cellmath__198_0_I141 (.Y(N350), .A(N1665), .B(N1678));
NOR2XL inst_cellmath__198_0_I142 (.Y(N352), .A(N1665), .B(N1684));
NOR2XL inst_cellmath__198_0_I143 (.Y(N354), .A(N1664), .B(N1689));
NOR2X2 inst_cellmath__198_0_I144 (.Y(N356), .A(N1664), .B(N1695));
NOR2XL inst_cellmath__198_0_I145 (.Y(N358), .A(N1664), .B(N1702));
NOR2XL inst_cellmath__198_0_I146 (.Y(N360), .A(N1664), .B(N1708));
NOR2XL inst_cellmath__198_0_I147 (.Y(N362), .A(N1664), .B(N1713));
NOR2XL inst_cellmath__198_0_I148 (.Y(N364), .A(N1665), .B(N1719));
OR2XL inst_cellmath__198_0_I149 (.Y(N604), .A(N1665), .B(N1725));
INVXL inst_cellmath__198_0_I154 (.Y(N378), .A(N1669));
NOR2XL inst_cellmath__198_0_I156 (.Y(N382), .A(N1669), .B(N1676));
NOR2XL inst_cellmath__198_0_I157 (.Y(N384), .A(N1669), .B(N1684));
NOR2X1 inst_cellmath__198_0_I158 (.Y(N386), .A(N1669), .B(N1689));
NOR2XL inst_cellmath__198_0_I159 (.Y(N388), .A(N1670), .B(N1695));
NOR2XL inst_cellmath__198_0_I160 (.Y(N390), .A(N1670), .B(N1702));
NOR2XL inst_cellmath__198_0_I161 (.Y(N392), .A(N1670), .B(N1708));
NOR2XL inst_cellmath__198_0_I162 (.Y(N394), .A(N1670), .B(N1713));
NOR2XL inst_cellmath__198_0_I163 (.Y(N396), .A(N1670), .B(N1719));
OR2XL inst_cellmath__198_0_I164 (.Y(N605), .A(N1669), .B(N1725));
INVXL inst_cellmath__198_0_I169 (.Y(N410), .A(N1676));
NOR2XL inst_cellmath__198_0_I171 (.Y(N414), .A(N1676), .B(N1684));
NOR2XL inst_cellmath__198_0_I172 (.Y(N416), .A(N1676), .B(N1689));
NOR2XL inst_cellmath__198_0_I173 (.Y(N418), .A(N1676), .B(N1695));
NOR2XL inst_cellmath__198_0_I174 (.Y(N420), .A(N1676), .B(N1702));
NOR2XL inst_cellmath__198_0_I175 (.Y(N422), .A(N1676), .B(N1708));
NOR2XL inst_cellmath__198_0_I176 (.Y(N424), .A(N1676), .B(N1713));
NOR2XL inst_cellmath__198_0_I177 (.Y(N426), .A(N1676), .B(N1719));
OR2XL inst_cellmath__198_0_I178 (.Y(N606), .A(N1676), .B(N1725));
INVXL inst_cellmath__198_0_I183 (.Y(N440), .A(N1684));
NOR2XL inst_cellmath__198_0_I185 (.Y(N444), .A(N1684), .B(N1689));
NOR2XL inst_cellmath__198_0_I186 (.Y(N446), .A(N1684), .B(N1695));
NOR2XL inst_cellmath__198_0_I187 (.Y(N448), .A(N1684), .B(N1702));
NOR2XL inst_cellmath__198_0_I188 (.Y(N450), .A(N1684), .B(N1708));
NOR2XL inst_cellmath__198_0_I189 (.Y(N452), .A(N1684), .B(N1713));
NOR2XL inst_cellmath__198_0_I190 (.Y(N454), .A(N1684), .B(N1719));
OR2XL inst_cellmath__198_0_I191 (.Y(N607), .A(N1684), .B(N1725));
INVXL inst_cellmath__198_0_I196 (.Y(N468), .A(N1690));
NOR2XL inst_cellmath__198_0_I198 (.Y(N472), .A(N1690), .B(N1695));
NOR2XL inst_cellmath__198_0_I199 (.Y(N474), .A(N1690), .B(N1702));
NOR2XL inst_cellmath__198_0_I200 (.Y(N476), .A(N1690), .B(N1708));
NOR2XL inst_cellmath__198_0_I201 (.Y(N478), .A(N1689), .B(N1713));
NOR2XL inst_cellmath__198_0_I202 (.Y(N480), .A(N1689), .B(N1719));
OR2XL inst_cellmath__198_0_I203 (.Y(N608), .A(N1690), .B(N1725));
INVXL inst_cellmath__198_0_I208 (.Y(N494), .A(N1695));
NOR2XL inst_cellmath__198_0_I210 (.Y(N498), .A(N1695), .B(N1702));
NOR2XL inst_cellmath__198_0_I211 (.Y(N500), .A(N1695), .B(N1708));
NOR2XL inst_cellmath__198_0_I212 (.Y(N502), .A(N1695), .B(N1713));
NOR2XL inst_cellmath__198_0_I213 (.Y(N504), .A(N1695), .B(N1719));
OR2XL inst_cellmath__198_0_I214 (.Y(N609), .A(N1695), .B(N1725));
INVXL inst_cellmath__198_0_I219 (.Y(N518), .A(N1702));
NOR2XL inst_cellmath__198_0_I221 (.Y(N522), .A(N1702), .B(N1708));
NOR2XL inst_cellmath__198_0_I222 (.Y(N524), .A(N1702), .B(N1713));
NOR2XL inst_cellmath__198_0_I223 (.Y(N526), .A(N1702), .B(N1719));
OR2XL inst_cellmath__198_0_I224 (.Y(N610), .A(N1702), .B(N1725));
INVXL inst_cellmath__198_0_I229 (.Y(N540), .A(N1708));
NOR2XL inst_cellmath__198_0_I231 (.Y(N544), .A(N1708), .B(N1713));
NOR2XL inst_cellmath__198_0_I232 (.Y(N546), .A(N1708), .B(N1719));
OR2XL inst_cellmath__198_0_I233 (.Y(N611), .A(N1708), .B(N1725));
INVXL inst_cellmath__198_0_I238 (.Y(N560), .A(N1713));
NOR2XL inst_cellmath__198_0_I240 (.Y(N564), .A(N1713), .B(N1719));
OR2XL inst_cellmath__198_0_I241 (.Y(N612), .A(N1713), .B(N1725));
INVXL inst_cellmath__198_0_I246 (.Y(N578), .A(N1719));
ADDHX1 inst_cellmath__198_0_I269 (.CO(N614), .S(N613), .A(N106), .B(N148));
INVXL inst_cellmath__198_0_I1054 (.Y(N1733), .A(N613));
ADDHX1 inst_cellmath__198_0_I270 (.CO(N616), .S(N615), .A(N108), .B(N150));
ADDHX1 inst_cellmath__198_0_I271 (.CO(N618), .S(N617), .A(N110), .B(N152));
ADDFX1 inst_cellmath__198_0_I272 (.CO(N620), .S(N619), .A(N192), .B(N230), .CI(N616));
ADDHX1 inst_cellmath__198_0_I273 (.CO(N622), .S(N621), .A(N112), .B(N154));
ADDFX1 inst_cellmath__198_0_I274 (.CO(N624), .S(N623), .A(N618), .B(N194), .CI(N621));
ADDHX1 inst_cellmath__198_0_I275 (.CO(N626), .S(N625), .A(N114), .B(N156));
ADDFX1 inst_cellmath__198_0_I276 (.CO(N628), .S(N627), .A(N270), .B(N234), .CI(N622));
ADDFX1 inst_cellmath__198_0_I277 (.CO(N630), .S(N629), .A(N625), .B(N196), .CI(N624));
ADDHX1 inst_cellmath__198_0_I278 (.CO(N632), .S(N631), .A(N116), .B(N158));
ADDFX1 inst_cellmath__198_0_I279 (.CO(N634), .S(N633), .A(N198), .B(N236), .CI(N626));
ADDFX1 inst_cellmath__198_0_I280 (.CO(N636), .S(N635), .A(N628), .B(N631), .CI(N633));
ADDHX1 inst_cellmath__198_0_I281 (.CO(N638), .S(N637), .A(N118), .B(N160));
ADDFX1 inst_cellmath__198_0_I282 (.CO(N640), .S(N639), .A(N238), .B(N308), .CI(N274));
ADDFX1 inst_cellmath__198_0_I283 (.CO(N642), .S(N641), .A(N632), .B(N200), .CI(N637));
ADDFX1 inst_cellmath__198_0_I284 (.CO(N644), .S(N643), .A(N639), .B(N634), .CI(N641));
ADDHX1 inst_cellmath__198_0_I285 (.CO(N646), .S(N645), .A(N120), .B(N162));
ADDFX1 inst_cellmath__198_0_I286 (.CO(N648), .S(N647), .A(N276), .B(N240), .CI(N638));
ADDFX1 inst_cellmath__198_0_I287 (.CO(N650), .S(N649), .A(N645), .B(N202), .CI(N640));
ADDFX1 inst_cellmath__198_0_I288 (.CO(N652), .S(N651), .A(N647), .B(N642), .CI(N649));
ADDHX1 inst_cellmath__198_0_I289 (.CO(N654), .S(N653), .A(N344), .B(N122));
ADDFX1 inst_cellmath__198_0_I290 (.CO(N656), .S(N655), .A(N164), .B(N312), .CI(N242));
ADDFX1 inst_cellmath__198_0_I291 (.CO(N658), .S(N657), .A(N646), .B(N278), .CI(N653));
ADDFX1 inst_cellmath__198_0_I292 (.CO(N660), .S(N659), .A(N648), .B(N204), .CI(N655));
ADDFX1 inst_cellmath__198_0_I293 (.CO(N662), .S(N661), .A(N650), .B(N657), .CI(N659));
ADDHX1 inst_cellmath__198_0_I294 (.CO(N664), .S(N663), .A(N124), .B(N166));
ADDFX1 inst_cellmath__198_0_I295 (.CO(N666), .S(N665), .A(N654), .B(N314), .CI(N244));
ADDFX1 inst_cellmath__198_0_I296 (.CO(N668), .S(N667), .A(N206), .B(N280), .CI(N663));
ADDFX1 inst_cellmath__198_0_I297 (.CO(N670), .S(N669), .A(N658), .B(N656), .CI(N665));
ADDFX1 inst_cellmath__198_0_I298 (.CO(N672), .S(N671), .A(N660), .B(N667), .CI(N669));
ADDHX1 inst_cellmath__198_0_I299 (.CO(N674), .S(N673), .A(N348), .B(N126));
ADDFX1 inst_cellmath__198_0_I300 (.CO(N676), .S(N675), .A(N316), .B(N378), .CI(N168));
ADDFX1 inst_cellmath__198_0_I301 (.CO(N678), .S(N677), .A(N282), .B(N246), .CI(N664));
ADDFX1 inst_cellmath__198_0_I302 (.CO(N680), .S(N679), .A(N673), .B(N208), .CI(N666));
ADDFX1 inst_cellmath__198_0_I303 (.CO(N682), .S(N681), .A(N668), .B(N675), .CI(N677));
ADDFX1 inst_cellmath__198_0_I304 (.CO(N684), .S(N683), .A(N670), .B(N679), .CI(N681));
ADDHX1 inst_cellmath__198_0_I305 (.CO(N686), .S(N685), .A(N350), .B(N128));
ADDFX1 inst_cellmath__198_0_I306 (.CO(N688), .S(N687), .A(N170), .B(N318), .CI(N248));
ADDFX1 inst_cellmath__198_0_I307 (.CO(N690), .S(N689), .A(N284), .B(N674), .CI(N210));
ADDFX1 inst_cellmath__198_0_I308 (.CO(N692), .S(N691), .A(N676), .B(N685), .CI(N678));
ADDFX1 inst_cellmath__198_0_I309 (.CO(N694), .S(N693), .A(N689), .B(N687), .CI(N680));
ADDFHXL inst_cellmath__198_0_I310 (.CO(N696), .S(N695), .A(N691), .B(N682), .CI(N693));
ADDHX1 inst_cellmath__198_0_I311 (.CO(N698), .S(N697), .A(N352), .B(N382));
ADDFX1 inst_cellmath__198_0_I312 (.CO(N700), .S(N699), .A(N320), .B(N130), .CI(N410));
ADDFX1 inst_cellmath__198_0_I313 (.CO(N702), .S(N701), .A(N250), .B(N172), .CI(N286));
ADDFX1 inst_cellmath__198_0_I314 (.CO(N704), .S(N703), .A(N686), .B(N212), .CI(N697));
ADDFX1 inst_cellmath__198_0_I315 (.CO(N706), .S(N705), .A(N688), .B(N699), .CI(N690));
ADDFX1 inst_cellmath__198_0_I316 (.CO(N708), .S(N707), .A(N703), .B(N701), .CI(N692));
ADDFX1 inst_cellmath__198_0_I317 (.CO(N710), .S(N709), .A(N694), .B(N705), .CI(N707));
XNOR2X1 hap1_A_I894 (.Y(N711), .A(N354), .B(N384));
OR2XL hap1_A_I895 (.Y(N712), .A(N354), .B(N384));
ADDFX1 inst_cellmath__198_0_I319 (.CO(N716), .S(N715), .A(N174), .B(N322), .CI(N598));
ADDFX1 inst_cellmath__198_0_I320 (.CO(N718), .S(N717), .A(N698), .B(N252), .CI(N288));
ADDFX1 inst_cellmath__198_0_I321 (.CO(N720), .S(N719), .A(N711), .B(N214), .CI(N700));
ADDFX1 inst_cellmath__198_0_I322 (.CO(N722), .S(N721), .A(N715), .B(N702), .CI(N704));
ADDFHXL inst_cellmath__198_0_I323 (.CO(N724), .S(N723), .A(N719), .B(N717), .CI(N706));
ADDFHXL inst_cellmath__198_0_I324 (.CO(N726), .S(N725), .A(N708), .B(N721), .CI(N723));
ADDFX1 inst_cellmath__198_0_I325 (.CO(N728), .S(N727), .A(N356), .B(N440), .CI(N386));
ADDFX1 inst_cellmath__198_0_I326 (.CO(N730), .S(N729), .A(N414), .B(N324), .CI(N599));
ADDFX1 inst_cellmath__198_0_I327 (.CO(N732), .S(N731), .A(N254), .B(N712), .CI(N290));
ADDFHXL inst_cellmath__198_0_I328 (.CO(N734), .S(N733), .A(N716), .B(N216), .CI(N727));
ADDFX1 inst_cellmath__198_0_I329 (.CO(N736), .S(N735), .A(N729), .B(N718), .CI(N720));
ADDFXL inst_cellmath__198_0_I330 (.CO(N738), .S(N737), .A(N733), .B(N731), .CI(N722));
ADDFHX1 inst_cellmath__198_0_I331 (.CO(N740), .S(N739), .A(N724), .B(N735), .CI(N737));
ADDFX1 inst_cellmath__198_0_I332 (.CO(N742), .S(N741), .A(N358), .B(N388), .CI(N326));
ADDFX1 inst_cellmath__198_0_I333 (.CO(N744), .S(N743), .A(N256), .B(N416), .CI(N292));
ADDFX1 inst_cellmath__198_0_I334 (.CO(N746), .S(N745), .A(N728), .B(N600), .CI(N730));
ADDFX1 inst_cellmath__198_0_I335 (.CO(N748), .S(N747), .A(N732), .B(N741), .CI(N743));
ADDFHXL inst_cellmath__198_0_I336 (.CO(N750), .S(N749), .A(N745), .B(N734), .CI(N736));
ADDFHXL inst_cellmath__198_0_I337 (.CO(N752), .S(N751), .A(N738), .B(N747), .CI(N749));
ADDFX1 inst_cellmath__198_0_I338 (.CO(N754), .S(N753), .A(N444), .B(N468), .CI(N390));
ADDFX1 inst_cellmath__198_0_I339 (.CO(N756), .S(N755), .A(N418), .B(N360), .CI(N328));
ADDFX1 inst_cellmath__198_0_I340 (.CO(N758), .S(N757), .A(N601), .B(N294), .CI(N742));
ADDFX1 inst_cellmath__198_0_I341 (.CO(N760), .S(N759), .A(N744), .B(N753), .CI(N755));
ADDFX1 inst_cellmath__198_0_I342 (.CO(N762), .S(N761), .A(N757), .B(N746), .CI(N748));
ADDFHX1 inst_cellmath__198_0_I343 (.CO(N764), .S(N763), .A(N750), .B(N759), .CI(N761));
ADDFX1 inst_cellmath__198_0_I344 (.CO(N766), .S(N765), .A(N392), .B(N446), .CI(N330));
ADDFX1 inst_cellmath__198_0_I345 (.CO(N768), .S(N767), .A(N362), .B(N420), .CI(N602));
ADDFX1 inst_cellmath__198_0_I346 (.CO(N770), .S(N769), .A(N756), .B(N754), .CI(N765));
ADDFX1 inst_cellmath__198_0_I347 (.CO(N772), .S(N771), .A(N758), .B(N767), .CI(N760));
ADDFX1 inst_cellmath__198_0_I348 (.CO(N774), .S(N773), .A(N762), .B(N769), .CI(N771));
ADDFX1 inst_cellmath__198_0_I349 (.CO(N776), .S(N775), .A(N472), .B(N494), .CI(N364));
ADDFX1 inst_cellmath__198_0_I350 (.CO(N778), .S(N777), .A(N422), .B(N448), .CI(N603));
ADDFX1 inst_cellmath__198_0_I351 (.CO(N780), .S(N779), .A(N766), .B(N394), .CI(N775));
ADDFX1 inst_cellmath__198_0_I352 (.CO(N782), .S(N781), .A(N777), .B(N768), .CI(N770));
ADDFX1 inst_cellmath__198_0_I353 (.CO(N784), .S(N783), .A(N772), .B(N779), .CI(N781));
ADDFX1 inst_cellmath__198_0_I354 (.CO(N786), .S(N785), .A(N474), .B(N396), .CI(N450));
ADDFX1 inst_cellmath__198_0_I355 (.CO(N788), .S(N787), .A(N424), .B(N604), .CI(N776));
ADDFX1 inst_cellmath__198_0_I356 (.CO(N790), .S(N789), .A(N785), .B(N778), .CI(N780));
ADDFX1 inst_cellmath__198_0_I357 (.CO(N792), .S(N791), .A(N782), .B(N787), .CI(N789));
ADDFX1 inst_cellmath__198_0_I358 (.CO(N794), .S(N793), .A(N498), .B(N518), .CI(N476));
ADDFX1 inst_cellmath__198_0_I359 (.CO(N796), .S(N795), .A(N605), .B(N426), .CI(N452));
ADDFX1 inst_cellmath__198_0_I360 (.CO(N798), .S(N797), .A(N793), .B(N786), .CI(N788));
ADDFX1 inst_cellmath__198_0_I361 (.CO(N800), .S(N799), .A(N790), .B(N795), .CI(N797));
ADDFX1 inst_cellmath__198_0_I362 (.CO(N802), .S(N801), .A(N500), .B(N454), .CI(N478));
ADDFX1 inst_cellmath__198_0_I363 (.CO(N804), .S(N803), .A(N794), .B(N606), .CI(N796));
ADDFX1 inst_cellmath__198_0_I364 (.CO(N806), .S(N805), .A(N798), .B(N801), .CI(N803));
ADDFX1 inst_cellmath__198_0_I365 (.CO(N808), .S(N807), .A(N480), .B(N540), .CI(N522));
ADDFX1 inst_cellmath__198_0_I366 (.CO(N810), .S(N809), .A(N502), .B(N607), .CI(N802));
ADDFX1 inst_cellmath__198_0_I367 (.CO(N812), .S(N811), .A(N804), .B(N807), .CI(N809));
ADDFX1 inst_cellmath__198_0_I368 (.CO(N814), .S(N813), .A(N608), .B(N504), .CI(N524));
ADDFX1 inst_cellmath__198_0_I369 (.CO(N816), .S(N815), .A(N813), .B(N808), .CI(N810));
ADDFX1 inst_cellmath__198_0_I370 (.CO(N818), .S(N817), .A(N560), .B(N526), .CI(N609));
ADDFX1 inst_cellmath__198_0_I371 (.CO(N820), .S(N819), .A(N814), .B(N544), .CI(N817));
ADDFX1 inst_cellmath__198_0_I372 (.CO(N822), .S(N821), .A(N610), .B(N546), .CI(N818));
ADDFX1 inst_cellmath__198_0_I373 (.CO(N824), .S(N823), .A(N564), .B(N578), .CI(N611));
NOR2XL inst_cellmath__198_0_I374 (.Y(N825), .A(N102), .B(N1636));
NOR2XL inst_cellmath__198_0_I378 (.Y(N829), .A(N614), .B(N615));
NAND2XL inst_cellmath__198_0_I379 (.Y(N830), .A(N614), .B(N615));
NOR2XL inst_cellmath__198_0_I380 (.Y(N831), .A(N617), .B(N619));
NAND2XL inst_cellmath__198_0_I381 (.Y(N832), .A(N617), .B(N619));
NOR2XL inst_cellmath__198_0_I382 (.Y(N833), .A(N620), .B(N623));
NAND2XL inst_cellmath__198_0_I383 (.Y(N834), .A(N620), .B(N623));
NOR2XL inst_cellmath__198_0_I384 (.Y(N835), .A(N627), .B(N629));
NAND2XL inst_cellmath__198_0_I385 (.Y(N836), .A(N627), .B(N629));
NOR2XL inst_cellmath__198_0_I386 (.Y(N837), .A(N630), .B(N635));
NAND2X1 inst_cellmath__198_0_I387 (.Y(N838), .A(N630), .B(N635));
NOR2X1 inst_cellmath__198_0_I388 (.Y(N839), .A(N636), .B(N643));
NAND2XL inst_cellmath__198_0_I389 (.Y(N840), .A(N636), .B(N643));
NOR2X1 inst_cellmath__198_0_I390 (.Y(N841), .A(N644), .B(N651));
NAND2X2 inst_cellmath__198_0_I391 (.Y(N842), .A(N644), .B(N651));
NOR2XL inst_cellmath__198_0_I392 (.Y(N843), .A(N652), .B(N661));
NAND2XL inst_cellmath__198_0_I393 (.Y(N844), .A(N652), .B(N661));
AND2XL inst_cellmath__198_0_I396 (.Y(N847), .A(N826), .B(N825));
AND2XL inst_cellmath__198_0_I1205 (.Y(N1734), .A(N1642), .B(N1733));
INVXL inst_cellmath__198_0_I1056 (.Y(N1735), .A(N1734));
OR2XL inst_cellmath__198_0_I1206 (.Y(N1736), .A(N1642), .B(N1733));
INVXL inst_cellmath__198_0_I1058 (.Y(N1737), .A(N1736));
OAI21X1 inst_cellmath__198_0_I404 (.Y(N857), .A0(N1737), .A1(N847), .B0(N1735));
AOI21X1 inst_cellmath__198_0_I412 (.Y(N865), .A0(N830), .A1(N857), .B0(N829));
INVXL inst_cellmath__198_0_I1064 (.Y(N1743), .A(N831));
INVXL inst_cellmath__198_0_I1065 (.Y(N1744), .A(N832));
OAI21X1 inst_cellmath__198_0_I424 (.Y(N877), .A0(N1744), .A1(N865), .B0(N1743));
AOI21X2 inst_cellmath__198_0_I436 (.Y(N889), .A0(N834), .A1(N877), .B0(N833));
INVXL inst_cellmath__198_0_I1075 (.Y(N1754), .A(N835));
INVXL inst_cellmath__198_0_I1076 (.Y(N1755), .A(N836));
OAI21X2 inst_cellmath__198_0_I452 (.Y(N905), .A0(N1755), .A1(N889), .B0(N1754));
AOI21X2 inst_cellmath__198_0_I468 (.Y(N921), .A0(N838), .A1(N905), .B0(N837));
AOI21X2 inst_cellmath__198_0_I472 (.Y(N925), .A0(N842), .A1(N839), .B0(N841));
NAND2X1 inst_cellmath__198_0_I473 (.Y(N926), .A(N842), .B(N840));
OAI21X2 inst_cellmath__198_0_I492 (.Y(N945), .A0(N926), .A1(N921), .B0(N925));
NOR2BX1 andori2bb1_A_I2439 (.Y(N1867), .AN(N840), .B(N921));
NOR2XL andori2bb1_A_I1309 (.Y(N1789), .A(N1867), .B(N839));
AOI21X2 inst_cellmath__198_0_I514 (.Y(N967), .A0(N844), .A1(N945), .B0(N843));
NAND2BXL inst_cellmath__198_0_I534 (.Y(N989), .AN(N1734), .B(N1736));
NAND2BXL inst_cellmath__198_0_I537 (.Y(N992), .AN(N829), .B(N830));
NAND2BXL inst_cellmath__198_0_I540 (.Y(N995), .AN(N831), .B(N832));
NAND2BXL inst_cellmath__198_0_I543 (.Y(N998), .AN(N833), .B(N834));
NAND2BXL inst_cellmath__198_0_I546 (.Y(N1001), .AN(N835), .B(N836));
NAND2BXL inst_cellmath__198_0_I549 (.Y(N1004), .AN(N837), .B(N838));
NAND2BXL inst_cellmath__198_0_I552 (.Y(N1007), .AN(N839), .B(N840));
NAND2BXL inst_cellmath__198_0_I555 (.Y(N1010), .AN(N841), .B(N842));
NAND2BXL inst_cellmath__198_0_I558 (.Y(N1013), .AN(N843), .B(N844));
XOR2XL inst_cellmath__198_0_I559 (.Y(inst_cellmath__198_0_out0[2]), .A(N102), .B(N1637));
XOR2XL inst_cellmath__198_0_I1209 (.Y(inst_cellmath__198_0_out0[3]), .A(N825), .B(N826));
XNOR2X1 inst_cellmath__198_0_I561 (.Y(inst_cellmath__198_0_out0[4]), .A(N847), .B(N989));
XOR2XL inst_cellmath__198_0_I1210 (.Y(inst_cellmath__198_0_out0[5]), .A(N857), .B(N992));
XNOR2X1 inst_cellmath__198_0_I563 (.Y(inst_cellmath__198_0_out0[6]), .A(N865), .B(N995));
XOR2XL inst_cellmath__198_0_I1211 (.Y(inst_cellmath__198_0_out0[7]), .A(N877), .B(N998));
XNOR2X1 inst_cellmath__198_0_I565 (.Y(inst_cellmath__198_0_out0[8]), .A(N889), .B(N1001));
XOR2XL inst_cellmath__198_0_I1212 (.Y(inst_cellmath__198_0_out0[9]), .A(N905), .B(N1004));
XNOR2X1 inst_cellmath__198_0_I567 (.Y(inst_cellmath__198_0_out0[10]), .A(N921), .B(N1007));
XNOR2X1 inst_cellmath__198_0_I568 (.Y(inst_cellmath__198_0_out0[11]), .A(N1789), .B(N1010));
XOR2XL inst_cellmath__198_0_I1213 (.Y(inst_cellmath__198_0_out0[12]), .A(N945), .B(N1013));
INVX2 inst_cellmath__198_0_I570 (.Y(N1025), .A(N967));
NOR2XL inst_cellmath__198_0_I571 (.Y(N1027), .A(N662), .B(N671));
NAND2X1 inst_cellmath__198_0_I572 (.Y(N1028), .A(N662), .B(N671));
NOR2X1 inst_cellmath__198_0_I573 (.Y(N1029), .A(N672), .B(N683));
NAND2XL inst_cellmath__198_0_I574 (.Y(N1030), .A(N672), .B(N683));
NOR2X1 inst_cellmath__198_0_I575 (.Y(N1031), .A(N684), .B(N695));
NAND2X2 inst_cellmath__198_0_I576 (.Y(N1032), .A(N684), .B(N695));
NOR2X2 inst_cellmath__198_0_I577 (.Y(N1033), .A(N696), .B(N709));
NAND2X2 inst_cellmath__198_0_I578 (.Y(N1034), .A(N696), .B(N709));
NOR2X1 inst_cellmath__198_0_I579 (.Y(N1035), .A(N710), .B(N725));
NAND2X4 inst_cellmath__198_0_I580 (.Y(N1036), .A(N710), .B(N725));
NOR2X2 inst_cellmath__198_0_I581 (.Y(N1037), .A(N726), .B(N739));
NAND2X2 inst_cellmath__198_0_I582 (.Y(N1038), .A(N726), .B(N739));
NOR2X1 inst_cellmath__198_0_I583 (.Y(N1039), .A(N740), .B(N751));
NAND2X4 inst_cellmath__198_0_I584 (.Y(N1040), .A(N740), .B(N751));
NOR2X2 inst_cellmath__198_0_I585 (.Y(N1041), .A(N752), .B(N763));
NAND2X2 inst_cellmath__198_0_I586 (.Y(N1042), .A(N752), .B(N763));
NOR2X1 inst_cellmath__198_0_I587 (.Y(N1043), .A(N764), .B(N773));
NAND2X4 inst_cellmath__198_0_I588 (.Y(N1044), .A(N764), .B(N773));
NOR2X1 inst_cellmath__198_0_I589 (.Y(N1045), .A(N774), .B(N783));
NAND2X2 inst_cellmath__198_0_I590 (.Y(N1046), .A(N774), .B(N783));
NOR2XL inst_cellmath__198_0_I591 (.Y(N1047), .A(N784), .B(N791));
NAND2X2 inst_cellmath__198_0_I592 (.Y(N1048), .A(N784), .B(N791));
NOR2X1 inst_cellmath__198_0_I593 (.Y(N1049), .A(N792), .B(N799));
NAND2XL inst_cellmath__198_0_I594 (.Y(N1050), .A(N792), .B(N799));
NOR2XL inst_cellmath__198_0_I595 (.Y(N1051), .A(N805), .B(N800));
NAND2XL inst_cellmath__198_0_I596 (.Y(N1052), .A(N805), .B(N800));
NOR2XL inst_cellmath__198_0_I597 (.Y(N1053), .A(N806), .B(N811));
NAND2XL inst_cellmath__198_0_I598 (.Y(N1054), .A(N806), .B(N811));
NOR2XL inst_cellmath__198_0_I599 (.Y(N1055), .A(N812), .B(N815));
NAND2XL inst_cellmath__198_0_I600 (.Y(N1056), .A(N812), .B(N815));
NOR2XL inst_cellmath__198_0_I601 (.Y(N1057), .A(N819), .B(N816));
NAND2XL inst_cellmath__198_0_I602 (.Y(N1058), .A(N819), .B(N816));
NOR2XL inst_cellmath__198_0_I603 (.Y(N1059), .A(N820), .B(N821));
NAND2XL inst_cellmath__198_0_I604 (.Y(N1060), .A(N820), .B(N821));
NOR2XL inst_cellmath__198_0_I605 (.Y(N1061), .A(N823), .B(N822));
NAND2XL inst_cellmath__198_0_I606 (.Y(N1062), .A(N823), .B(N822));
NOR2XL inst_cellmath__198_0_I607 (.Y(N1063), .A(N612), .B(N824));
NAND2XL inst_cellmath__198_0_I608 (.Y(N1064), .A(N612), .B(N824));
AOI21X4 inst_cellmath__198_0_I613 (.Y(N1069), .A0(N1028), .A1(N1025), .B0(N1027));
AOI21X4 inst_cellmath__198_0_I617 (.Y(N1073), .A0(N1032), .A1(N1029), .B0(N1031));
NAND2X2 inst_cellmath__198_0_I618 (.Y(N1074), .A(N1032), .B(N1030));
AOI21X4 inst_cellmath__198_0_I621 (.Y(N1077), .A0(N1036), .A1(N1033), .B0(N1035));
NAND2X4 inst_cellmath__198_0_I622 (.Y(N1078), .A(N1036), .B(N1034));
AOI21X4 inst_cellmath__198_0_I625 (.Y(N1081), .A0(N1040), .A1(N1037), .B0(N1039));
NAND2X4 inst_cellmath__198_0_I626 (.Y(N1082), .A(N1040), .B(N1038));
AOI21X4 inst_cellmath__198_0_I629 (.Y(N1085), .A0(N1044), .A1(N1041), .B0(N1043));
NAND2X4 inst_cellmath__198_0_I630 (.Y(N1086), .A(N1044), .B(N1042));
AOI21X2 inst_cellmath__198_0_I633 (.Y(N1089), .A0(N1048), .A1(N1045), .B0(N1047));
NAND2X2 inst_cellmath__198_0_I634 (.Y(N1090), .A(N1048), .B(N1046));
AOI21X1 inst_cellmath__198_0_I637 (.Y(N1093), .A0(N1052), .A1(N1049), .B0(N1051));
NAND2XL inst_cellmath__198_0_I638 (.Y(N1094), .A(N1052), .B(N1050));
INVXL inst_cellmath__198_0_I1128 (.Y(N1807), .A(N1053));
INVXL inst_cellmath__198_0_I1129 (.Y(N1808), .A(N1054));
AOI21XL inst_cellmath__198_0_I641 (.Y(N1097), .A0(N1056), .A1(N1053), .B0(N1055));
NAND2XL inst_cellmath__198_0_I642 (.Y(N1098), .A(N1056), .B(N1054));
OAI21XL inst_cellmath__198_0_I647 (.Y(N1103), .A0(N1808), .A1(N1093), .B0(N1807));
AOI21XL inst_cellmath__198_0_I653 (.Y(N1109), .A0(N1060), .A1(N1057), .B0(N1059));
NAND2XL inst_cellmath__198_0_I654 (.Y(N1110), .A(N1060), .B(N1058));
INVXL inst_cellmath__198_0_I1136 (.Y(N1815), .A(N1061));
INVXL inst_cellmath__198_0_I1137 (.Y(N1816), .A(N1062));
AOI21XL inst_cellmath__198_0_I657 (.Y(N1113), .A0(N1064), .A1(N1061), .B0(N1063));
NAND2XL inst_cellmath__198_0_I658 (.Y(N1114), .A(N1064), .B(N1062));
OAI21XL inst_cellmath__198_0_I663 (.Y(N1119), .A0(N1816), .A1(N1109), .B0(N1815));
OA21X1 inst_cellmath__198_0_I1296 (.Y(N1827), .A0(N1098), .A1(N1093), .B0(N1097));
OR2XL inst_cellmath__198_0_I1241 (.Y(N1828), .A(N1098), .B(N1094));
OA21X1 inst_cellmath__198_0_I1217 (.Y(N1835), .A0(N1114), .A1(N1109), .B0(N1113));
OR2XL inst_cellmath__198_0_I1218 (.Y(N1836), .A(N1114), .B(N1110));
INVX1 inst_cellmath__198_0_I1158 (.Y(N1837), .A(N1069));
OAI21X2 inst_cellmath__198_0_I687 (.Y(N1143), .A0(N1074), .A1(N1069), .B0(N1073));
OAI21X2 inst_cellmath__198_0_I689 (.Y(N1145), .A0(N1078), .A1(N1073), .B0(N1077));
NOR2X1 inst_cellmath__198_0_I690 (.Y(N1146), .A(N1078), .B(N1074));
OAI21X4 inst_cellmath__198_0_I691 (.Y(N1147), .A0(N1082), .A1(N1077), .B0(N1081));
NOR2X1 inst_cellmath__198_0_I692 (.Y(N1148), .A(N1082), .B(N1078));
OAI21X2 inst_cellmath__198_0_I693 (.Y(N1149), .A0(N1086), .A1(N1081), .B0(N1085));
NOR2X2 inst_cellmath__198_0_I694 (.Y(N1150), .A(N1086), .B(N1082));
OAI21X2 inst_cellmath__198_0_I695 (.Y(N1151), .A0(N1090), .A1(N1085), .B0(N1089));
NOR2X2 inst_cellmath__198_0_I696 (.Y(N1152), .A(N1090), .B(N1086));
OAI21XL inst_cellmath__198_0_I697 (.Y(N1153), .A0(N1828), .A1(N1089), .B0(N1827));
NOR2XL inst_cellmath__198_0_I698 (.Y(N1154), .A(N1828), .B(N1090));
OAI21XL inst_cellmath__198_0_I699 (.Y(N1155), .A0(N1836), .A1(N1827), .B0(N1835));
NOR2XL inst_cellmath__198_0_I700 (.Y(N1156), .A(N1836), .B(N1828));
INVXL inst_cellmath__198_0_I1159 (.Y(N1838), .A(N1837));
INVX2 inst_cellmath__198_0_I1160 (.Y(N1839), .A(N1143));
AOI21X2 inst_cellmath__198_0_I705 (.Y(N1161), .A0(N1146), .A1(N1837), .B0(N1145));
AOI21X2 inst_cellmath__198_0_I707 (.Y(N1163), .A0(N1148), .A1(N1143), .B0(N1147));
AOI21X2 inst_cellmath__198_0_I709 (.Y(N1165), .A0(N1150), .A1(N1145), .B0(N1149));
NAND2X1 inst_cellmath__198_0_I710 (.Y(N1166), .A(N1150), .B(N1146));
AOI21X4 inst_cellmath__198_0_I711 (.Y(N1167), .A0(N1152), .A1(N1147), .B0(N1151));
NAND2X2 inst_cellmath__198_0_I712 (.Y(N1168), .A(N1152), .B(N1148));
AOI21X1 inst_cellmath__198_0_I713 (.Y(N1169), .A0(N1154), .A1(N1149), .B0(N1153));
NAND2XL inst_cellmath__198_0_I714 (.Y(N1170), .A(N1154), .B(N1150));
AOI21X1 inst_cellmath__198_0_I715 (.Y(N1171), .A0(N1156), .A1(N1151), .B0(N1155));
NAND2XL inst_cellmath__198_0_I716 (.Y(N1172), .A(N1156), .B(N1152));
OAI21X2 inst_cellmath__198_0_I725 (.Y(N1181), .A0(N1166), .A1(N1838), .B0(N1165));
OAI21X4 inst_cellmath__198_0_I727 (.Y(N1183), .A0(N1168), .A1(N1839), .B0(N1167));
OAI21X2 inst_cellmath__198_0_I729 (.Y(N1185), .A0(N1170), .A1(N1161), .B0(N1169));
OAI21X1 inst_cellmath__198_0_I731 (.Y(N1187), .A0(N1172), .A1(N1163), .B0(N1171));
INVXL inst_cellmath__198_0_I1177 (.Y(N1856), .A(N1093));
INVXL inst_cellmath__198_0_I1183 (.Y(N1862), .A(N1109));
NAND2BXL inst_cellmath__198_0_I764 (.Y(N1220), .AN(N1027), .B(N1028));
NAND2BXL inst_cellmath__198_0_I767 (.Y(N1223), .AN(N1029), .B(N1030));
NAND2BXL inst_cellmath__198_0_I770 (.Y(N1226), .AN(N1031), .B(N1032));
NAND2BXL inst_cellmath__198_0_I773 (.Y(N1229), .AN(N1033), .B(N1034));
NAND2BXL inst_cellmath__198_0_I776 (.Y(N1232), .AN(N1035), .B(N1036));
NAND2BXL inst_cellmath__198_0_I779 (.Y(N1235), .AN(N1037), .B(N1038));
NAND2BXL inst_cellmath__198_0_I782 (.Y(N1238), .AN(N1039), .B(N1040));
NAND2BXL inst_cellmath__198_0_I785 (.Y(N1241), .AN(N1041), .B(N1042));
NAND2BXL inst_cellmath__198_0_I788 (.Y(N1244), .AN(N1043), .B(N1044));
NAND2BXL inst_cellmath__198_0_I791 (.Y(N1247), .AN(N1045), .B(N1046));
NAND2BXL inst_cellmath__198_0_I794 (.Y(N1250), .AN(N1047), .B(N1048));
NAND2BXL inst_cellmath__198_0_I797 (.Y(N1253), .AN(N1049), .B(N1050));
NAND2BXL inst_cellmath__198_0_I800 (.Y(N1256), .AN(N1051), .B(N1052));
NAND2BXL inst_cellmath__198_0_I803 (.Y(N1259), .AN(N1053), .B(N1054));
NAND2BXL inst_cellmath__198_0_I806 (.Y(N1262), .AN(N1055), .B(N1056));
NAND2BXL inst_cellmath__198_0_I809 (.Y(N1265), .AN(N1057), .B(N1058));
NAND2BXL inst_cellmath__198_0_I812 (.Y(N1268), .AN(N1059), .B(N1060));
NAND2BXL inst_cellmath__198_0_I815 (.Y(N1271), .AN(N1061), .B(N1062));
NAND2BXL inst_cellmath__198_0_I818 (.Y(N1274), .AN(N1063), .B(N1064));
AND2XL inst_cellmath__198_0_I1270 (.Y(N1277), .A(N1719), .B(inst_cellmath__198_0_in1[0]));
XOR2XL inst_cellmath__198_0_I1220 (.Y(inst_cellmath__198_0_out0[13]), .A(N1025), .B(N1220));
XNOR2X1 inst_cellmath__198_0_I824 (.Y(inst_cellmath__198_0_out0[14]), .A(N1838), .B(N1223));
XNOR2X1 inst_cellmath__198_0_I825 (.Y(inst_cellmath__198_0_out0[16]), .A(N1839), .B(N1229));
XNOR2X1 inst_cellmath__198_0_I826 (.Y(inst_cellmath__198_0_out0[18]), .A(N1161), .B(N1235));
XNOR2X1 inst_cellmath__198_0_I1221 (.Y(inst_cellmath__198_0_out0[20]), .A(N1163), .B(N1241));
XOR2XL inst_cellmath__198_0_I828 (.Y(inst_cellmath__198_0_out0[22]), .A(N1181), .B(N1247));
XOR2XL inst_cellmath__198_0_I829 (.Y(inst_cellmath__198_0_out0[24]), .A(N1183), .B(N1253));
XOR2XL inst_cellmath__198_0_I830 (.Y(inst_cellmath__198_0_out0[28]), .A(N1185), .B(N1265));
XOR2XL inst_cellmath__198_0_I2441 (.Y(inst_cellmath__198_0_out0[32]), .A(N1187), .B(N1277));
XNOR2X1 node_cs_reduced_local_A_I900 (.Y(N1288), .A(N1226), .B(N1030));
XNOR2X1 node_cs_reduced_local_A_I901 (.Y(N1289), .A(N1226), .B(N1029));
MXI2XL inst_cellmath__198_0_I833 (.Y(inst_cellmath__198_0_out0[15]), .A(N1288), .B(N1289), .S0(N1838));
XNOR2X1 node_cs_reduced_local_A_I902 (.Y(N1291), .A(N1232), .B(N1034));
XNOR2X1 node_cs_reduced_local_A_I903 (.Y(N1292), .A(N1232), .B(N1033));
MXI2XL inst_cellmath__198_0_I835 (.Y(inst_cellmath__198_0_out0[17]), .A(N1291), .B(N1292), .S0(N1839));
XNOR2X1 node_cs_reduced_local_A_I904 (.Y(N1294), .A(N1238), .B(N1038));
XNOR2X1 node_cs_reduced_local_A_I905 (.Y(N1295), .A(N1238), .B(N1037));
MXI2X1 inst_cellmath__198_0_I837 (.Y(inst_cellmath__198_0_out0[19]), .A(N1294), .B(N1295), .S0(N1161));
XNOR2X1 node_cs_reduced_local_A_I906 (.Y(N1297), .A(N1244), .B(N1042));
XNOR2X1 node_cs_reduced_local_A_I907 (.Y(N1298), .A(N1244), .B(N1041));
MXI2XL inst_cellmath__198_0_I839 (.Y(inst_cellmath__198_0_out0[21]), .A(N1297), .B(N1298), .S0(N1163));
XNOR2X1 node_cs_reduced_local_A_I908 (.Y(N1300), .A(N1250), .B(N1046));
XNOR2X1 node_cs_reduced_local_A_I909 (.Y(N1301), .A(N1250), .B(N1045));
MXI2XL inst_cellmath__198_0_I841 (.Y(inst_cellmath__198_0_out0[23]), .A(N1301), .B(N1300), .S0(N1181));
XNOR2X1 node_cs_reduced_local_A_I910 (.Y(N1303), .A(N1256), .B(N1050));
XNOR2X1 node_cs_reduced_local_A_I911 (.Y(N1304), .A(N1256), .B(N1049));
MXI2XL inst_cellmath__198_0_I843 (.Y(inst_cellmath__198_0_out0[25]), .A(N1304), .B(N1303), .S0(N1183));
XNOR2X1 node_cs_local_A_I912 (.Y(N1306), .A(N1259), .B(N1856));
NOR2BX1 node_cs_local_A_I1223 (.Y(N1546), .AN(N1094), .B(N1856));
XOR2XL node_cs_local_A_I914 (.Y(N1307), .A(N1259), .B(N1546));
MXI2XL inst_cellmath__198_0_I845 (.Y(inst_cellmath__198_0_out0[26]), .A(N1306), .B(N1307), .S0(N1183));
XNOR2X1 node_cs_local_A_I915 (.Y(N1309), .A(N1262), .B(N1103));
NOR2XL andori2bb1_A_I1310 (.Y(N1874), .A(N1808), .B(N1094));
NOR2XL andori2bb1_A_I1311 (.Y(N1555), .A(N1874), .B(N1103));
XOR2XL node_cs_local_A_I917 (.Y(N1310), .A(N1262), .B(N1555));
MXI2XL inst_cellmath__198_0_I847 (.Y(inst_cellmath__198_0_out0[27]), .A(N1309), .B(N1310), .S0(N1183));
XNOR2X1 node_cs_reduced_local_A_I918 (.Y(N1312), .A(N1268), .B(N1058));
XNOR2X1 node_cs_reduced_local_A_I919 (.Y(N1313), .A(N1268), .B(N1057));
MXI2X1 inst_cellmath__198_0_I849 (.Y(inst_cellmath__198_0_out0[29]), .A(N1313), .B(N1312), .S0(N1185));
XNOR2X1 node_cs_local_A_I920 (.Y(N1315), .A(N1271), .B(N1862));
NOR2BX1 node_cs_local_A_I1225 (.Y(N1571), .AN(N1110), .B(N1862));
XOR2XL node_cs_local_A_I922 (.Y(N1316), .A(N1271), .B(N1571));
MXI2XL inst_cellmath__198_0_I851 (.Y(inst_cellmath__198_0_out0[30]), .A(N1315), .B(N1316), .S0(N1185));
XNOR2X1 node_cs_local_A_I923 (.Y(N1318), .A(N1274), .B(N1119));
NOR2XL andori2bb1_A_I1312 (.Y(N1881), .A(N1816), .B(N1110));
NOR2XL andori2bb1_A_I1313 (.Y(N1580), .A(N1881), .B(N1119));
XOR2XL node_cs_local_A_I925 (.Y(N1319), .A(N1274), .B(N1580));
MXI2XL inst_cellmath__198_0_I853 (.Y(inst_cellmath__198_0_out0[31]), .A(N1318), .B(N1319), .S0(N1185));
assign inst_cellmath__198_0_out0[1] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__203_0_bdw1157874770_bdw (
	inst_cellmath__203_0_out0,
	inst_cellmath__203_0_out1,
	inst_cellmath__203_0_in0,
	inst_cellmath__203_0_in1,
	inst_cellmath__203_0_in2,
	inst_cellmath__203_0_in3,
	inst_cellmath__203_0_in4
	); /* architecture "gate_level" */ 
output [46:0] inst_cellmath__203_0_out0,
	inst_cellmath__203_0_out1;
input [15:0] inst_cellmath__203_0_in0;
input [32:17] inst_cellmath__203_0_in1;
input [42:23] inst_cellmath__203_0_in2;
input [21:0] inst_cellmath__203_0_in3;
input [0:0] inst_cellmath__203_0_in4;
wire N518,N520,N522,N524,N526,N528,N530 
	,N532,N534,N536,N538,N540,N542,N544,N546 
	,N548,N550,N552,N554,N560,N567,N568,N569 
	,N570,N571,N572,N573,N574,N575,N576,N577 
	,N578,N579,N580,N581,N582,N583,N584,N585 
	,N591,N596,N597,N598,N599,N600,N601,N602 
	,N603,N604,N605,N606,N607,N608,N609,N610 
	,N611,N612,N613,N614,N615,N621,N625,N626 
	,N627,N628,N629,N630,N631,N632,N633,N634 
	,N635,N636,N637,N638,N639,N640,N641,N642 
	,N643,N644,N645,N651,N655,N656,N657,N658 
	,N659,N660,N661,N662,N663,N664,N665,N666 
	,N667,N668,N669,N670,N671,N672,N673,N674 
	,N675,N681,N685,N686,N687,N688,N689,N690 
	,N691,N692,N693,N694,N695,N696,N697,N698 
	,N699,N700,N701,N702,N703,N704,N705,N711 
	,N715,N716,N717,N718,N719,N720,N721,N722 
	,N723,N724,N725,N726,N727,N728,N729,N730 
	,N731,N732,N733,N734,N735,N741,N745,N746 
	,N747,N748,N749,N750,N751,N752,N753,N754 
	,N755,N756,N757,N758,N759,N760,N761,N762 
	,N763,N764,N765,N768,N770,N779,N781,N783 
	,N785,N787,N789,N791,N793,N795,N797,N799 
	,N801,N803,N805,N807,N809,N811,N813,N815 
	,N817,N819,N1025,N1027,N1029,N1031,N1033,N1035 
	,N1037,N1039,N1041,N1043,N1045,N1047,N1049,N1051 
	,N1053,N1055,N1059,N1061,N1067,N1077,N1078,N1079 
	,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087 
	,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095 
	,N1096,N1097,N1098,N1099,N1103,N1105,N1109,N1110 
	,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118 
	,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126 
	,N1127,N1128,N1129,N1130,N1131,N1135,N1137,N1141 
	,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149 
	,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157 
	,N1158,N1159,N1160,N1161,N1162,N1163,N1167,N1169 
	,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180 
	,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188 
	,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1199 
	,N1201,N1205,N1206,N1207,N1208,N1209,N1210,N1211 
	,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219 
	,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227 
	,N1231,N1233,N1237,N1238,N1239,N1240,N1241,N1242 
	,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250 
	,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258 
	,N1259,N1263,N1265,N1269,N1270,N1271,N1272,N1273 
	,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281 
	,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289 
	,N1290,N1295,N1297,N1301,N1302,N1303,N1304,N1305 
	,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313 
	,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321 
	,N1322,N1366,N1376,N1378,N1379,N1380,N1382,N1384 
	,N1386,N1387,N1388,N1389,N1390,N1392,N1395,N1396 
	,N1397,N1398,N1399,N1400,N1403,N1404,N1405,N1406 
	,N1407,N1408,N1409,N1410,N1411,N1412,N1415,N1416 
	,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424 
	,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434 
	,N1435,N1436,N1437,N1438,N1439,N1440,N1443,N1444 
	,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452 
	,N1453,N1454,N1455,N1456,N1459,N1460,N1461,N1462 
	,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470 
	,N1471,N1472,N1473,N1474,N1475,N1476,N1479,N1480 
	,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488 
	,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496 
	,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506 
	,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514 
	,N1515,N1516,N1517,N1518,N1519,N1520,N1523,N1524 
	,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532 
	,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540 
	,N1541,N1542,N1543,N1544,N1547,N1548,N1549,N1550 
	,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558 
	,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566 
	,N1567,N1568,N1569,N1570,N1571,N1572,N1575,N1576 
	,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584 
	,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592 
	,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600 
	,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610 
	,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618 
	,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626 
	,N1627,N1628,N1629,N1630,N1633,N1634,N1635,N1636 
	,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644 
	,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652 
	,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660 
	,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670 
	,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678 
	,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686 
	,N1687,N1688,N1689,N1690,N1691,N1692,N1695,N1696 
	,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706 
	,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714 
	,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722 
	,N1723,N1724,N1725,N1726,N1729,N1730,N1732,N1733 
	,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741 
	,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749 
	,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757 
	,N1758,N1759,N1760,N1763,N1764,N1765,N1766,N1767 
	,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775 
	,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783 
	,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791 
	,N1792,N1795,N1796,N1798,N1799,N1800,N1801,N1802 
	,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810 
	,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818 
	,N1819,N1820,N1821,N1822,N1823,N1824,N1827,N1828 
	,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837 
	,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845 
	,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853 
	,N1854,N1855,N1856,N1859,N1860,N1863,N1864,N1865 
	,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873 
	,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881 
	,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1891 
	,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899 
	,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907 
	,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915 
	,N1916,N1919,N1920,N1923,N1924,N1925,N1926,N1927 
	,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935 
	,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943 
	,N1944,N1947,N1948,N1951,N1952,N1953,N1954,N1955 
	,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963 
	,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1973 
	,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981 
	,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989 
	,N1990,N1991,N1992,N1995,N1996,N1999,N2000,N2001 
	,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009 
	,N2010,N2011,N2012,N2013,N2014,N2017,N2018,N2019 
	,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027 
	,N2028,N2029,N2030,N2031,N2032,N2035,N2036,N2039 
	,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047 
	,N2048,N2049,N2050,N2053,N2054,N2055,N2056,N2057 
	,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2067 
	,N2068,N2071,N2072,N2073,N2074,N2075,N2076,N2077 
	,N2078,N2081,N2082,N2083,N2084,N2085,N2086,N2087 
	,N2088,N2091,N2092,N2095,N2096,N2097,N2098,N2101 
	,N2102,N2103,N2104,N2107,N2108,N2111,N2112,N2234 
	,N2243,N2252,N2261,N2270,N2279,N2288,N2297,N2306 
	,N2315,N2324,N2333,N2342,N2351,N2360,N2369,N2378 
	,N2387,N2396,N2405,N2414,N2423,N2425,N2436,N2445 
	,N2454,N2463,N2472,N2481,N2490,N2499,N2508,N2517 
	,N2526,N2535,N2544,N2553,N2562,N2571,N2580,N2589 
	,N2598,N2607,N2616,N2625,N2627,N2638,N2647,N2656 
	,N2665,N2674,N2683,N2692,N2701,N2710,N2719,N2728 
	,N2737,N2746,N2755,N2764,N2773,N2782,N2791,N2800 
	,N2809,N2818,N2827,N2829,N2840,N2849,N2858,N2867 
	,N2876,N2885,N2894,N2903,N2912,N2921,N2930,N2939 
	,N2948,N2957,N2966,N2975,N2984,N2993,N3002,N3011 
	,N3020,N3029,N3031,N3042,N3051,N3060,N3069,N3078 
	,N3087,N3096,N3105,N3114,N3123,N3132,N3141,N3150 
	,N3159,N3168,N3177,N3186,N3195,N3204,N3213,N3222 
	,N3231,N3233,N3244,N3253,N3262,N3271,N3280,N3289 
	,N3298,N3307,N3316,N3325,N3334,N3343,N3352,N3361 
	,N3370,N3379,N3388,N3397,N3406,N3415,N3424,N3433 
	,N3435,N3446,N3455,N3464,N3473,N3482,N3491,N3500 
	,N3509,N3518,N3527,N3536,N3545,N3554,N3563,N3572 
	,N3581,N3590,N3599,N3608,N3617,N3626,N3648,N3657 
	,N3666,N3675,N3684,N3693,N3702,N3711,N3720,N3729 
	,N3738,N3747,N3756,N3765,N3774,N3783,N3792,N3801 
	,N3810,N3819,N3828,N3837,N3846,N3855,N3857,N3868 
	,N3877,N3886,N3895,N3904,N3913,N3922,N3931,N3940 
	,N3949,N3958,N3967,N3976,N3985,N3994,N4003,N4012 
	,N4021,N4030,N4039,N4048,N4057,N4066,N4075,N4077 
	,N4088,N4097,N4106,N4115,N4124,N4133,N4142,N4151 
	,N4160,N4169,N4178,N4187,N4196,N4205,N4214,N4223 
	,N4232,N4241,N4250,N4259,N4268,N4277,N4286,N4295 
	,N4297,N4308,N4317,N4326,N4335,N4344,N4353,N4362 
	,N4371,N4380,N4389,N4398,N4407,N4416,N4425,N4434 
	,N4443,N4452,N4461,N4470,N4479,N4488,N4497,N4506 
	,N4515,N4517,N4528,N4537,N4546,N4555,N4564,N4573 
	,N4582,N4591,N4600,N4609,N4618,N4627,N4636,N4645 
	,N4654,N4663,N4672,N4681,N4690,N4699,N4708,N4717 
	,N4726,N4735,N4737,N4748,N4757,N4766,N4775,N4784 
	,N4793,N4802,N4811,N4820,N4829,N4838,N4847,N4856 
	,N4865,N4874,N4883,N4892,N4901,N4910,N4919,N4928 
	,N4937,N4946,N4955,N4957,N4968,N4977,N4986,N4995 
	,N5004,N5013,N5022,N5031,N5040,N5049,N5058,N5067 
	,N5076,N5085,N5094,N5103,N5112,N5121,N5130,N5139 
	,N5148,N5157,N5166,N5175,N5177,N5188,N5197,N5206 
	,N5215,N5224,N5233,N5242,N5251,N5260,N5269,N5278 
	,N5287,N5296,N5305,N5314,N5323,N5332,N5341,N5350 
	,N5359,N5368,N5377,N5386,N5395,N5413,N5422,N5443 
	,N5452,N5461,N5470,N5479,N5627,N5628,N5629,N5630 
	,N5631,N5632,N5633,N5634,N5635,N5636,N5637,N5638 
	,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646 
	,N5654,N5662,N5670,N5671,N5674,N5678,N5687,N5688 
	,N5691,N5696,N5705,N5706,N5707,N5711,N5712,N5720 
	,N5721,N5722,N5727,N5728,N5736,N5737,N5738,N5742 
	,N5751,N5752,N5753,N5758,N5759,N5767,N5768,N5769 
	,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777 
	,N5778,N5779,N5780,N5781,N5782,N5783,N5784,N5785 
	,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793 
	,N5794,N5804,N5820,N5839,N5848,N5865,N5874,N5891 
	,N5900,N5917,N5926,N5941,N5949,N5966,N5974,N5989 
	;
INVXL inst_cellmath__203_0_I1822 (.Y(N5627), .A(inst_cellmath__203_0_in2[23]));
INVXL inst_cellmath__203_0_I1823 (.Y(N5628), .A(inst_cellmath__203_0_in2[24]));
INVXL inst_cellmath__203_0_I1824 (.Y(N5629), .A(inst_cellmath__203_0_in2[25]));
INVXL inst_cellmath__203_0_I1825 (.Y(N5630), .A(inst_cellmath__203_0_in2[26]));
INVXL inst_cellmath__203_0_I1826 (.Y(N5631), .A(inst_cellmath__203_0_in2[27]));
INVXL inst_cellmath__203_0_I1827 (.Y(N5632), .A(inst_cellmath__203_0_in2[28]));
INVXL inst_cellmath__203_0_I1828 (.Y(N5633), .A(inst_cellmath__203_0_in2[29]));
INVXL inst_cellmath__203_0_I1829 (.Y(N5634), .A(inst_cellmath__203_0_in2[30]));
INVXL inst_cellmath__203_0_I1830 (.Y(N5635), .A(inst_cellmath__203_0_in2[31]));
INVXL inst_cellmath__203_0_I1831 (.Y(N5636), .A(inst_cellmath__203_0_in2[32]));
INVXL inst_cellmath__203_0_I1832 (.Y(N5637), .A(inst_cellmath__203_0_in2[33]));
INVXL inst_cellmath__203_0_I1833 (.Y(N5638), .A(inst_cellmath__203_0_in2[34]));
INVXL inst_cellmath__203_0_I1834 (.Y(N5639), .A(inst_cellmath__203_0_in2[35]));
INVXL inst_cellmath__203_0_I1835 (.Y(N5640), .A(inst_cellmath__203_0_in2[36]));
INVXL inst_cellmath__203_0_I1836 (.Y(N5641), .A(inst_cellmath__203_0_in2[37]));
INVXL inst_cellmath__203_0_I1837 (.Y(N5642), .A(inst_cellmath__203_0_in2[38]));
INVXL inst_cellmath__203_0_I1838 (.Y(N5643), .A(inst_cellmath__203_0_in2[39]));
INVXL inst_cellmath__203_0_I1839 (.Y(N5644), .A(inst_cellmath__203_0_in2[40]));
INVXL inst_cellmath__203_0_I1840 (.Y(N5645), .A(inst_cellmath__203_0_in2[41]));
INVXL inst_cellmath__203_0_I1841 (.Y(N5646), .A(inst_cellmath__203_0_in2[42]));
INVXL inst_cellmath__203_0_I1849 (.Y(N5654), .A(inst_cellmath__203_0_in1[17]));
NOR2XL inst_cellmath__203_0_I71 (.Y(inst_cellmath__203_0_out1[0]), .A(N5654), .B(N5627));
NOR2XL inst_cellmath__203_0_I72 (.Y(N518), .A(N5654), .B(N5628));
NOR2XL inst_cellmath__203_0_I73 (.Y(N520), .A(N5654), .B(N5629));
NOR2XL inst_cellmath__203_0_I74 (.Y(N522), .A(N5654), .B(N5630));
NOR2XL inst_cellmath__203_0_I75 (.Y(N524), .A(N5654), .B(N5631));
NOR2XL inst_cellmath__203_0_I76 (.Y(N526), .A(N5654), .B(N5632));
NOR2XL inst_cellmath__203_0_I77 (.Y(N528), .A(N5654), .B(N5633));
NOR2XL inst_cellmath__203_0_I78 (.Y(N530), .A(N5654), .B(N5634));
NOR2XL inst_cellmath__203_0_I79 (.Y(N532), .A(N5654), .B(N5635));
NOR2XL inst_cellmath__203_0_I80 (.Y(N534), .A(N5654), .B(N5636));
NOR2XL inst_cellmath__203_0_I81 (.Y(N536), .A(N5654), .B(N5637));
NOR2XL inst_cellmath__203_0_I82 (.Y(N538), .A(N5654), .B(N5638));
NOR2XL inst_cellmath__203_0_I83 (.Y(N540), .A(N5654), .B(N5639));
NOR2XL inst_cellmath__203_0_I84 (.Y(N542), .A(N5654), .B(N5640));
NOR2XL inst_cellmath__203_0_I85 (.Y(N544), .A(N5654), .B(N5641));
NOR2XL inst_cellmath__203_0_I86 (.Y(N546), .A(N5654), .B(N5642));
NOR2XL inst_cellmath__203_0_I87 (.Y(N548), .A(N5654), .B(N5643));
NOR2XL inst_cellmath__203_0_I88 (.Y(N550), .A(N5654), .B(N5644));
NOR2XL inst_cellmath__203_0_I89 (.Y(N552), .A(N5654), .B(N5645));
NOR2XL inst_cellmath__203_0_I90 (.Y(N554), .A(N5654), .B(N5646));
NOR2BX1 inst_cellmath__203_0_I1821 (.Y(N560), .AN(inst_cellmath__203_0_in1[18]), .B(inst_cellmath__203_0_in1[19]));
INVXL inst_cellmath__203_0_I1857 (.Y(N5662), .A(inst_cellmath__203_0_in1[18]));
INVXL inst_cellmath__203_0_I1865 (.Y(N5670), .A(N560));
INVXL inst_cellmath__203_0_I1866 (.Y(N5671), .A(inst_cellmath__203_0_in1[19]));
NOR2XL addgen2_A_I1063 (.Y(N2234), .A(N5627), .B(N5662));
MXI2XL addgen2_A_I1064 (.Y(inst_cellmath__203_0_out0[1]), .A(N5671), .B(N5670), .S0(N2234));
MXI2XL inst_cellmath__203_0_I1065 (.Y(N2243), .A(N5628), .B(N5627), .S0(N5662));
MXI2XL inst_cellmath__203_0_I4809 (.Y(inst_cellmath__203_0_out1[2]), .A(N5671), .B(N5670), .S0(N2243));
MXI2XL addgen2_A_I1067 (.Y(N2252), .A(N5629), .B(N5628), .S0(N5662));
MXI2XL addgen2_A_I1068 (.Y(N567), .A(N5671), .B(N5670), .S0(N2252));
MXI2XL addgen2_A_I1069 (.Y(N2261), .A(N5630), .B(N5629), .S0(N5662));
MXI2XL addgen2_A_I1070 (.Y(N568), .A(N5671), .B(N5670), .S0(N2261));
MXI2XL addgen2_A_I1071 (.Y(N2270), .A(N5631), .B(N5630), .S0(N5662));
MXI2XL addgen2_A_I1072 (.Y(N569), .A(N5671), .B(N5670), .S0(N2270));
MXI2XL addgen2_A_I1073 (.Y(N2279), .A(N5632), .B(N5631), .S0(N5662));
MXI2XL addgen2_A_I1074 (.Y(N570), .A(N5671), .B(N5670), .S0(N2279));
MXI2XL addgen2_A_I1075 (.Y(N2288), .A(N5633), .B(N5632), .S0(N5662));
MXI2XL addgen2_A_I1076 (.Y(N571), .A(N5671), .B(N5670), .S0(N2288));
MXI2XL addgen2_A_I1077 (.Y(N2297), .A(N5634), .B(N5633), .S0(N5662));
MXI2XL addgen2_A_I1078 (.Y(N572), .A(N5671), .B(N5670), .S0(N2297));
MXI2XL addgen2_A_I1079 (.Y(N2306), .A(N5635), .B(N5634), .S0(N5662));
MXI2XL addgen2_A_I1080 (.Y(N573), .A(N5671), .B(N5670), .S0(N2306));
MXI2XL addgen2_A_I1081 (.Y(N2315), .A(N5636), .B(N5635), .S0(N5662));
MXI2XL addgen2_A_I1082 (.Y(N574), .A(N5671), .B(N5670), .S0(N2315));
MXI2XL addgen2_A_I1083 (.Y(N2324), .A(N5637), .B(N5636), .S0(N5662));
MXI2XL addgen2_A_I1084 (.Y(N575), .A(N5671), .B(N5670), .S0(N2324));
MXI2XL addgen2_A_I1085 (.Y(N2333), .A(N5638), .B(N5637), .S0(N5662));
MXI2XL addgen2_A_I1086 (.Y(N576), .A(N5671), .B(N5670), .S0(N2333));
MXI2XL addgen2_A_I1087 (.Y(N2342), .A(N5639), .B(N5638), .S0(N5662));
MXI2XL addgen2_A_I1088 (.Y(N577), .A(N5671), .B(N5670), .S0(N2342));
MXI2XL addgen2_A_I1089 (.Y(N2351), .A(N5640), .B(N5639), .S0(N5662));
MXI2XL addgen2_A_I1090 (.Y(N578), .A(N5671), .B(N5670), .S0(N2351));
MXI2XL addgen2_A_I1091 (.Y(N2360), .A(N5641), .B(N5640), .S0(N5662));
MXI2XL addgen2_A_I1092 (.Y(N579), .A(N5671), .B(N5670), .S0(N2360));
MXI2XL addgen2_A_I1093 (.Y(N2369), .A(N5642), .B(N5641), .S0(N5662));
MXI2XL addgen2_A_I1094 (.Y(N580), .A(N5671), .B(N5670), .S0(N2369));
MXI2XL addgen2_A_I1095 (.Y(N2378), .A(N5643), .B(N5642), .S0(N5662));
MXI2XL addgen2_A_I1096 (.Y(N581), .A(N5671), .B(N5670), .S0(N2378));
MXI2XL addgen2_A_I1097 (.Y(N2387), .A(N5644), .B(N5643), .S0(N5662));
MXI2XL addgen2_A_I1098 (.Y(N582), .A(N5671), .B(N5670), .S0(N2387));
MXI2XL addgen2_A_I1099 (.Y(N2396), .A(N5645), .B(N5644), .S0(N5662));
MXI2XL addgen2_A_I1100 (.Y(N583), .A(N5671), .B(N5670), .S0(N2396));
MXI2XL addgen2_A_I1101 (.Y(N2405), .A(N5646), .B(N5645), .S0(N5662));
MXI2XL addgen2_A_I1102 (.Y(N584), .A(N5671), .B(N5670), .S0(N2405));
NAND2XL addgen2_A_I1103 (.Y(N2414), .A(N5646), .B(N5662));
MXI2XL addgen2_A_I1104 (.Y(N585), .A(N5671), .B(N5670), .S0(N2414));
NAND2XL enc2_A_I1106 (.Y(N2423), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
NOR2XL enc2_A_I1107 (.Y(N2425), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
AND2XL enc2_A_I1108 (.Y(N591), .A(N2423), .B(inst_cellmath__203_0_in1[21]));
XOR2XL inst_cellmath__203_0_I2195 (.Y(N5674), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
INVX1 inst_cellmath__203_0_I1873 (.Y(N5678), .A(N5674));
OR2XL inst_cellmath__203_0_I4810 (.Y(N5687), .A(N2425), .B(inst_cellmath__203_0_in1[21]));
INVXL inst_cellmath__203_0_I1883 (.Y(N5688), .A(N591));
NOR2XL inst_cellmath__203_0_I1110 (.Y(N2436), .A(N5627), .B(N5678));
MXI2XL inst_cellmath__203_0_I4811 (.Y(inst_cellmath__203_0_out1[3]), .A(N5688), .B(N5687), .S0(N2436));
MXI2XL addgen2_A_I2202 (.Y(N2445), .A(N5627), .B(N5628), .S0(N5674));
MXI2XL addgen2_A_I1113 (.Y(N596), .A(N5688), .B(N5687), .S0(N2445));
MXI2XL addgen2_A_I1114 (.Y(N2454), .A(N5629), .B(N5628), .S0(N5678));
MXI2XL addgen2_A_I1115 (.Y(N597), .A(N5688), .B(N5687), .S0(N2454));
MXI2XL addgen2_A_I1116 (.Y(N2463), .A(N5630), .B(N5629), .S0(N5678));
MXI2XL addgen2_A_I1117 (.Y(N598), .A(N5688), .B(N5687), .S0(N2463));
MXI2XL addgen2_A_I1118 (.Y(N2472), .A(N5631), .B(N5630), .S0(N5678));
MXI2XL addgen2_A_I1119 (.Y(N599), .A(N5688), .B(N5687), .S0(N2472));
MXI2XL addgen2_A_I1120 (.Y(N2481), .A(N5632), .B(N5631), .S0(N5678));
MXI2XL addgen2_A_I1121 (.Y(N600), .A(N5688), .B(N5687), .S0(N2481));
MXI2XL addgen2_A_I1122 (.Y(N2490), .A(N5633), .B(N5632), .S0(N5678));
MXI2XL addgen2_A_I1123 (.Y(N601), .A(N5688), .B(N5687), .S0(N2490));
MXI2XL addgen2_A_I1124 (.Y(N2499), .A(N5634), .B(N5633), .S0(N5678));
MXI2XL addgen2_A_I1125 (.Y(N602), .A(N5688), .B(N5687), .S0(N2499));
MXI2XL addgen2_A_I1126 (.Y(N2508), .A(N5635), .B(N5634), .S0(N5678));
MXI2XL addgen2_A_I1127 (.Y(N603), .A(N5688), .B(N5687), .S0(N2508));
MXI2XL addgen2_A_I1128 (.Y(N2517), .A(N5636), .B(N5635), .S0(N5678));
MXI2XL addgen2_A_I1129 (.Y(N604), .A(N5688), .B(N5687), .S0(N2517));
MXI2XL addgen2_A_I1130 (.Y(N2526), .A(N5637), .B(N5636), .S0(N5678));
MXI2XL addgen2_A_I1131 (.Y(N605), .A(N5688), .B(N5687), .S0(N2526));
MXI2XL addgen2_A_I1132 (.Y(N2535), .A(N5638), .B(N5637), .S0(N5678));
MXI2XL addgen2_A_I1133 (.Y(N606), .A(N5688), .B(N5687), .S0(N2535));
MXI2XL addgen2_A_I1134 (.Y(N2544), .A(N5639), .B(N5638), .S0(N5678));
MXI2XL addgen2_A_I1135 (.Y(N607), .A(N5688), .B(N5687), .S0(N2544));
MXI2XL addgen2_A_I1136 (.Y(N2553), .A(N5640), .B(N5639), .S0(N5678));
MXI2XL addgen2_A_I1137 (.Y(N608), .A(N5688), .B(N5687), .S0(N2553));
MXI2XL addgen2_A_I1138 (.Y(N2562), .A(N5641), .B(N5640), .S0(N5678));
MXI2XL addgen2_A_I1139 (.Y(N609), .A(N5688), .B(N5687), .S0(N2562));
MXI2XL addgen2_A_I1140 (.Y(N2571), .A(N5642), .B(N5641), .S0(N5678));
MXI2XL addgen2_A_I1141 (.Y(N610), .A(N5688), .B(N5687), .S0(N2571));
MXI2XL addgen2_A_I1142 (.Y(N2580), .A(N5643), .B(N5642), .S0(N5678));
MXI2XL addgen2_A_I1143 (.Y(N611), .A(N5688), .B(N5687), .S0(N2580));
MXI2XL addgen2_A_I1144 (.Y(N2589), .A(N5644), .B(N5643), .S0(N5678));
MXI2XL addgen2_A_I1145 (.Y(N612), .A(N5688), .B(N5687), .S0(N2589));
MXI2XL addgen2_A_I1146 (.Y(N2598), .A(N5645), .B(N5644), .S0(N5678));
MXI2XL addgen2_A_I1147 (.Y(N613), .A(N5688), .B(N5687), .S0(N2598));
MXI2XL addgen2_A_I1148 (.Y(N2607), .A(N5646), .B(N5645), .S0(N5678));
MXI2XL addgen2_A_I1149 (.Y(N614), .A(N5688), .B(N5687), .S0(N2607));
NAND2XL addgen2_A_I1150 (.Y(N2616), .A(N5646), .B(N5678));
MXI2XL addgen2_A_I1151 (.Y(N615), .A(N5688), .B(N5687), .S0(N2616));
NAND2XL enc2_A_I1153 (.Y(N2625), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
NOR2XL enc2_A_I1154 (.Y(N2627), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
AND2XL enc2_A_I1155 (.Y(N621), .A(N2625), .B(inst_cellmath__203_0_in1[23]));
XOR2XL inst_cellmath__203_0_I2203 (.Y(N5691), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
INVX1 inst_cellmath__203_0_I1891 (.Y(N5696), .A(N5691));
OR2XL inst_cellmath__203_0_I4812 (.Y(N5705), .A(N2627), .B(inst_cellmath__203_0_in1[23]));
INVXL inst_cellmath__203_0_I1901 (.Y(N5706), .A(N621));
NOR2XL addgen2_A_I1157 (.Y(N2638), .A(N5627), .B(N5696));
MXI2XL addgen2_A_I1158 (.Y(N625), .A(N5706), .B(N5705), .S0(N2638));
MXI2XL addgen2_A_I2204 (.Y(N2647), .A(N5627), .B(N5628), .S0(N5691));
MXI2XL addgen2_A_I1160 (.Y(N626), .A(N5706), .B(N5705), .S0(N2647));
MXI2XL addgen2_A_I1161 (.Y(N2656), .A(N5629), .B(N5628), .S0(N5696));
MXI2XL addgen2_A_I1162 (.Y(N627), .A(N5706), .B(N5705), .S0(N2656));
MXI2XL addgen2_A_I1163 (.Y(N2665), .A(N5630), .B(N5629), .S0(N5696));
MXI2XL addgen2_A_I1164 (.Y(N628), .A(N5706), .B(N5705), .S0(N2665));
MXI2XL addgen2_A_I1165 (.Y(N2674), .A(N5631), .B(N5630), .S0(N5696));
MXI2XL addgen2_A_I1166 (.Y(N629), .A(N5706), .B(N5705), .S0(N2674));
MXI2XL addgen2_A_I1167 (.Y(N2683), .A(N5632), .B(N5631), .S0(N5696));
MXI2XL addgen2_A_I1168 (.Y(N630), .A(N5706), .B(N5705), .S0(N2683));
MXI2XL addgen2_A_I1169 (.Y(N2692), .A(N5633), .B(N5632), .S0(N5696));
MXI2XL addgen2_A_I1170 (.Y(N631), .A(N5706), .B(N5705), .S0(N2692));
MXI2XL addgen2_A_I1171 (.Y(N2701), .A(N5634), .B(N5633), .S0(N5696));
MXI2XL addgen2_A_I1172 (.Y(N632), .A(N5706), .B(N5705), .S0(N2701));
MXI2XL addgen2_A_I1173 (.Y(N2710), .A(N5635), .B(N5634), .S0(N5696));
MXI2XL addgen2_A_I1174 (.Y(N633), .A(N5706), .B(N5705), .S0(N2710));
MXI2XL addgen2_A_I1175 (.Y(N2719), .A(N5636), .B(N5635), .S0(N5696));
MXI2XL addgen2_A_I1176 (.Y(N634), .A(N5706), .B(N5705), .S0(N2719));
MXI2XL addgen2_A_I1177 (.Y(N2728), .A(N5637), .B(N5636), .S0(N5696));
MXI2XL addgen2_A_I1178 (.Y(N635), .A(N5706), .B(N5705), .S0(N2728));
MXI2XL addgen2_A_I1179 (.Y(N2737), .A(N5638), .B(N5637), .S0(N5696));
MXI2XL addgen2_A_I1180 (.Y(N636), .A(N5706), .B(N5705), .S0(N2737));
MXI2XL addgen2_A_I1181 (.Y(N2746), .A(N5639), .B(N5638), .S0(N5696));
MXI2XL addgen2_A_I1182 (.Y(N637), .A(N5706), .B(N5705), .S0(N2746));
MXI2XL addgen2_A_I1183 (.Y(N2755), .A(N5640), .B(N5639), .S0(N5696));
MXI2XL addgen2_A_I1184 (.Y(N638), .A(N5706), .B(N5705), .S0(N2755));
MXI2XL addgen2_A_I1185 (.Y(N2764), .A(N5641), .B(N5640), .S0(N5696));
MXI2XL addgen2_A_I1186 (.Y(N639), .A(N5706), .B(N5705), .S0(N2764));
MXI2XL addgen2_A_I1187 (.Y(N2773), .A(N5642), .B(N5641), .S0(N5696));
MXI2XL addgen2_A_I1188 (.Y(N640), .A(N5706), .B(N5705), .S0(N2773));
MXI2XL addgen2_A_I1189 (.Y(N2782), .A(N5643), .B(N5642), .S0(N5696));
MXI2XL addgen2_A_I1190 (.Y(N641), .A(N5706), .B(N5705), .S0(N2782));
MXI2XL addgen2_A_I1191 (.Y(N2791), .A(N5644), .B(N5643), .S0(N5696));
MXI2XL addgen2_A_I1192 (.Y(N642), .A(N5706), .B(N5705), .S0(N2791));
MXI2XL addgen2_A_I1193 (.Y(N2800), .A(N5645), .B(N5644), .S0(N5696));
MXI2XL addgen2_A_I1194 (.Y(N643), .A(N5706), .B(N5705), .S0(N2800));
MXI2XL addgen2_A_I1195 (.Y(N2809), .A(N5646), .B(N5645), .S0(N5696));
MXI2XL addgen2_A_I1196 (.Y(N644), .A(N5706), .B(N5705), .S0(N2809));
NAND2XL addgen2_A_I1197 (.Y(N2818), .A(N5646), .B(N5696));
MXI2XL addgen2_A_I1198 (.Y(N645), .A(N5706), .B(N5705), .S0(N2818));
NAND2XL enc2_A_I1200 (.Y(N2827), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
NOR2XL enc2_A_I1201 (.Y(N2829), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
AND2XL enc2_A_I1202 (.Y(N651), .A(N2827), .B(inst_cellmath__203_0_in1[25]));
XOR2XL inst_cellmath__203_0_I2205 (.Y(N5707), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
INVXL inst_cellmath__203_0_I1907 (.Y(N5712), .A(N5707));
INVXL inst_cellmath__203_0_I1906 (.Y(N5711), .A(N5707));
OR2XL inst_cellmath__203_0_I4813 (.Y(N5720), .A(N2829), .B(inst_cellmath__203_0_in1[25]));
INVXL inst_cellmath__203_0_I1916 (.Y(N5721), .A(N651));
NOR2XL addgen2_A_I1204 (.Y(N2840), .A(N5627), .B(N5712));
MXI2XL addgen2_A_I1205 (.Y(N655), .A(N5721), .B(N5720), .S0(N2840));
MXI2XL addgen2_A_I1206 (.Y(N2849), .A(N5628), .B(N5627), .S0(N5712));
MXI2XL addgen2_A_I1207 (.Y(N656), .A(N5721), .B(N5720), .S0(N2849));
MXI2XL addgen2_A_I1208 (.Y(N2858), .A(N5629), .B(N5628), .S0(N5711));
MXI2XL addgen2_A_I1209 (.Y(N657), .A(N5721), .B(N5720), .S0(N2858));
MXI2XL addgen2_A_I1210 (.Y(N2867), .A(N5630), .B(N5629), .S0(N5711));
MXI2XL addgen2_A_I1211 (.Y(N658), .A(N5721), .B(N5720), .S0(N2867));
MXI2XL addgen2_A_I1212 (.Y(N2876), .A(N5631), .B(N5630), .S0(N5711));
MXI2XL addgen2_A_I1213 (.Y(N659), .A(N5721), .B(N5720), .S0(N2876));
MXI2XL addgen2_A_I1214 (.Y(N2885), .A(N5632), .B(N5631), .S0(N5711));
MXI2XL addgen2_A_I1215 (.Y(N660), .A(N5721), .B(N5720), .S0(N2885));
MXI2XL addgen2_A_I1216 (.Y(N2894), .A(N5633), .B(N5632), .S0(N5711));
MXI2XL addgen2_A_I1217 (.Y(N661), .A(N5721), .B(N5720), .S0(N2894));
MXI2XL addgen2_A_I1218 (.Y(N2903), .A(N5634), .B(N5633), .S0(N5711));
MXI2XL addgen2_A_I1219 (.Y(N662), .A(N5721), .B(N5720), .S0(N2903));
MXI2XL addgen2_A_I1220 (.Y(N2912), .A(N5635), .B(N5634), .S0(N5711));
MXI2XL addgen2_A_I1221 (.Y(N663), .A(N5721), .B(N5720), .S0(N2912));
MXI2XL addgen2_A_I1222 (.Y(N2921), .A(N5636), .B(N5635), .S0(N5711));
MXI2XL addgen2_A_I1223 (.Y(N664), .A(N5721), .B(N5720), .S0(N2921));
MXI2XL addgen2_A_I1224 (.Y(N2930), .A(N5637), .B(N5636), .S0(N5711));
MXI2XL addgen2_A_I1225 (.Y(N665), .A(N5721), .B(N5720), .S0(N2930));
MXI2XL addgen2_A_I1226 (.Y(N2939), .A(N5638), .B(N5637), .S0(N5711));
MXI2XL addgen2_A_I1227 (.Y(N666), .A(N5721), .B(N5720), .S0(N2939));
MXI2XL addgen2_A_I1228 (.Y(N2948), .A(N5639), .B(N5638), .S0(N5712));
MXI2XL addgen2_A_I1229 (.Y(N667), .A(N5721), .B(N5720), .S0(N2948));
MXI2XL addgen2_A_I1230 (.Y(N2957), .A(N5640), .B(N5639), .S0(N5712));
MXI2XL addgen2_A_I1231 (.Y(N668), .A(N5721), .B(N5720), .S0(N2957));
MXI2XL addgen2_A_I1232 (.Y(N2966), .A(N5641), .B(N5640), .S0(N5712));
MXI2XL addgen2_A_I1233 (.Y(N669), .A(N5721), .B(N5720), .S0(N2966));
MXI2XL addgen2_A_I1234 (.Y(N2975), .A(N5642), .B(N5641), .S0(N5712));
MXI2XL addgen2_A_I1235 (.Y(N670), .A(N5721), .B(N5720), .S0(N2975));
MXI2XL addgen2_A_I1236 (.Y(N2984), .A(N5643), .B(N5642), .S0(N5712));
MXI2XL addgen2_A_I1237 (.Y(N671), .A(N5721), .B(N5720), .S0(N2984));
MXI2XL addgen2_A_I1238 (.Y(N2993), .A(N5644), .B(N5643), .S0(N5712));
MXI2XL addgen2_A_I1239 (.Y(N672), .A(N5721), .B(N5720), .S0(N2993));
MXI2XL addgen2_A_I1240 (.Y(N3002), .A(N5645), .B(N5644), .S0(N5712));
MXI2XL addgen2_A_I1241 (.Y(N673), .A(N5721), .B(N5720), .S0(N3002));
MXI2XL addgen2_A_I1242 (.Y(N3011), .A(N5646), .B(N5645), .S0(N5712));
MXI2XL addgen2_A_I1243 (.Y(N674), .A(N5721), .B(N5720), .S0(N3011));
NAND2XL addgen2_A_I1244 (.Y(N3020), .A(N5646), .B(N5712));
MXI2XL addgen2_A_I1245 (.Y(N675), .A(N5721), .B(N5720), .S0(N3020));
NAND2XL enc2_A_I1247 (.Y(N3029), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
NOR2XL enc2_A_I1248 (.Y(N3031), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
AND2XL enc2_A_I1249 (.Y(N681), .A(N3029), .B(inst_cellmath__203_0_in1[27]));
XOR2XL inst_cellmath__203_0_I2206 (.Y(N5722), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
INVXL inst_cellmath__203_0_I1923 (.Y(N5728), .A(N5722));
INVXL inst_cellmath__203_0_I1922 (.Y(N5727), .A(N5722));
OR2XL inst_cellmath__203_0_I4814 (.Y(N5736), .A(N3031), .B(inst_cellmath__203_0_in1[27]));
INVXL inst_cellmath__203_0_I1932 (.Y(N5737), .A(N681));
NOR2XL addgen2_A_I1251 (.Y(N3042), .A(N5627), .B(N5728));
MXI2XL addgen2_A_I1252 (.Y(N685), .A(N5737), .B(N5736), .S0(N3042));
MXI2XL addgen2_A_I1253 (.Y(N3051), .A(N5628), .B(N5627), .S0(N5728));
MXI2XL addgen2_A_I1254 (.Y(N686), .A(N5737), .B(N5736), .S0(N3051));
MXI2XL addgen2_A_I1255 (.Y(N3060), .A(N5629), .B(N5628), .S0(N5727));
MXI2XL addgen2_A_I1256 (.Y(N687), .A(N5737), .B(N5736), .S0(N3060));
MXI2XL addgen2_A_I1257 (.Y(N3069), .A(N5630), .B(N5629), .S0(N5727));
MXI2XL addgen2_A_I1258 (.Y(N688), .A(N5737), .B(N5736), .S0(N3069));
MXI2XL addgen2_A_I1259 (.Y(N3078), .A(N5631), .B(N5630), .S0(N5727));
MXI2XL addgen2_A_I1260 (.Y(N689), .A(N5737), .B(N5736), .S0(N3078));
MXI2XL addgen2_A_I1261 (.Y(N3087), .A(N5632), .B(N5631), .S0(N5727));
MXI2XL addgen2_A_I1262 (.Y(N690), .A(N5737), .B(N5736), .S0(N3087));
MXI2XL addgen2_A_I1263 (.Y(N3096), .A(N5633), .B(N5632), .S0(N5727));
MXI2XL addgen2_A_I1264 (.Y(N691), .A(N5737), .B(N5736), .S0(N3096));
MXI2XL addgen2_A_I1265 (.Y(N3105), .A(N5634), .B(N5633), .S0(N5727));
MXI2XL addgen2_A_I1266 (.Y(N692), .A(N5737), .B(N5736), .S0(N3105));
MXI2XL addgen2_A_I1267 (.Y(N3114), .A(N5635), .B(N5634), .S0(N5727));
MXI2XL addgen2_A_I1268 (.Y(N693), .A(N5737), .B(N5736), .S0(N3114));
MXI2XL addgen2_A_I1269 (.Y(N3123), .A(N5636), .B(N5635), .S0(N5727));
MXI2XL addgen2_A_I1270 (.Y(N694), .A(N5737), .B(N5736), .S0(N3123));
MXI2XL addgen2_A_I1271 (.Y(N3132), .A(N5637), .B(N5636), .S0(N5728));
MXI2XL addgen2_A_I1272 (.Y(N695), .A(N5737), .B(N5736), .S0(N3132));
MXI2XL addgen2_A_I1273 (.Y(N3141), .A(N5638), .B(N5637), .S0(N5728));
MXI2XL addgen2_A_I1274 (.Y(N696), .A(N5737), .B(N5736), .S0(N3141));
MXI2XL addgen2_A_I1275 (.Y(N3150), .A(N5639), .B(N5638), .S0(N5728));
MXI2XL addgen2_A_I1276 (.Y(N697), .A(N5737), .B(N5736), .S0(N3150));
MXI2XL addgen2_A_I1277 (.Y(N3159), .A(N5640), .B(N5639), .S0(N5728));
MXI2XL addgen2_A_I1278 (.Y(N698), .A(N5737), .B(N5736), .S0(N3159));
MXI2XL addgen2_A_I1279 (.Y(N3168), .A(N5641), .B(N5640), .S0(N5728));
MXI2XL addgen2_A_I1280 (.Y(N699), .A(N5737), .B(N5736), .S0(N3168));
MXI2XL addgen2_A_I1281 (.Y(N3177), .A(N5642), .B(N5641), .S0(N5728));
MXI2XL addgen2_A_I1282 (.Y(N700), .A(N5737), .B(N5736), .S0(N3177));
MXI2XL addgen2_A_I1283 (.Y(N3186), .A(N5643), .B(N5642), .S0(N5728));
MXI2XL addgen2_A_I1284 (.Y(N701), .A(N5737), .B(N5736), .S0(N3186));
MXI2XL addgen2_A_I1285 (.Y(N3195), .A(N5644), .B(N5643), .S0(N5728));
MXI2XL addgen2_A_I1286 (.Y(N702), .A(N5737), .B(N5736), .S0(N3195));
MXI2XL addgen2_A_I1287 (.Y(N3204), .A(N5645), .B(N5644), .S0(N5728));
MXI2XL addgen2_A_I1288 (.Y(N703), .A(N5737), .B(N5736), .S0(N3204));
MXI2XL addgen2_A_I1289 (.Y(N3213), .A(N5646), .B(N5645), .S0(N5728));
MXI2XL addgen2_A_I1290 (.Y(N704), .A(N5737), .B(N5736), .S0(N3213));
NAND2XL addgen2_A_I1291 (.Y(N3222), .A(N5646), .B(N5728));
MXI2XL addgen2_A_I1292 (.Y(N705), .A(N5737), .B(N5736), .S0(N3222));
NAND2XL enc2_A_I1294 (.Y(N3231), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
NOR2XL enc2_A_I1295 (.Y(N3233), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
AND2XL enc2_A_I1296 (.Y(N711), .A(N3231), .B(inst_cellmath__203_0_in1[29]));
XOR2XL inst_cellmath__203_0_I4815 (.Y(N5738), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
INVX1 inst_cellmath__203_0_I1937 (.Y(N5742), .A(N5738));
OR2XL inst_cellmath__203_0_I2208 (.Y(N5751), .A(N3233), .B(inst_cellmath__203_0_in1[29]));
INVXL inst_cellmath__203_0_I1947 (.Y(N5752), .A(N711));
NOR2XL addgen2_A_I1298 (.Y(N3244), .A(N5627), .B(N5742));
MXI2XL addgen2_A_I1299 (.Y(N715), .A(N5752), .B(N5751), .S0(N3244));
MXI2XL addgen2_A_I2209 (.Y(N3253), .A(N5627), .B(N5628), .S0(N5738));
MXI2XL addgen2_A_I1301 (.Y(N716), .A(N5752), .B(N5751), .S0(N3253));
MXI2XL addgen2_A_I1302 (.Y(N3262), .A(N5629), .B(N5628), .S0(N5742));
MXI2XL addgen2_A_I1303 (.Y(N717), .A(N5752), .B(N5751), .S0(N3262));
MXI2XL addgen2_A_I1304 (.Y(N3271), .A(N5630), .B(N5629), .S0(N5742));
MXI2XL addgen2_A_I1305 (.Y(N718), .A(N5752), .B(N5751), .S0(N3271));
MXI2XL addgen2_A_I1306 (.Y(N3280), .A(N5631), .B(N5630), .S0(N5742));
MXI2XL addgen2_A_I1307 (.Y(N719), .A(N5752), .B(N5751), .S0(N3280));
MXI2XL addgen2_A_I1308 (.Y(N3289), .A(N5632), .B(N5631), .S0(N5742));
MXI2XL addgen2_A_I1309 (.Y(N720), .A(N5752), .B(N5751), .S0(N3289));
MXI2XL addgen2_A_I1310 (.Y(N3298), .A(N5633), .B(N5632), .S0(N5742));
MXI2XL addgen2_A_I1311 (.Y(N721), .A(N5752), .B(N5751), .S0(N3298));
MXI2XL addgen2_A_I1312 (.Y(N3307), .A(N5634), .B(N5633), .S0(N5742));
MXI2XL addgen2_A_I1313 (.Y(N722), .A(N5752), .B(N5751), .S0(N3307));
MXI2XL addgen2_A_I1314 (.Y(N3316), .A(N5635), .B(N5634), .S0(N5742));
MXI2XL addgen2_A_I1315 (.Y(N723), .A(N5752), .B(N5751), .S0(N3316));
MXI2XL addgen2_A_I1316 (.Y(N3325), .A(N5636), .B(N5635), .S0(N5742));
MXI2XL addgen2_A_I1317 (.Y(N724), .A(N5752), .B(N5751), .S0(N3325));
MXI2XL addgen2_A_I1318 (.Y(N3334), .A(N5637), .B(N5636), .S0(N5742));
MXI2XL addgen2_A_I1319 (.Y(N725), .A(N5752), .B(N5751), .S0(N3334));
MXI2XL addgen2_A_I1320 (.Y(N3343), .A(N5638), .B(N5637), .S0(N5742));
MXI2XL addgen2_A_I1321 (.Y(N726), .A(N5752), .B(N5751), .S0(N3343));
MXI2XL addgen2_A_I1322 (.Y(N3352), .A(N5639), .B(N5638), .S0(N5742));
MXI2XL addgen2_A_I1323 (.Y(N727), .A(N5752), .B(N5751), .S0(N3352));
MXI2XL addgen2_A_I1324 (.Y(N3361), .A(N5640), .B(N5639), .S0(N5742));
MXI2XL addgen2_A_I1325 (.Y(N728), .A(N5752), .B(N5751), .S0(N3361));
MXI2XL addgen2_A_I1326 (.Y(N3370), .A(N5641), .B(N5640), .S0(N5742));
MXI2XL addgen2_A_I1327 (.Y(N729), .A(N5752), .B(N5751), .S0(N3370));
MXI2XL addgen2_A_I1328 (.Y(N3379), .A(N5642), .B(N5641), .S0(N5742));
MXI2XL addgen2_A_I1329 (.Y(N730), .A(N5752), .B(N5751), .S0(N3379));
MXI2XL addgen2_A_I1330 (.Y(N3388), .A(N5643), .B(N5642), .S0(N5742));
MXI2XL addgen2_A_I1331 (.Y(N731), .A(N5752), .B(N5751), .S0(N3388));
MXI2XL addgen2_A_I1332 (.Y(N3397), .A(N5644), .B(N5643), .S0(N5742));
MXI2XL addgen2_A_I1333 (.Y(N732), .A(N5752), .B(N5751), .S0(N3397));
MXI2XL addgen2_A_I1334 (.Y(N3406), .A(N5645), .B(N5644), .S0(N5742));
MXI2XL addgen2_A_I1335 (.Y(N733), .A(N5752), .B(N5751), .S0(N3406));
MXI2XL addgen2_A_I1336 (.Y(N3415), .A(N5646), .B(N5645), .S0(N5742));
MXI2XL addgen2_A_I1337 (.Y(N734), .A(N5752), .B(N5751), .S0(N3415));
NAND2XL addgen2_A_I1338 (.Y(N3424), .A(N5646), .B(N5742));
MXI2XL addgen2_A_I1339 (.Y(N735), .A(N5752), .B(N5751), .S0(N3424));
NAND2XL enc2_A_I1341 (.Y(N3433), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
NOR2XL enc2_A_I1342 (.Y(N3435), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
AND2XL enc2_A_I1343 (.Y(N741), .A(N3433), .B(inst_cellmath__203_0_in1[31]));
XOR2XL inst_cellmath__203_0_I2210 (.Y(N5753), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
INVXL inst_cellmath__203_0_I1954 (.Y(N5759), .A(N5753));
INVXL inst_cellmath__203_0_I1953 (.Y(N5758), .A(N5753));
OR2XL inst_cellmath__203_0_I2211 (.Y(N5767), .A(N3435), .B(inst_cellmath__203_0_in1[31]));
INVXL inst_cellmath__203_0_I1963 (.Y(N5768), .A(N741));
NOR2XL addgen2_A_I1345 (.Y(N3446), .A(N5627), .B(N5758));
MXI2XL addgen2_A_I1346 (.Y(N745), .A(N5768), .B(N5767), .S0(N3446));
MXI2XL addgen2_A_I1347 (.Y(N3455), .A(N5628), .B(N5627), .S0(N5759));
MXI2XL addgen2_A_I1348 (.Y(N746), .A(N5768), .B(N5767), .S0(N3455));
MXI2XL addgen2_A_I1349 (.Y(N3464), .A(N5629), .B(N5628), .S0(N5758));
MXI2XL addgen2_A_I1350 (.Y(N747), .A(N5768), .B(N5767), .S0(N3464));
MXI2XL addgen2_A_I1351 (.Y(N3473), .A(N5630), .B(N5629), .S0(N5758));
MXI2XL addgen2_A_I1352 (.Y(N748), .A(N5768), .B(N5767), .S0(N3473));
MXI2XL addgen2_A_I1353 (.Y(N3482), .A(N5631), .B(N5630), .S0(N5758));
MXI2XL addgen2_A_I1354 (.Y(N749), .A(N5768), .B(N5767), .S0(N3482));
MXI2XL addgen2_A_I1355 (.Y(N3491), .A(N5632), .B(N5631), .S0(N5758));
MXI2XL addgen2_A_I1356 (.Y(N750), .A(N5768), .B(N5767), .S0(N3491));
MXI2XL addgen2_A_I1357 (.Y(N3500), .A(N5633), .B(N5632), .S0(N5758));
MXI2XL addgen2_A_I1358 (.Y(N751), .A(N5768), .B(N5767), .S0(N3500));
MXI2XL addgen2_A_I1359 (.Y(N3509), .A(N5634), .B(N5633), .S0(N5758));
MXI2XL addgen2_A_I1360 (.Y(N752), .A(N5768), .B(N5767), .S0(N3509));
MXI2XL addgen2_A_I1361 (.Y(N3518), .A(N5635), .B(N5634), .S0(N5758));
MXI2XL addgen2_A_I1362 (.Y(N753), .A(N5768), .B(N5767), .S0(N3518));
MXI2XL addgen2_A_I1363 (.Y(N3527), .A(N5636), .B(N5635), .S0(N5758));
MXI2XL addgen2_A_I1364 (.Y(N754), .A(N5768), .B(N5767), .S0(N3527));
MXI2XL addgen2_A_I1365 (.Y(N3536), .A(N5637), .B(N5636), .S0(N5758));
MXI2XL addgen2_A_I1366 (.Y(N755), .A(N5768), .B(N5767), .S0(N3536));
MXI2XL addgen2_A_I1367 (.Y(N3545), .A(N5638), .B(N5637), .S0(N5758));
MXI2XL addgen2_A_I1368 (.Y(N756), .A(N5768), .B(N5767), .S0(N3545));
MXI2XL addgen2_A_I1369 (.Y(N3554), .A(N5639), .B(N5638), .S0(N5758));
MXI2XL addgen2_A_I1370 (.Y(N757), .A(N5768), .B(N5767), .S0(N3554));
MXI2XL addgen2_A_I1371 (.Y(N3563), .A(N5640), .B(N5639), .S0(N5758));
MXI2XL addgen2_A_I1372 (.Y(N758), .A(N5768), .B(N5767), .S0(N3563));
MXI2XL addgen2_A_I1373 (.Y(N3572), .A(N5641), .B(N5640), .S0(N5759));
MXI2XL addgen2_A_I1374 (.Y(N759), .A(N5768), .B(N5767), .S0(N3572));
MXI2XL addgen2_A_I1375 (.Y(N3581), .A(N5642), .B(N5641), .S0(N5759));
MXI2XL addgen2_A_I1376 (.Y(N760), .A(N5768), .B(N5767), .S0(N3581));
MXI2XL addgen2_A_I1377 (.Y(N3590), .A(N5643), .B(N5642), .S0(N5759));
MXI2XL addgen2_A_I1378 (.Y(N761), .A(N5768), .B(N5767), .S0(N3590));
MXI2XL addgen2_A_I1379 (.Y(N3599), .A(N5644), .B(N5643), .S0(N5759));
MXI2XL addgen2_A_I1380 (.Y(N762), .A(N5768), .B(N5767), .S0(N3599));
MXI2XL addgen2_A_I1381 (.Y(N3608), .A(N5645), .B(N5644), .S0(N5758));
MXI2XL addgen2_A_I1382 (.Y(N763), .A(N5768), .B(N5767), .S0(N3608));
MXI2XL addgen2_A_I1383 (.Y(N3617), .A(N5646), .B(N5645), .S0(N5758));
MXI2XL addgen2_A_I1384 (.Y(N764), .A(N5768), .B(N5767), .S0(N3617));
NAND2XL addgen2_A_I1385 (.Y(N3626), .A(N5646), .B(N5758));
MXI2XL addgen2_A_I1386 (.Y(N765), .A(N5768), .B(N5767), .S0(N3626));
ADDHX1 inst_cellmath__203_0_I281 (.CO(N770), .S(N768), .A(inst_cellmath__203_0_in1[32]), .B(inst_cellmath__203_0_in1[31]));
INVXL inst_cellmath__203_0_I1964 (.Y(N5769), .A(N768));
INVXL inst_cellmath__203_0_I1965 (.Y(N5770), .A(N770));
NOR2XL inst_cellmath__203_0_I285 (.Y(N779), .A(N5769), .B(N5627));
OAI22XL inst_cellmath__203_0_I286 (.Y(N781), .A0(N5627), .A1(N5770), .B0(N5769), .B1(N5628));
OAI22XL inst_cellmath__203_0_I287 (.Y(N783), .A0(N5628), .A1(N5770), .B0(N5769), .B1(N5629));
OAI22XL inst_cellmath__203_0_I288 (.Y(N785), .A0(N5629), .A1(N5770), .B0(N5769), .B1(N5630));
OAI22XL inst_cellmath__203_0_I289 (.Y(N787), .A0(N5630), .A1(N5770), .B0(N5769), .B1(N5631));
OAI22XL inst_cellmath__203_0_I290 (.Y(N789), .A0(N5631), .A1(N5770), .B0(N5769), .B1(N5632));
OAI22XL inst_cellmath__203_0_I291 (.Y(N791), .A0(N5632), .A1(N5770), .B0(N5769), .B1(N5633));
OAI22XL inst_cellmath__203_0_I292 (.Y(N793), .A0(N5633), .A1(N5770), .B0(N5769), .B1(N5634));
OAI22XL inst_cellmath__203_0_I293 (.Y(N795), .A0(N5634), .A1(N5770), .B0(N5769), .B1(N5635));
OAI22XL inst_cellmath__203_0_I294 (.Y(N797), .A0(N5635), .A1(N5770), .B0(N5769), .B1(N5636));
OAI22XL inst_cellmath__203_0_I295 (.Y(N799), .A0(N5636), .A1(N5770), .B0(N5769), .B1(N5637));
OAI22XL inst_cellmath__203_0_I296 (.Y(N801), .A0(N5637), .A1(N5770), .B0(N5769), .B1(N5638));
OAI22XL inst_cellmath__203_0_I297 (.Y(N803), .A0(N5638), .A1(N5770), .B0(N5769), .B1(N5639));
OAI22XL inst_cellmath__203_0_I298 (.Y(N805), .A0(N5639), .A1(N5770), .B0(N5769), .B1(N5640));
OAI22XL inst_cellmath__203_0_I299 (.Y(N807), .A0(N5640), .A1(N5770), .B0(N5769), .B1(N5641));
OAI22XL inst_cellmath__203_0_I300 (.Y(N809), .A0(N5641), .A1(N5770), .B0(N5769), .B1(N5642));
OAI22XL inst_cellmath__203_0_I301 (.Y(N811), .A0(N5642), .A1(N5770), .B0(N5769), .B1(N5643));
OAI22XL inst_cellmath__203_0_I302 (.Y(N813), .A0(N5643), .A1(N5770), .B0(N5769), .B1(N5644));
OAI22XL inst_cellmath__203_0_I303 (.Y(N815), .A0(N5644), .A1(N5770), .B0(N5769), .B1(N5645));
OAI22XL inst_cellmath__203_0_I304 (.Y(N817), .A0(N5645), .A1(N5770), .B0(N5769), .B1(N5646));
OAI21XL inst_cellmath__203_0_I305 (.Y(N819), .A0(N5770), .A1(N5646), .B0(N5769));
AND2XL inst_cellmath__203_0_I306 (.Y(N1366), .A(N5770), .B(N5769));
INVXL inst_cellmath__203_0_I1966 (.Y(N5771), .A(inst_cellmath__203_0_in3[0]));
INVXL inst_cellmath__203_0_I1967 (.Y(N5772), .A(inst_cellmath__203_0_in3[1]));
INVXL inst_cellmath__203_0_I1968 (.Y(N5773), .A(inst_cellmath__203_0_in3[2]));
INVXL inst_cellmath__203_0_I1969 (.Y(N5774), .A(inst_cellmath__203_0_in3[3]));
INVXL inst_cellmath__203_0_I1970 (.Y(N5775), .A(inst_cellmath__203_0_in3[4]));
INVXL inst_cellmath__203_0_I1971 (.Y(N5776), .A(inst_cellmath__203_0_in3[5]));
INVXL inst_cellmath__203_0_I1972 (.Y(N5777), .A(inst_cellmath__203_0_in3[6]));
INVXL inst_cellmath__203_0_I1973 (.Y(N5778), .A(inst_cellmath__203_0_in3[7]));
INVXL inst_cellmath__203_0_I1974 (.Y(N5779), .A(inst_cellmath__203_0_in3[8]));
INVXL inst_cellmath__203_0_I1975 (.Y(N5780), .A(inst_cellmath__203_0_in3[9]));
INVXL inst_cellmath__203_0_I1976 (.Y(N5781), .A(inst_cellmath__203_0_in3[10]));
INVXL inst_cellmath__203_0_I1977 (.Y(N5782), .A(inst_cellmath__203_0_in3[11]));
INVXL inst_cellmath__203_0_I1978 (.Y(N5783), .A(inst_cellmath__203_0_in3[12]));
INVXL inst_cellmath__203_0_I1979 (.Y(N5784), .A(inst_cellmath__203_0_in3[13]));
INVXL inst_cellmath__203_0_I1980 (.Y(N5785), .A(inst_cellmath__203_0_in3[14]));
INVXL inst_cellmath__203_0_I1981 (.Y(N5786), .A(inst_cellmath__203_0_in3[15]));
INVXL inst_cellmath__203_0_I1982 (.Y(N5787), .A(inst_cellmath__203_0_in3[16]));
INVXL inst_cellmath__203_0_I1983 (.Y(N5788), .A(inst_cellmath__203_0_in3[17]));
INVXL inst_cellmath__203_0_I1984 (.Y(N5789), .A(inst_cellmath__203_0_in3[18]));
INVXL inst_cellmath__203_0_I1985 (.Y(N5790), .A(inst_cellmath__203_0_in3[19]));
INVXL inst_cellmath__203_0_I1986 (.Y(N5791), .A(inst_cellmath__203_0_in3[20]));
INVXL inst_cellmath__203_0_I1987 (.Y(N5792), .A(inst_cellmath__203_0_in3[21]));
INVXL inst_cellmath__203_0_I1988 (.Y(N5793), .A(inst_cellmath__203_0_in0[0]));
NOR2XL inst_cellmath__203_0_I382 (.Y(N1025), .A(N5793), .B(N5771));
NOR2XL inst_cellmath__203_0_I383 (.Y(N1027), .A(N5793), .B(N5772));
NOR2XL inst_cellmath__203_0_I384 (.Y(N1029), .A(N5793), .B(N5773));
NOR2XL inst_cellmath__203_0_I385 (.Y(N1031), .A(N5793), .B(N5774));
NOR2XL inst_cellmath__203_0_I386 (.Y(N1033), .A(N5793), .B(N5775));
NOR2XL inst_cellmath__203_0_I387 (.Y(N1035), .A(N5793), .B(N5776));
NOR2XL inst_cellmath__203_0_I388 (.Y(N1037), .A(N5793), .B(N5777));
NOR2XL inst_cellmath__203_0_I389 (.Y(N1039), .A(N5793), .B(N5778));
NOR2XL inst_cellmath__203_0_I390 (.Y(N1041), .A(N5793), .B(N5779));
NOR2XL inst_cellmath__203_0_I391 (.Y(N1043), .A(N5793), .B(N5780));
NOR2XL inst_cellmath__203_0_I392 (.Y(N1045), .A(N5793), .B(N5781));
NOR2XL inst_cellmath__203_0_I393 (.Y(N1047), .A(N5793), .B(N5782));
NOR2XL inst_cellmath__203_0_I394 (.Y(N1049), .A(N5793), .B(N5783));
NOR2XL inst_cellmath__203_0_I395 (.Y(N1051), .A(N5793), .B(N5784));
NOR2XL inst_cellmath__203_0_I396 (.Y(N1053), .A(N5793), .B(N5785));
NOR2XL inst_cellmath__203_0_I397 (.Y(N1055), .A(N5793), .B(N5786));
NOR2XL inst_cellmath__203_0_I398 (.Y(N1732), .A(N5793), .B(N5787));
NOR2XL inst_cellmath__203_0_I399 (.Y(N1059), .A(N5793), .B(N5788));
NOR2XL inst_cellmath__203_0_I400 (.Y(N1061), .A(N5793), .B(N5789));
NOR2XL inst_cellmath__203_0_I401 (.Y(N1798), .A(N5793), .B(N5790));
NOR2XL inst_cellmath__203_0_I402 (.Y(N1830), .A(N5793), .B(N5791));
NOR2XL inst_cellmath__203_0_I403 (.Y(N1067), .A(N5793), .B(N5792));
INVXL inst_cellmath__203_0_I1989 (.Y(N5794), .A(inst_cellmath__203_0_in0[1]));
OR2XL inst_cellmath__203_0_I2213 (.Y(N5804), .A(N5794), .B(inst_cellmath__203_0_in0[2]));
INVXL inst_cellmath__203_0_I2015 (.Y(N5820), .A(inst_cellmath__203_0_in0[2]));
NOR2XL addgen2_A_I1392 (.Y(N3648), .A(N5771), .B(N5794));
MXI2XL addgen2_A_I1393 (.Y(N1077), .A(N5820), .B(N5804), .S0(N3648));
MXI2XL addgen2_A_I1394 (.Y(N3657), .A(N5772), .B(N5771), .S0(N5794));
MXI2XL addgen2_A_I1395 (.Y(N1078), .A(N5820), .B(N5804), .S0(N3657));
MXI2XL addgen2_A_I1396 (.Y(N3666), .A(N5773), .B(N5772), .S0(N5794));
MXI2XL addgen2_A_I1397 (.Y(N1079), .A(N5820), .B(N5804), .S0(N3666));
MXI2XL addgen2_A_I1398 (.Y(N3675), .A(N5774), .B(N5773), .S0(N5794));
MXI2XL addgen2_A_I1399 (.Y(N1080), .A(N5820), .B(N5804), .S0(N3675));
MXI2XL addgen2_A_I1400 (.Y(N3684), .A(N5775), .B(N5774), .S0(N5794));
MXI2XL addgen2_A_I1401 (.Y(N1081), .A(N5820), .B(N5804), .S0(N3684));
MXI2XL addgen2_A_I1402 (.Y(N3693), .A(N5776), .B(N5775), .S0(N5794));
MXI2XL addgen2_A_I1403 (.Y(N1082), .A(N5820), .B(N5804), .S0(N3693));
MXI2XL addgen2_A_I1404 (.Y(N3702), .A(N5777), .B(N5776), .S0(N5794));
MXI2XL addgen2_A_I1405 (.Y(N1083), .A(N5820), .B(N5804), .S0(N3702));
MXI2XL addgen2_A_I1406 (.Y(N3711), .A(N5778), .B(N5777), .S0(N5794));
MXI2XL addgen2_A_I1407 (.Y(N1084), .A(N5820), .B(N5804), .S0(N3711));
MXI2XL addgen2_A_I1408 (.Y(N3720), .A(N5779), .B(N5778), .S0(N5794));
MXI2XL addgen2_A_I1409 (.Y(N1085), .A(N5820), .B(N5804), .S0(N3720));
MXI2XL addgen2_A_I1410 (.Y(N3729), .A(N5780), .B(N5779), .S0(N5794));
MXI2XL addgen2_A_I1411 (.Y(N1086), .A(N5820), .B(N5804), .S0(N3729));
MXI2XL addgen2_A_I1412 (.Y(N3738), .A(N5781), .B(N5780), .S0(N5794));
MXI2XL addgen2_A_I1413 (.Y(N1087), .A(N5820), .B(N5804), .S0(N3738));
MXI2XL addgen2_A_I1414 (.Y(N3747), .A(N5782), .B(N5781), .S0(N5794));
MXI2XL addgen2_A_I1415 (.Y(N1088), .A(N5820), .B(N5804), .S0(N3747));
MXI2XL addgen2_A_I1416 (.Y(N3756), .A(N5783), .B(N5782), .S0(N5794));
MXI2XL addgen2_A_I1417 (.Y(N1089), .A(N5820), .B(N5804), .S0(N3756));
MXI2XL addgen2_A_I1418 (.Y(N3765), .A(N5784), .B(N5783), .S0(N5794));
MXI2XL addgen2_A_I1419 (.Y(N1090), .A(N5820), .B(N5804), .S0(N3765));
MXI2XL addgen2_A_I1420 (.Y(N3774), .A(N5785), .B(N5784), .S0(N5794));
MXI2XL addgen2_A_I1421 (.Y(N1091), .A(N5820), .B(N5804), .S0(N3774));
MXI2XL addgen2_A_I1422 (.Y(N3783), .A(N5786), .B(N5785), .S0(N5794));
MXI2XL addgen2_A_I1423 (.Y(N1092), .A(N5820), .B(N5804), .S0(N3783));
MXI2XL addgen2_A_I1424 (.Y(N3792), .A(N5787), .B(N5786), .S0(N5794));
MXI2XL addgen2_A_I1425 (.Y(N1093), .A(N5820), .B(N5804), .S0(N3792));
MXI2XL addgen2_A_I1426 (.Y(N3801), .A(N5788), .B(N5787), .S0(N5794));
MXI2XL addgen2_A_I1427 (.Y(N1094), .A(N5820), .B(N5804), .S0(N3801));
MXI2XL addgen2_A_I1428 (.Y(N3810), .A(N5789), .B(N5788), .S0(N5794));
MXI2XL addgen2_A_I1429 (.Y(N1095), .A(N5820), .B(N5804), .S0(N3810));
MXI2XL addgen2_A_I1430 (.Y(N3819), .A(N5790), .B(N5789), .S0(N5794));
MXI2XL addgen2_A_I1431 (.Y(N1096), .A(N5820), .B(N5804), .S0(N3819));
MXI2XL addgen2_A_I1432 (.Y(N3828), .A(N5791), .B(N5790), .S0(N5794));
MXI2XL addgen2_A_I1433 (.Y(N1097), .A(N5820), .B(N5804), .S0(N3828));
MXI2XL addgen2_A_I1434 (.Y(N3837), .A(N5792), .B(N5791), .S0(N5794));
MXI2XL addgen2_A_I1435 (.Y(N1098), .A(N5820), .B(N5804), .S0(N3837));
NOR2BX1 addgen2_A_I1436 (.Y(N3846), .AN(N5794), .B(N5792));
MXI2XL addgen2_A_I1437 (.Y(N1099), .A(N5820), .B(N5804), .S0(N3846));
XNOR2X1 enc2_A_I1438 (.Y(N1103), .A(inst_cellmath__203_0_in0[3]), .B(inst_cellmath__203_0_in0[2]));
NAND2XL enc2_A_I1439 (.Y(N3855), .A(inst_cellmath__203_0_in0[3]), .B(inst_cellmath__203_0_in0[2]));
NOR2XL enc2_A_I1440 (.Y(N3857), .A(inst_cellmath__203_0_in0[3]), .B(inst_cellmath__203_0_in0[2]));
AND2XL enc2_A_I1441 (.Y(N1105), .A(N3855), .B(inst_cellmath__203_0_in0[4]));
OR2XL inst_cellmath__203_0_I2216 (.Y(N5839), .A(N3857), .B(inst_cellmath__203_0_in0[4]));
INVXL inst_cellmath__203_0_I2043 (.Y(N5848), .A(N1105));
NOR2XL addgen2_A_I1443 (.Y(N3868), .A(N5771), .B(N1103));
MXI2XL addgen2_A_I1444 (.Y(N1109), .A(N5848), .B(N5839), .S0(N3868));
MXI2XL addgen2_A_I1445 (.Y(N3877), .A(N5772), .B(N5771), .S0(N1103));
MXI2XL addgen2_A_I1446 (.Y(N1110), .A(N5848), .B(N5839), .S0(N3877));
MXI2XL addgen2_A_I1447 (.Y(N3886), .A(N5773), .B(N5772), .S0(N1103));
MXI2XL addgen2_A_I1448 (.Y(N1111), .A(N5848), .B(N5839), .S0(N3886));
MXI2XL addgen2_A_I1449 (.Y(N3895), .A(N5774), .B(N5773), .S0(N1103));
MXI2XL addgen2_A_I1450 (.Y(N1112), .A(N5848), .B(N5839), .S0(N3895));
MXI2XL addgen2_A_I1451 (.Y(N3904), .A(N5775), .B(N5774), .S0(N1103));
MXI2XL addgen2_A_I1452 (.Y(N1113), .A(N5848), .B(N5839), .S0(N3904));
MXI2XL addgen2_A_I1453 (.Y(N3913), .A(N5776), .B(N5775), .S0(N1103));
MXI2XL addgen2_A_I1454 (.Y(N1114), .A(N5848), .B(N5839), .S0(N3913));
MXI2XL addgen2_A_I1455 (.Y(N3922), .A(N5777), .B(N5776), .S0(N1103));
MXI2XL addgen2_A_I1456 (.Y(N1115), .A(N5848), .B(N5839), .S0(N3922));
MXI2XL addgen2_A_I1457 (.Y(N3931), .A(N5778), .B(N5777), .S0(N1103));
MXI2XL addgen2_A_I1458 (.Y(N1116), .A(N5848), .B(N5839), .S0(N3931));
MXI2XL addgen2_A_I1459 (.Y(N3940), .A(N5779), .B(N5778), .S0(N1103));
MXI2XL addgen2_A_I1460 (.Y(N1117), .A(N5848), .B(N5839), .S0(N3940));
MXI2XL addgen2_A_I1461 (.Y(N3949), .A(N5780), .B(N5779), .S0(N1103));
MXI2XL addgen2_A_I1462 (.Y(N1118), .A(N5848), .B(N5839), .S0(N3949));
MXI2XL addgen2_A_I1463 (.Y(N3958), .A(N5781), .B(N5780), .S0(N1103));
MXI2XL addgen2_A_I1464 (.Y(N1119), .A(N5848), .B(N5839), .S0(N3958));
MXI2XL addgen2_A_I1465 (.Y(N3967), .A(N5782), .B(N5781), .S0(N1103));
MXI2XL addgen2_A_I1466 (.Y(N1120), .A(N5848), .B(N5839), .S0(N3967));
MXI2XL addgen2_A_I1467 (.Y(N3976), .A(N5783), .B(N5782), .S0(N1103));
MXI2XL addgen2_A_I1468 (.Y(N1121), .A(N5848), .B(N5839), .S0(N3976));
MXI2XL addgen2_A_I1469 (.Y(N3985), .A(N5784), .B(N5783), .S0(N1103));
MXI2XL addgen2_A_I1470 (.Y(N1122), .A(N5848), .B(N5839), .S0(N3985));
MXI2XL addgen2_A_I1471 (.Y(N3994), .A(N5785), .B(N5784), .S0(N1103));
MXI2XL addgen2_A_I1472 (.Y(N1123), .A(N5848), .B(N5839), .S0(N3994));
MXI2XL addgen2_A_I1473 (.Y(N4003), .A(N5786), .B(N5785), .S0(N1103));
MXI2XL addgen2_A_I1474 (.Y(N1124), .A(N5848), .B(N5839), .S0(N4003));
MXI2XL addgen2_A_I1475 (.Y(N4012), .A(N5787), .B(N5786), .S0(N1103));
MXI2XL addgen2_A_I1476 (.Y(N1125), .A(N5848), .B(N5839), .S0(N4012));
MXI2XL addgen2_A_I1477 (.Y(N4021), .A(N5788), .B(N5787), .S0(N1103));
MXI2XL addgen2_A_I1478 (.Y(N1126), .A(N5848), .B(N5839), .S0(N4021));
MXI2XL addgen2_A_I1479 (.Y(N4030), .A(N5789), .B(N5788), .S0(N1103));
MXI2XL addgen2_A_I1480 (.Y(N1127), .A(N5848), .B(N5839), .S0(N4030));
MXI2XL addgen2_A_I1481 (.Y(N4039), .A(N5790), .B(N5789), .S0(N1103));
MXI2XL addgen2_A_I1482 (.Y(N1128), .A(N5848), .B(N5839), .S0(N4039));
MXI2XL addgen2_A_I1483 (.Y(N4048), .A(N5791), .B(N5790), .S0(N1103));
MXI2XL addgen2_A_I1484 (.Y(N1129), .A(N5848), .B(N5839), .S0(N4048));
MXI2XL addgen2_A_I1485 (.Y(N4057), .A(N5792), .B(N5791), .S0(N1103));
MXI2XL addgen2_A_I1486 (.Y(N1130), .A(N5848), .B(N5839), .S0(N4057));
NOR2BX1 addgen2_A_I1487 (.Y(N4066), .AN(N1103), .B(N5792));
MXI2XL addgen2_A_I1488 (.Y(N1131), .A(N5848), .B(N5839), .S0(N4066));
XNOR2X1 enc2_A_I1489 (.Y(N1135), .A(inst_cellmath__203_0_in0[5]), .B(inst_cellmath__203_0_in0[4]));
NAND2XL enc2_A_I1490 (.Y(N4075), .A(inst_cellmath__203_0_in0[5]), .B(inst_cellmath__203_0_in0[4]));
NOR2XL enc2_A_I1491 (.Y(N4077), .A(inst_cellmath__203_0_in0[5]), .B(inst_cellmath__203_0_in0[4]));
AND2XL enc2_A_I1492 (.Y(N1137), .A(N4075), .B(inst_cellmath__203_0_in0[6]));
OR2XL inst_cellmath__203_0_I2218 (.Y(N5865), .A(N4077), .B(inst_cellmath__203_0_in0[6]));
INVXL inst_cellmath__203_0_I2069 (.Y(N5874), .A(N1137));
NOR2XL addgen2_A_I1494 (.Y(N4088), .A(N5771), .B(N1135));
MXI2XL addgen2_A_I1495 (.Y(N1141), .A(N5874), .B(N5865), .S0(N4088));
MXI2XL addgen2_A_I1496 (.Y(N4097), .A(N5772), .B(N5771), .S0(N1135));
MXI2XL addgen2_A_I1497 (.Y(N1142), .A(N5874), .B(N5865), .S0(N4097));
MXI2XL addgen2_A_I1498 (.Y(N4106), .A(N5773), .B(N5772), .S0(N1135));
MXI2XL addgen2_A_I1499 (.Y(N1143), .A(N5874), .B(N5865), .S0(N4106));
MXI2XL addgen2_A_I1500 (.Y(N4115), .A(N5774), .B(N5773), .S0(N1135));
MXI2XL addgen2_A_I1501 (.Y(N1144), .A(N5874), .B(N5865), .S0(N4115));
MXI2XL addgen2_A_I1502 (.Y(N4124), .A(N5775), .B(N5774), .S0(N1135));
MXI2XL addgen2_A_I1503 (.Y(N1145), .A(N5874), .B(N5865), .S0(N4124));
MXI2XL addgen2_A_I1504 (.Y(N4133), .A(N5776), .B(N5775), .S0(N1135));
MXI2XL addgen2_A_I1505 (.Y(N1146), .A(N5874), .B(N5865), .S0(N4133));
MXI2XL addgen2_A_I1506 (.Y(N4142), .A(N5777), .B(N5776), .S0(N1135));
MXI2XL addgen2_A_I1507 (.Y(N1147), .A(N5874), .B(N5865), .S0(N4142));
MXI2XL addgen2_A_I1508 (.Y(N4151), .A(N5778), .B(N5777), .S0(N1135));
MXI2XL addgen2_A_I1509 (.Y(N1148), .A(N5874), .B(N5865), .S0(N4151));
MXI2XL addgen2_A_I1510 (.Y(N4160), .A(N5779), .B(N5778), .S0(N1135));
MXI2XL addgen2_A_I1511 (.Y(N1149), .A(N5874), .B(N5865), .S0(N4160));
MXI2XL addgen2_A_I1512 (.Y(N4169), .A(N5780), .B(N5779), .S0(N1135));
MXI2XL addgen2_A_I1513 (.Y(N1150), .A(N5874), .B(N5865), .S0(N4169));
MXI2XL addgen2_A_I1514 (.Y(N4178), .A(N5781), .B(N5780), .S0(N1135));
MXI2XL addgen2_A_I1515 (.Y(N1151), .A(N5874), .B(N5865), .S0(N4178));
MXI2XL addgen2_A_I1516 (.Y(N4187), .A(N5782), .B(N5781), .S0(N1135));
MXI2XL addgen2_A_I1517 (.Y(N1152), .A(N5874), .B(N5865), .S0(N4187));
MXI2XL addgen2_A_I1518 (.Y(N4196), .A(N5783), .B(N5782), .S0(N1135));
MXI2XL addgen2_A_I1519 (.Y(N1153), .A(N5874), .B(N5865), .S0(N4196));
MXI2XL addgen2_A_I1520 (.Y(N4205), .A(N5784), .B(N5783), .S0(N1135));
MXI2XL addgen2_A_I1521 (.Y(N1154), .A(N5874), .B(N5865), .S0(N4205));
MXI2XL addgen2_A_I1522 (.Y(N4214), .A(N5785), .B(N5784), .S0(N1135));
MXI2XL addgen2_A_I1523 (.Y(N1155), .A(N5874), .B(N5865), .S0(N4214));
MXI2XL addgen2_A_I1524 (.Y(N4223), .A(N5786), .B(N5785), .S0(N1135));
MXI2XL addgen2_A_I1525 (.Y(N1156), .A(N5874), .B(N5865), .S0(N4223));
MXI2XL addgen2_A_I1526 (.Y(N4232), .A(N5787), .B(N5786), .S0(N1135));
MXI2XL addgen2_A_I1527 (.Y(N1157), .A(N5874), .B(N5865), .S0(N4232));
MXI2XL addgen2_A_I1528 (.Y(N4241), .A(N5788), .B(N5787), .S0(N1135));
MXI2XL addgen2_A_I1529 (.Y(N1158), .A(N5874), .B(N5865), .S0(N4241));
MXI2XL addgen2_A_I1530 (.Y(N4250), .A(N5789), .B(N5788), .S0(N1135));
MXI2XL addgen2_A_I1531 (.Y(N1159), .A(N5874), .B(N5865), .S0(N4250));
MXI2XL addgen2_A_I1532 (.Y(N4259), .A(N5790), .B(N5789), .S0(N1135));
MXI2XL addgen2_A_I1533 (.Y(N1160), .A(N5874), .B(N5865), .S0(N4259));
MXI2XL addgen2_A_I1534 (.Y(N4268), .A(N5791), .B(N5790), .S0(N1135));
MXI2XL addgen2_A_I1535 (.Y(N1161), .A(N5874), .B(N5865), .S0(N4268));
MXI2XL addgen2_A_I1536 (.Y(N4277), .A(N5792), .B(N5791), .S0(N1135));
MXI2XL addgen2_A_I1537 (.Y(N1162), .A(N5874), .B(N5865), .S0(N4277));
NOR2BX1 addgen2_A_I1538 (.Y(N4286), .AN(N1135), .B(N5792));
MXI2XL addgen2_A_I1539 (.Y(N1163), .A(N5874), .B(N5865), .S0(N4286));
XNOR2X1 enc2_A_I1540 (.Y(N1167), .A(inst_cellmath__203_0_in0[7]), .B(inst_cellmath__203_0_in0[6]));
NAND2XL enc2_A_I1541 (.Y(N4295), .A(inst_cellmath__203_0_in0[7]), .B(inst_cellmath__203_0_in0[6]));
NOR2XL enc2_A_I1542 (.Y(N4297), .A(inst_cellmath__203_0_in0[7]), .B(inst_cellmath__203_0_in0[6]));
AND2XL enc2_A_I1543 (.Y(N1169), .A(N4295), .B(inst_cellmath__203_0_in0[8]));
OR2XL inst_cellmath__203_0_I2220 (.Y(N5891), .A(N4297), .B(inst_cellmath__203_0_in0[8]));
INVXL inst_cellmath__203_0_I2095 (.Y(N5900), .A(N1169));
NOR2XL addgen2_A_I1545 (.Y(N4308), .A(N5771), .B(N1167));
MXI2XL addgen2_A_I1546 (.Y(N1173), .A(N5900), .B(N5891), .S0(N4308));
MXI2XL addgen2_A_I1547 (.Y(N4317), .A(N5772), .B(N5771), .S0(N1167));
MXI2XL addgen2_A_I1548 (.Y(N1174), .A(N5900), .B(N5891), .S0(N4317));
MXI2XL addgen2_A_I1549 (.Y(N4326), .A(N5773), .B(N5772), .S0(N1167));
MXI2XL addgen2_A_I1550 (.Y(N1175), .A(N5900), .B(N5891), .S0(N4326));
MXI2XL addgen2_A_I1551 (.Y(N4335), .A(N5774), .B(N5773), .S0(N1167));
MXI2XL addgen2_A_I1552 (.Y(N1176), .A(N5900), .B(N5891), .S0(N4335));
MXI2XL addgen2_A_I1553 (.Y(N4344), .A(N5775), .B(N5774), .S0(N1167));
MXI2XL addgen2_A_I1554 (.Y(N1177), .A(N5900), .B(N5891), .S0(N4344));
MXI2XL addgen2_A_I1555 (.Y(N4353), .A(N5776), .B(N5775), .S0(N1167));
MXI2XL addgen2_A_I1556 (.Y(N1178), .A(N5900), .B(N5891), .S0(N4353));
MXI2XL addgen2_A_I1557 (.Y(N4362), .A(N5777), .B(N5776), .S0(N1167));
MXI2XL addgen2_A_I1558 (.Y(N1179), .A(N5900), .B(N5891), .S0(N4362));
MXI2XL addgen2_A_I1559 (.Y(N4371), .A(N5778), .B(N5777), .S0(N1167));
MXI2XL addgen2_A_I1560 (.Y(N1180), .A(N5900), .B(N5891), .S0(N4371));
MXI2XL addgen2_A_I1561 (.Y(N4380), .A(N5779), .B(N5778), .S0(N1167));
MXI2XL addgen2_A_I1562 (.Y(N1181), .A(N5900), .B(N5891), .S0(N4380));
MXI2XL addgen2_A_I1563 (.Y(N4389), .A(N5780), .B(N5779), .S0(N1167));
MXI2XL addgen2_A_I1564 (.Y(N1182), .A(N5900), .B(N5891), .S0(N4389));
MXI2XL addgen2_A_I1565 (.Y(N4398), .A(N5781), .B(N5780), .S0(N1167));
MXI2XL addgen2_A_I1566 (.Y(N1183), .A(N5900), .B(N5891), .S0(N4398));
MXI2XL addgen2_A_I1567 (.Y(N4407), .A(N5782), .B(N5781), .S0(N1167));
MXI2XL addgen2_A_I1568 (.Y(N1184), .A(N5900), .B(N5891), .S0(N4407));
MXI2XL addgen2_A_I1569 (.Y(N4416), .A(N5783), .B(N5782), .S0(N1167));
MXI2XL addgen2_A_I1570 (.Y(N1185), .A(N5900), .B(N5891), .S0(N4416));
MXI2XL addgen2_A_I1571 (.Y(N4425), .A(N5784), .B(N5783), .S0(N1167));
MXI2XL addgen2_A_I1572 (.Y(N1186), .A(N5900), .B(N5891), .S0(N4425));
MXI2XL addgen2_A_I1573 (.Y(N4434), .A(N5785), .B(N5784), .S0(N1167));
MXI2XL addgen2_A_I1574 (.Y(N1187), .A(N5900), .B(N5891), .S0(N4434));
MXI2XL addgen2_A_I1575 (.Y(N4443), .A(N5786), .B(N5785), .S0(N1167));
MXI2XL addgen2_A_I1576 (.Y(N1188), .A(N5900), .B(N5891), .S0(N4443));
MXI2XL addgen2_A_I1577 (.Y(N4452), .A(N5787), .B(N5786), .S0(N1167));
MXI2XL addgen2_A_I1578 (.Y(N1189), .A(N5900), .B(N5891), .S0(N4452));
MXI2XL addgen2_A_I1579 (.Y(N4461), .A(N5788), .B(N5787), .S0(N1167));
MXI2XL addgen2_A_I1580 (.Y(N1190), .A(N5900), .B(N5891), .S0(N4461));
MXI2XL addgen2_A_I1581 (.Y(N4470), .A(N5789), .B(N5788), .S0(N1167));
MXI2XL addgen2_A_I1582 (.Y(N1191), .A(N5900), .B(N5891), .S0(N4470));
MXI2XL addgen2_A_I1583 (.Y(N4479), .A(N5790), .B(N5789), .S0(N1167));
MXI2XL addgen2_A_I1584 (.Y(N1192), .A(N5900), .B(N5891), .S0(N4479));
MXI2XL addgen2_A_I1585 (.Y(N4488), .A(N5791), .B(N5790), .S0(N1167));
MXI2XL addgen2_A_I1586 (.Y(N1193), .A(N5900), .B(N5891), .S0(N4488));
MXI2XL addgen2_A_I1587 (.Y(N4497), .A(N5792), .B(N5791), .S0(N1167));
MXI2XL addgen2_A_I1588 (.Y(N1194), .A(N5900), .B(N5891), .S0(N4497));
NOR2BX1 addgen2_A_I1589 (.Y(N4506), .AN(N1167), .B(N5792));
MXI2XL addgen2_A_I1590 (.Y(N1195), .A(N5900), .B(N5891), .S0(N4506));
XNOR2X1 enc2_A_I1591 (.Y(N1199), .A(inst_cellmath__203_0_in0[9]), .B(inst_cellmath__203_0_in0[8]));
NAND2XL enc2_A_I1592 (.Y(N4515), .A(inst_cellmath__203_0_in0[9]), .B(inst_cellmath__203_0_in0[8]));
NOR2XL enc2_A_I1593 (.Y(N4517), .A(inst_cellmath__203_0_in0[9]), .B(inst_cellmath__203_0_in0[8]));
AND2XL enc2_A_I1594 (.Y(N1201), .A(N4515), .B(inst_cellmath__203_0_in0[10]));
OR2XL inst_cellmath__203_0_I2222 (.Y(N5917), .A(N4517), .B(inst_cellmath__203_0_in0[10]));
INVXL inst_cellmath__203_0_I2121 (.Y(N5926), .A(N1201));
NOR2XL addgen2_A_I1596 (.Y(N4528), .A(N5771), .B(N1199));
MXI2XL addgen2_A_I1597 (.Y(N1205), .A(N5926), .B(N5917), .S0(N4528));
MXI2XL addgen2_A_I1598 (.Y(N4537), .A(N5772), .B(N5771), .S0(N1199));
MXI2XL addgen2_A_I1599 (.Y(N1206), .A(N5926), .B(N5917), .S0(N4537));
MXI2XL addgen2_A_I1600 (.Y(N4546), .A(N5773), .B(N5772), .S0(N1199));
MXI2XL addgen2_A_I1601 (.Y(N1207), .A(N5926), .B(N5917), .S0(N4546));
MXI2XL addgen2_A_I1602 (.Y(N4555), .A(N5774), .B(N5773), .S0(N1199));
MXI2XL addgen2_A_I1603 (.Y(N1208), .A(N5926), .B(N5917), .S0(N4555));
MXI2XL addgen2_A_I1604 (.Y(N4564), .A(N5775), .B(N5774), .S0(N1199));
MXI2XL addgen2_A_I1605 (.Y(N1209), .A(N5926), .B(N5917), .S0(N4564));
MXI2XL addgen2_A_I1606 (.Y(N4573), .A(N5776), .B(N5775), .S0(N1199));
MXI2XL addgen2_A_I1607 (.Y(N1210), .A(N5926), .B(N5917), .S0(N4573));
MXI2XL addgen2_A_I1608 (.Y(N4582), .A(N5777), .B(N5776), .S0(N1199));
MXI2XL addgen2_A_I1609 (.Y(N1211), .A(N5926), .B(N5917), .S0(N4582));
MXI2XL addgen2_A_I1610 (.Y(N4591), .A(N5778), .B(N5777), .S0(N1199));
MXI2XL addgen2_A_I1611 (.Y(N1212), .A(N5926), .B(N5917), .S0(N4591));
MXI2XL addgen2_A_I1612 (.Y(N4600), .A(N5779), .B(N5778), .S0(N1199));
MXI2XL addgen2_A_I1613 (.Y(N1213), .A(N5926), .B(N5917), .S0(N4600));
MXI2XL addgen2_A_I1614 (.Y(N4609), .A(N5780), .B(N5779), .S0(N1199));
MXI2XL addgen2_A_I1615 (.Y(N1214), .A(N5926), .B(N5917), .S0(N4609));
MXI2XL addgen2_A_I1616 (.Y(N4618), .A(N5781), .B(N5780), .S0(N1199));
MXI2XL addgen2_A_I1617 (.Y(N1215), .A(N5926), .B(N5917), .S0(N4618));
MXI2XL addgen2_A_I1618 (.Y(N4627), .A(N5782), .B(N5781), .S0(N1199));
MXI2XL addgen2_A_I1619 (.Y(N1216), .A(N5926), .B(N5917), .S0(N4627));
MXI2XL addgen2_A_I1620 (.Y(N4636), .A(N5783), .B(N5782), .S0(N1199));
MXI2XL addgen2_A_I1621 (.Y(N1217), .A(N5926), .B(N5917), .S0(N4636));
MXI2XL addgen2_A_I1622 (.Y(N4645), .A(N5784), .B(N5783), .S0(N1199));
MXI2XL addgen2_A_I1623 (.Y(N1218), .A(N5926), .B(N5917), .S0(N4645));
MXI2XL addgen2_A_I1624 (.Y(N4654), .A(N5785), .B(N5784), .S0(N1199));
MXI2XL addgen2_A_I1625 (.Y(N1219), .A(N5926), .B(N5917), .S0(N4654));
MXI2XL addgen2_A_I1626 (.Y(N4663), .A(N5786), .B(N5785), .S0(N1199));
MXI2XL addgen2_A_I1627 (.Y(N1220), .A(N5926), .B(N5917), .S0(N4663));
MXI2XL addgen2_A_I1628 (.Y(N4672), .A(N5787), .B(N5786), .S0(N1199));
MXI2XL addgen2_A_I1629 (.Y(N1221), .A(N5926), .B(N5917), .S0(N4672));
MXI2XL addgen2_A_I1630 (.Y(N4681), .A(N5788), .B(N5787), .S0(N1199));
MXI2XL addgen2_A_I1631 (.Y(N1222), .A(N5926), .B(N5917), .S0(N4681));
MXI2XL addgen2_A_I1632 (.Y(N4690), .A(N5789), .B(N5788), .S0(N1199));
MXI2XL addgen2_A_I1633 (.Y(N1223), .A(N5926), .B(N5917), .S0(N4690));
MXI2XL addgen2_A_I1634 (.Y(N4699), .A(N5790), .B(N5789), .S0(N1199));
MXI2XL addgen2_A_I1635 (.Y(N1224), .A(N5926), .B(N5917), .S0(N4699));
MXI2XL addgen2_A_I1636 (.Y(N4708), .A(N5791), .B(N5790), .S0(N1199));
MXI2XL addgen2_A_I1637 (.Y(N1225), .A(N5926), .B(N5917), .S0(N4708));
MXI2XL addgen2_A_I1638 (.Y(N4717), .A(N5792), .B(N5791), .S0(N1199));
MXI2XL addgen2_A_I1639 (.Y(N1226), .A(N5926), .B(N5917), .S0(N4717));
NOR2BX1 addgen2_A_I1640 (.Y(N4726), .AN(N1199), .B(N5792));
MXI2XL addgen2_A_I1641 (.Y(N1227), .A(N5926), .B(N5917), .S0(N4726));
XNOR2X1 enc2_A_I1642 (.Y(N1231), .A(inst_cellmath__203_0_in0[11]), .B(inst_cellmath__203_0_in0[10]));
NAND2XL enc2_A_I1643 (.Y(N4735), .A(inst_cellmath__203_0_in0[11]), .B(inst_cellmath__203_0_in0[10]));
NOR2XL enc2_A_I1644 (.Y(N4737), .A(inst_cellmath__203_0_in0[11]), .B(inst_cellmath__203_0_in0[10]));
AND2XL enc2_A_I1645 (.Y(N1233), .A(N4735), .B(inst_cellmath__203_0_in0[12]));
OR2XL inst_cellmath__203_0_I2223 (.Y(N5941), .A(N4737), .B(inst_cellmath__203_0_in0[12]));
INVXL inst_cellmath__203_0_I2144 (.Y(N5949), .A(N1233));
NOR2XL addgen2_A_I1647 (.Y(N4748), .A(N5771), .B(N1231));
MXI2XL addgen2_A_I1648 (.Y(N1237), .A(N5949), .B(N5941), .S0(N4748));
MXI2XL addgen2_A_I1649 (.Y(N4757), .A(N5772), .B(N5771), .S0(N1231));
MXI2XL addgen2_A_I1650 (.Y(N1238), .A(N5949), .B(N5941), .S0(N4757));
MXI2XL addgen2_A_I1651 (.Y(N4766), .A(N5773), .B(N5772), .S0(N1231));
MXI2XL addgen2_A_I1652 (.Y(N1239), .A(N5949), .B(N5941), .S0(N4766));
MXI2XL addgen2_A_I1653 (.Y(N4775), .A(N5774), .B(N5773), .S0(N1231));
MXI2XL addgen2_A_I1654 (.Y(N1240), .A(N5949), .B(N5941), .S0(N4775));
MXI2XL addgen2_A_I1655 (.Y(N4784), .A(N5775), .B(N5774), .S0(N1231));
MXI2XL addgen2_A_I1656 (.Y(N1241), .A(N5949), .B(N5941), .S0(N4784));
MXI2XL addgen2_A_I1657 (.Y(N4793), .A(N5776), .B(N5775), .S0(N1231));
MXI2XL addgen2_A_I1658 (.Y(N1242), .A(N5949), .B(N5941), .S0(N4793));
MXI2XL addgen2_A_I1659 (.Y(N4802), .A(N5777), .B(N5776), .S0(N1231));
MXI2XL addgen2_A_I1660 (.Y(N1243), .A(N5949), .B(N5941), .S0(N4802));
MXI2XL addgen2_A_I1661 (.Y(N4811), .A(N5778), .B(N5777), .S0(N1231));
MXI2XL addgen2_A_I1662 (.Y(N1244), .A(N5949), .B(N5941), .S0(N4811));
MXI2XL addgen2_A_I1663 (.Y(N4820), .A(N5779), .B(N5778), .S0(N1231));
MXI2XL addgen2_A_I1664 (.Y(N1245), .A(N5949), .B(N5941), .S0(N4820));
MXI2XL addgen2_A_I1665 (.Y(N4829), .A(N5780), .B(N5779), .S0(N1231));
MXI2XL addgen2_A_I1666 (.Y(N1246), .A(N5949), .B(N5941), .S0(N4829));
MXI2XL addgen2_A_I1667 (.Y(N4838), .A(N5781), .B(N5780), .S0(N1231));
MXI2XL addgen2_A_I1668 (.Y(N1247), .A(N5949), .B(N5941), .S0(N4838));
MXI2XL addgen2_A_I1669 (.Y(N4847), .A(N5782), .B(N5781), .S0(N1231));
MXI2XL addgen2_A_I1670 (.Y(N1248), .A(N5949), .B(N5941), .S0(N4847));
MXI2XL addgen2_A_I1671 (.Y(N4856), .A(N5783), .B(N5782), .S0(N1231));
MXI2XL addgen2_A_I1672 (.Y(N1249), .A(N5949), .B(N5941), .S0(N4856));
MXI2XL addgen2_A_I1673 (.Y(N4865), .A(N5784), .B(N5783), .S0(N1231));
MXI2XL addgen2_A_I1674 (.Y(N1250), .A(N5949), .B(N5941), .S0(N4865));
MXI2XL addgen2_A_I1675 (.Y(N4874), .A(N5785), .B(N5784), .S0(N1231));
MXI2XL addgen2_A_I1676 (.Y(N1251), .A(N5949), .B(N5941), .S0(N4874));
MXI2XL addgen2_A_I1677 (.Y(N4883), .A(N5786), .B(N5785), .S0(N1231));
MXI2XL addgen2_A_I1678 (.Y(N1252), .A(N5949), .B(N5941), .S0(N4883));
MXI2XL addgen2_A_I1679 (.Y(N4892), .A(N5787), .B(N5786), .S0(N1231));
MXI2XL addgen2_A_I1680 (.Y(N1253), .A(N5949), .B(N5941), .S0(N4892));
MXI2XL addgen2_A_I1681 (.Y(N4901), .A(N5788), .B(N5787), .S0(N1231));
MXI2XL addgen2_A_I1682 (.Y(N1254), .A(N5949), .B(N5941), .S0(N4901));
MXI2XL addgen2_A_I1683 (.Y(N4910), .A(N5789), .B(N5788), .S0(N1231));
MXI2XL addgen2_A_I1684 (.Y(N1255), .A(N5949), .B(N5941), .S0(N4910));
MXI2XL addgen2_A_I1685 (.Y(N4919), .A(N5790), .B(N5789), .S0(N1231));
MXI2XL addgen2_A_I1686 (.Y(N1256), .A(N5949), .B(N5941), .S0(N4919));
MXI2XL addgen2_A_I1687 (.Y(N4928), .A(N5791), .B(N5790), .S0(N1231));
MXI2XL addgen2_A_I1688 (.Y(N1257), .A(N5949), .B(N5941), .S0(N4928));
MXI2XL addgen2_A_I1689 (.Y(N4937), .A(N5792), .B(N5791), .S0(N1231));
MXI2XL addgen2_A_I1690 (.Y(N1258), .A(N5949), .B(N5941), .S0(N4937));
NOR2BX1 addgen2_A_I1691 (.Y(N4946), .AN(N1231), .B(N5792));
MXI2XL addgen2_A_I1692 (.Y(N1259), .A(N5949), .B(N5941), .S0(N4946));
XNOR2X1 enc2_A_I1693 (.Y(N1263), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
NAND2XL enc2_A_I1694 (.Y(N4955), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
NOR2XL enc2_A_I1695 (.Y(N4957), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
AND2XL enc2_A_I1696 (.Y(N1265), .A(N4955), .B(inst_cellmath__203_0_in0[14]));
OR2XL inst_cellmath__203_0_I2225 (.Y(N5966), .A(N4957), .B(inst_cellmath__203_0_in0[14]));
INVXL inst_cellmath__203_0_I2169 (.Y(N5974), .A(N1265));
NOR2XL addgen2_A_I1698 (.Y(N4968), .A(N5771), .B(N1263));
MXI2XL addgen2_A_I1699 (.Y(N1269), .A(N5974), .B(N5966), .S0(N4968));
MXI2XL addgen2_A_I1700 (.Y(N4977), .A(N5772), .B(N5771), .S0(N1263));
MXI2XL addgen2_A_I1701 (.Y(N1270), .A(N5974), .B(N5966), .S0(N4977));
MXI2XL addgen2_A_I1702 (.Y(N4986), .A(N5773), .B(N5772), .S0(N1263));
MXI2XL addgen2_A_I1703 (.Y(N1271), .A(N5974), .B(N5966), .S0(N4986));
MXI2XL addgen2_A_I1704 (.Y(N4995), .A(N5774), .B(N5773), .S0(N1263));
MXI2XL addgen2_A_I1705 (.Y(N1272), .A(N5974), .B(N5966), .S0(N4995));
MXI2XL addgen2_A_I1706 (.Y(N5004), .A(N5775), .B(N5774), .S0(N1263));
MXI2XL addgen2_A_I1707 (.Y(N1273), .A(N5974), .B(N5966), .S0(N5004));
MXI2XL addgen2_A_I1708 (.Y(N5013), .A(N5776), .B(N5775), .S0(N1263));
MXI2XL addgen2_A_I1709 (.Y(N1274), .A(N5974), .B(N5966), .S0(N5013));
MXI2XL addgen2_A_I1710 (.Y(N5022), .A(N5777), .B(N5776), .S0(N1263));
MXI2XL addgen2_A_I1711 (.Y(N1275), .A(N5974), .B(N5966), .S0(N5022));
MXI2XL addgen2_A_I1712 (.Y(N5031), .A(N5778), .B(N5777), .S0(N1263));
MXI2XL addgen2_A_I1713 (.Y(N1276), .A(N5974), .B(N5966), .S0(N5031));
MXI2XL addgen2_A_I1714 (.Y(N5040), .A(N5779), .B(N5778), .S0(N1263));
MXI2XL addgen2_A_I1715 (.Y(N1277), .A(N5974), .B(N5966), .S0(N5040));
MXI2XL addgen2_A_I1716 (.Y(N5049), .A(N5780), .B(N5779), .S0(N1263));
MXI2XL addgen2_A_I1717 (.Y(N1278), .A(N5974), .B(N5966), .S0(N5049));
MXI2XL addgen2_A_I1718 (.Y(N5058), .A(N5781), .B(N5780), .S0(N1263));
MXI2XL addgen2_A_I1719 (.Y(N1279), .A(N5974), .B(N5966), .S0(N5058));
MXI2XL addgen2_A_I1720 (.Y(N5067), .A(N5782), .B(N5781), .S0(N1263));
MXI2XL addgen2_A_I1721 (.Y(N1280), .A(N5974), .B(N5966), .S0(N5067));
MXI2XL addgen2_A_I1722 (.Y(N5076), .A(N5783), .B(N5782), .S0(N1263));
MXI2XL addgen2_A_I1723 (.Y(N1281), .A(N5974), .B(N5966), .S0(N5076));
MXI2XL addgen2_A_I1724 (.Y(N5085), .A(N5784), .B(N5783), .S0(N1263));
MXI2XL addgen2_A_I1725 (.Y(N1282), .A(N5974), .B(N5966), .S0(N5085));
MXI2XL addgen2_A_I1726 (.Y(N5094), .A(N5785), .B(N5784), .S0(N1263));
MXI2XL addgen2_A_I1727 (.Y(N1283), .A(N5974), .B(N5966), .S0(N5094));
MXI2XL addgen2_A_I1728 (.Y(N5103), .A(N5786), .B(N5785), .S0(N1263));
MXI2XL addgen2_A_I1729 (.Y(N1284), .A(N5974), .B(N5966), .S0(N5103));
MXI2XL addgen2_A_I1730 (.Y(N5112), .A(N5787), .B(N5786), .S0(N1263));
MXI2XL addgen2_A_I1731 (.Y(N1285), .A(N5974), .B(N5966), .S0(N5112));
MXI2XL addgen2_A_I1732 (.Y(N5121), .A(N5788), .B(N5787), .S0(N1263));
MXI2XL addgen2_A_I1733 (.Y(N1286), .A(N5974), .B(N5966), .S0(N5121));
MXI2XL addgen2_A_I1734 (.Y(N5130), .A(N5789), .B(N5788), .S0(N1263));
MXI2XL addgen2_A_I1735 (.Y(N1287), .A(N5974), .B(N5966), .S0(N5130));
MXI2XL addgen2_A_I1736 (.Y(N5139), .A(N5790), .B(N5789), .S0(N1263));
MXI2XL addgen2_A_I1737 (.Y(N1288), .A(N5974), .B(N5966), .S0(N5139));
MXI2XL addgen2_A_I1738 (.Y(N5148), .A(N5791), .B(N5790), .S0(N1263));
MXI2XL addgen2_A_I1739 (.Y(N1289), .A(N5974), .B(N5966), .S0(N5148));
MXI2XL addgen2_A_I1740 (.Y(N5157), .A(N5792), .B(N5791), .S0(N1263));
MXI2XL addgen2_A_I1741 (.Y(N1290), .A(N5974), .B(N5966), .S0(N5157));
NOR2BX1 addgen2_A_I1742 (.Y(N5166), .AN(N1263), .B(N5792));
MXI2XL addgen2_A_I1743 (.Y(N2112), .A(N5974), .B(N5966), .S0(N5166));
XNOR2X1 enc2_A_I1744 (.Y(N1295), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
NAND2XL enc2_A_I1745 (.Y(N5175), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
NOR2XL enc2_A_I1746 (.Y(N5177), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
AND2XL enc2_A_I1747 (.Y(N1297), .A(N5175), .B(inst_cellmath__203_0_in4[0]));
OR2XL inst_cellmath__203_0_I2226 (.Y(N5989), .A(N5177), .B(inst_cellmath__203_0_in4[0]));
INVXL inst_cellmath__203_0_I2192 (.Y(inst_cellmath__203_0_out1[42]), .A(N1297));
NOR2XL addgen2_A_I1749 (.Y(N5188), .A(N5771), .B(N1295));
MXI2XL addgen2_A_I1750 (.Y(N1301), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5188));
MXI2XL addgen2_A_I1751 (.Y(N5197), .A(N5772), .B(N5771), .S0(N1295));
MXI2XL addgen2_A_I1752 (.Y(N1302), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5197));
MXI2XL addgen2_A_I1753 (.Y(N5206), .A(N5773), .B(N5772), .S0(N1295));
MXI2XL addgen2_A_I1754 (.Y(N1303), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5206));
MXI2XL addgen2_A_I1755 (.Y(N5215), .A(N5774), .B(N5773), .S0(N1295));
MXI2XL addgen2_A_I1756 (.Y(N1304), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5215));
MXI2XL addgen2_A_I1757 (.Y(N5224), .A(N5775), .B(N5774), .S0(N1295));
MXI2XL addgen2_A_I1758 (.Y(N1305), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5224));
MXI2XL addgen2_A_I1759 (.Y(N5233), .A(N5776), .B(N5775), .S0(N1295));
MXI2XL addgen2_A_I1760 (.Y(N1306), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5233));
MXI2XL addgen2_A_I1761 (.Y(N5242), .A(N5777), .B(N5776), .S0(N1295));
MXI2XL addgen2_A_I1762 (.Y(N1307), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5242));
MXI2XL addgen2_A_I1763 (.Y(N5251), .A(N5778), .B(N5777), .S0(N1295));
MXI2XL addgen2_A_I1764 (.Y(N1308), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5251));
MXI2XL addgen2_A_I1765 (.Y(N5260), .A(N5779), .B(N5778), .S0(N1295));
MXI2XL addgen2_A_I1766 (.Y(N1309), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5260));
MXI2XL addgen2_A_I1767 (.Y(N5269), .A(N5780), .B(N5779), .S0(N1295));
MXI2XL addgen2_A_I1768 (.Y(N1310), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5269));
MXI2XL addgen2_A_I1769 (.Y(N5278), .A(N5781), .B(N5780), .S0(N1295));
MXI2XL addgen2_A_I1770 (.Y(N1311), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5278));
MXI2XL addgen2_A_I1771 (.Y(N5287), .A(N5782), .B(N5781), .S0(N1295));
MXI2XL addgen2_A_I1772 (.Y(N1312), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5287));
MXI2XL addgen2_A_I1773 (.Y(N5296), .A(N5783), .B(N5782), .S0(N1295));
MXI2XL addgen2_A_I1774 (.Y(N1313), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5296));
MXI2XL addgen2_A_I1775 (.Y(N5305), .A(N5784), .B(N5783), .S0(N1295));
MXI2XL addgen2_A_I1776 (.Y(N1314), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5305));
MXI2XL addgen2_A_I1777 (.Y(N5314), .A(N5785), .B(N5784), .S0(N1295));
MXI2XL addgen2_A_I1778 (.Y(N1315), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5314));
MXI2XL addgen2_A_I1779 (.Y(N5323), .A(N5786), .B(N5785), .S0(N1295));
MXI2XL addgen2_A_I1780 (.Y(N1316), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5323));
MXI2XL addgen2_A_I1781 (.Y(N5332), .A(N5787), .B(N5786), .S0(N1295));
MXI2XL addgen2_A_I1782 (.Y(N1317), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5332));
MXI2XL addgen2_A_I1783 (.Y(N5341), .A(N5788), .B(N5787), .S0(N1295));
MXI2XL addgen2_A_I1784 (.Y(N1318), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5341));
MXI2XL addgen2_A_I1785 (.Y(N5350), .A(N5789), .B(N5788), .S0(N1295));
MXI2XL addgen2_A_I1786 (.Y(N1319), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5350));
MXI2XL addgen2_A_I1787 (.Y(N5359), .A(N5790), .B(N5789), .S0(N1295));
MXI2XL addgen2_A_I1788 (.Y(N1320), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5359));
MXI2XL addgen2_A_I1789 (.Y(N5368), .A(N5791), .B(N5790), .S0(N1295));
MXI2XL addgen2_A_I1790 (.Y(N1321), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5368));
MXI2XL addgen2_A_I1791 (.Y(N5377), .A(N5792), .B(N5791), .S0(N1295));
MXI2XL addgen2_A_I1792 (.Y(N1322), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5377));
NOR2BX1 addgen2_A_I1793 (.Y(N5386), .AN(N1295), .B(N5792));
MXI2XL addgen2_A_I1794 (.Y(inst_cellmath__203_0_out0[42]), .A(inst_cellmath__203_0_out1[42]), .B(N5989), .S0(N5386));
ADDHX1 inst_cellmath__203_0_I684 (.CO(N1376), .S(inst_cellmath__203_0_out1[1]), .A(N518), .B(inst_cellmath__203_0_in1[19]));
ADDHX1 inst_cellmath__203_0_I685 (.CO(N1378), .S(inst_cellmath__203_0_out0[2]), .A(N520), .B(N1376));
ADDHX1 inst_cellmath__203_0_I686 (.CO(N1380), .S(N1379), .A(N522), .B(N591));
ADDFX1 inst_cellmath__203_0_I687 (.CO(N1382), .S(inst_cellmath__203_0_out0[3]), .A(N1379), .B(N567), .CI(N1378));
ADDFX1 inst_cellmath__203_0_I688 (.CO(N1384), .S(inst_cellmath__203_0_out1[4]), .A(N524), .B(N1025), .CI(N568));
ADDFX1 inst_cellmath__203_0_I689 (.CO(N1386), .S(inst_cellmath__203_0_out0[4]), .A(N596), .B(N1380), .CI(N1382));
ADDFX1 inst_cellmath__203_0_I690 (.CO(N1388), .S(N1387), .A(N1027), .B(inst_cellmath__203_0_in0[2]), .CI(N1077));
ADDFX1 inst_cellmath__203_0_I691 (.CO(N1390), .S(N1389), .A(N526), .B(N1387), .CI(N621));
ADDFX1 inst_cellmath__203_0_I692 (.CO(N1392), .S(inst_cellmath__203_0_out1[5]), .A(N597), .B(N569), .CI(N625));
ADDFX1 inst_cellmath__203_0_I693 (.CO(inst_cellmath__203_0_out1[6]), .S(inst_cellmath__203_0_out0[5]), .A(N1384), .B(N1389), .CI(N1386));
ADDFX1 inst_cellmath__203_0_I694 (.CO(N1396), .S(N1395), .A(N1078), .B(N1029), .CI(N1388));
ADDFX1 inst_cellmath__203_0_I695 (.CO(N1398), .S(N1397), .A(N528), .B(N1395), .CI(N570));
ADDFX1 inst_cellmath__203_0_I696 (.CO(N1400), .S(N1399), .A(N598), .B(N1390), .CI(N626));
ADDFX1 inst_cellmath__203_0_I697 (.CO(inst_cellmath__203_0_out1[7]), .S(inst_cellmath__203_0_out0[6]), .A(N1392), .B(N1397), .CI(N1399));
ADDFX1 inst_cellmath__203_0_I698 (.CO(N1404), .S(N1403), .A(N1031), .B(N1105), .CI(N1109));
ADDFX1 inst_cellmath__203_0_I699 (.CO(N1406), .S(N1405), .A(N1403), .B(N1079), .CI(N1396));
ADDFX1 inst_cellmath__203_0_I700 (.CO(N1408), .S(N1407), .A(N1405), .B(N530), .CI(N651));
ADDFX1 inst_cellmath__203_0_I701 (.CO(N1410), .S(N1409), .A(N599), .B(N571), .CI(N627));
ADDFX1 inst_cellmath__203_0_I702 (.CO(N1412), .S(N1411), .A(N1407), .B(N655), .CI(N1398));
ADDFX1 inst_cellmath__203_0_I703 (.CO(inst_cellmath__203_0_out1[8]), .S(inst_cellmath__203_0_out0[7]), .A(N1409), .B(N1400), .CI(N1411));
ADDFX1 inst_cellmath__203_0_I704 (.CO(N1416), .S(N1415), .A(N1110), .B(N1033), .CI(N1080));
ADDFX1 inst_cellmath__203_0_I705 (.CO(N1418), .S(N1417), .A(N1415), .B(N1404), .CI(N1406));
ADDFX1 inst_cellmath__203_0_I706 (.CO(N1420), .S(N1419), .A(N1417), .B(N532), .CI(N572));
ADDFX1 inst_cellmath__203_0_I707 (.CO(N1422), .S(N1421), .A(N600), .B(N1408), .CI(N628));
ADDFX1 inst_cellmath__203_0_I708 (.CO(N1424), .S(N1423), .A(N1419), .B(N656), .CI(N1410));
ADDFX1 inst_cellmath__203_0_I709 (.CO(inst_cellmath__203_0_out1[9]), .S(inst_cellmath__203_0_out0[8]), .A(N1421), .B(N1412), .CI(N1423));
ADDFX1 inst_cellmath__203_0_I710 (.CO(N1428), .S(N1427), .A(N1035), .B(N1137), .CI(N1141));
ADDFX1 inst_cellmath__203_0_I711 (.CO(N1430), .S(N1429), .A(N1081), .B(N1111), .CI(N1416));
ADDFX1 inst_cellmath__203_0_I712 (.CO(N1432), .S(N1431), .A(N1429), .B(N1427), .CI(N534));
ADDFX1 inst_cellmath__203_0_I713 (.CO(N1434), .S(N1433), .A(N681), .B(N1418), .CI(N1431));
ADDFX1 inst_cellmath__203_0_I714 (.CO(N1436), .S(N1435), .A(N685), .B(N573), .CI(N601));
ADDFX1 inst_cellmath__203_0_I715 (.CO(N1438), .S(N1437), .A(N657), .B(N629), .CI(N1433));
ADDFX1 inst_cellmath__203_0_I716 (.CO(N1440), .S(N1439), .A(N1422), .B(N1420), .CI(N1435));
ADDFX1 inst_cellmath__203_0_I717 (.CO(inst_cellmath__203_0_out1[10]), .S(inst_cellmath__203_0_out0[9]), .A(N1424), .B(N1437), .CI(N1439));
ADDFX1 inst_cellmath__203_0_I718 (.CO(N1444), .S(N1443), .A(N1142), .B(N1037), .CI(N1112));
ADDFX1 inst_cellmath__203_0_I719 (.CO(N1446), .S(N1445), .A(N1428), .B(N1082), .CI(N1443));
ADDFX1 inst_cellmath__203_0_I720 (.CO(N1448), .S(N1447), .A(N1445), .B(N1430), .CI(N536));
ADDFX1 inst_cellmath__203_0_I721 (.CO(N1450), .S(N1449), .A(N1447), .B(N1432), .CI(N574));
ADDFX1 inst_cellmath__203_0_I722 (.CO(N1452), .S(N1451), .A(N1434), .B(N686), .CI(N602));
ADDFX1 inst_cellmath__203_0_I723 (.CO(N1454), .S(N1453), .A(N658), .B(N630), .CI(N1449));
ADDFX1 inst_cellmath__203_0_I724 (.CO(N1456), .S(N1455), .A(N1438), .B(N1436), .CI(N1451));
ADDFX1 inst_cellmath__203_0_I725 (.CO(inst_cellmath__203_0_out1[11]), .S(inst_cellmath__203_0_out0[10]), .A(N1440), .B(N1453), .CI(N1455));
ADDFX1 inst_cellmath__203_0_I726 (.CO(N1460), .S(N1459), .A(N1039), .B(N1169), .CI(N1173));
ADDFX1 inst_cellmath__203_0_I727 (.CO(N1462), .S(N1461), .A(N1113), .B(N1143), .CI(N1083));
ADDFX1 inst_cellmath__203_0_I728 (.CO(N1464), .S(N1463), .A(N1459), .B(N1444), .CI(N1461));
ADDFX1 inst_cellmath__203_0_I729 (.CO(N1466), .S(N1465), .A(N538), .B(N1446), .CI(N1463));
ADDFX1 inst_cellmath__203_0_I730 (.CO(N1468), .S(N1467), .A(N711), .B(N1448), .CI(N1465));
ADDFX1 inst_cellmath__203_0_I731 (.CO(N1470), .S(N1469), .A(N687), .B(N575), .CI(N603));
ADDFX1 inst_cellmath__203_0_I732 (.CO(N1472), .S(N1471), .A(N659), .B(N631), .CI(N715));
ADDFX1 inst_cellmath__203_0_I733 (.CO(N1474), .S(N1473), .A(N1467), .B(N1450), .CI(N1452));
ADDFX1 inst_cellmath__203_0_I734 (.CO(N1476), .S(N1475), .A(N1471), .B(N1469), .CI(N1454));
ADDFX1 inst_cellmath__203_0_I735 (.CO(inst_cellmath__203_0_out1[12]), .S(inst_cellmath__203_0_out0[11]), .A(N1456), .B(N1473), .CI(N1475));
ADDFX1 inst_cellmath__203_0_I736 (.CO(N1480), .S(N1479), .A(N1174), .B(N1041), .CI(N1144));
ADDFX1 inst_cellmath__203_0_I737 (.CO(N1482), .S(N1481), .A(N1084), .B(N1114), .CI(N1460));
ADDFX1 inst_cellmath__203_0_I738 (.CO(N1484), .S(N1483), .A(N1479), .B(N1462), .CI(N1481));
ADDFX1 inst_cellmath__203_0_I739 (.CO(N1486), .S(N1485), .A(N540), .B(N1464), .CI(N1483));
ADDFX1 inst_cellmath__203_0_I740 (.CO(N1488), .S(N1487), .A(N576), .B(N1466), .CI(N1485));
ADDFX1 inst_cellmath__203_0_I741 (.CO(N1490), .S(N1489), .A(N604), .B(N688), .CI(N632));
ADDFX1 inst_cellmath__203_0_I742 (.CO(N1492), .S(N1491), .A(N1468), .B(N660), .CI(N716));
ADDFX1 inst_cellmath__203_0_I743 (.CO(N1494), .S(N1493), .A(N1487), .B(N1470), .CI(N1472));
ADDFX1 inst_cellmath__203_0_I744 (.CO(N1496), .S(N1495), .A(N1491), .B(N1489), .CI(N1474));
ADDFX1 inst_cellmath__203_0_I745 (.CO(inst_cellmath__203_0_out1[13]), .S(inst_cellmath__203_0_out0[12]), .A(N1476), .B(N1493), .CI(N1495));
ADDFX1 inst_cellmath__203_0_I746 (.CO(N1500), .S(N1499), .A(N1043), .B(N1201), .CI(N1205));
ADDFX1 inst_cellmath__203_0_I747 (.CO(N1502), .S(N1501), .A(N1085), .B(N1175), .CI(N1145));
ADDFX1 inst_cellmath__203_0_I748 (.CO(N1504), .S(N1503), .A(N1480), .B(N1115), .CI(N1499));
ADDFX1 inst_cellmath__203_0_I749 (.CO(N1506), .S(N1505), .A(N1482), .B(N1501), .CI(N1503));
ADDFX1 inst_cellmath__203_0_I750 (.CO(N1508), .S(N1507), .A(N1484), .B(N542), .CI(N1505));
ADDFX1 inst_cellmath__203_0_I751 (.CO(N1510), .S(N1509), .A(N741), .B(N1486), .CI(N577));
ADDFX1 inst_cellmath__203_0_I752 (.CO(N1512), .S(N1511), .A(N1507), .B(N689), .CI(N605));
ADDFX1 inst_cellmath__203_0_I753 (.CO(N1514), .S(N1513), .A(N661), .B(N633), .CI(N717));
ADDFX1 inst_cellmath__203_0_I754 (.CO(N1516), .S(N1515), .A(N1488), .B(N745), .CI(N1509));
ADDFX1 inst_cellmath__203_0_I755 (.CO(N1518), .S(N1517), .A(N1492), .B(N1490), .CI(N1511));
ADDFX1 inst_cellmath__203_0_I756 (.CO(N1520), .S(N1519), .A(N1494), .B(N1513), .CI(N1515));
ADDFX1 inst_cellmath__203_0_I757 (.CO(inst_cellmath__203_0_out1[14]), .S(inst_cellmath__203_0_out0[13]), .A(N1517), .B(N1496), .CI(N1519));
ADDFX1 inst_cellmath__203_0_I758 (.CO(N1524), .S(N1523), .A(N1206), .B(N1045), .CI(N1176));
ADDFX1 inst_cellmath__203_0_I759 (.CO(N1526), .S(N1525), .A(N1086), .B(N1146), .CI(N1116));
ADDFX1 inst_cellmath__203_0_I760 (.CO(N1528), .S(N1527), .A(N1502), .B(N1500), .CI(N1523));
ADDFX1 inst_cellmath__203_0_I761 (.CO(N1530), .S(N1529), .A(N1504), .B(N1525), .CI(N1527));
ADDFX1 inst_cellmath__203_0_I762 (.CO(N1532), .S(N1531), .A(N1506), .B(N544), .CI(N1529));
ADDFX1 inst_cellmath__203_0_I763 (.CO(N1534), .S(N1533), .A(N1508), .B(N578), .CI(N690));
ADDFX1 inst_cellmath__203_0_I764 (.CO(N1536), .S(N1535), .A(N634), .B(N606), .CI(N662));
ADDFX1 inst_cellmath__203_0_I765 (.CO(N1538), .S(N1537), .A(N718), .B(N1531), .CI(N746));
ADDFX1 inst_cellmath__203_0_I766 (.CO(N1540), .S(N1539), .A(N1512), .B(N1510), .CI(N1514));
ADDFX1 inst_cellmath__203_0_I767 (.CO(N1542), .S(N1541), .A(N1535), .B(N1533), .CI(N1516));
ADDFX1 inst_cellmath__203_0_I768 (.CO(N1544), .S(N1543), .A(N1518), .B(N1537), .CI(N1539));
ADDFX1 inst_cellmath__203_0_I769 (.CO(inst_cellmath__203_0_out1[15]), .S(inst_cellmath__203_0_out0[14]), .A(N1520), .B(N1541), .CI(N1543));
ADDHX1 inst_cellmath__203_0_I770 (.CO(N1548), .S(N1547), .A(N1233), .B(N1047));
ADDFX1 inst_cellmath__203_0_I771 (.CO(N1550), .S(N1549), .A(N1547), .B(N1237), .CI(N1207));
ADDFX1 inst_cellmath__203_0_I772 (.CO(N1552), .S(N1551), .A(N1177), .B(N1117), .CI(N1147));
ADDFX1 inst_cellmath__203_0_I773 (.CO(N1554), .S(N1553), .A(N1524), .B(N1087), .CI(N1526));
ADDFX1 inst_cellmath__203_0_I774 (.CO(N1556), .S(N1555), .A(N1551), .B(N1549), .CI(N1528));
ADDFX1 inst_cellmath__203_0_I775 (.CO(N1558), .S(N1557), .A(N546), .B(N1553), .CI(N1530));
ADDFX1 inst_cellmath__203_0_I776 (.CO(N1560), .S(N1559), .A(N779), .B(N1555), .CI(N579));
ADDFX1 inst_cellmath__203_0_I777 (.CO(N1562), .S(N1561), .A(N1557), .B(N1532), .CI(N691));
ADDFX1 inst_cellmath__203_0_I778 (.CO(N1564), .S(N1563), .A(N635), .B(N607), .CI(N663));
ADDFX1 inst_cellmath__203_0_I779 (.CO(N1566), .S(N1565), .A(N747), .B(N719), .CI(N1534));
ADDFX1 inst_cellmath__203_0_I780 (.CO(N1568), .S(N1567), .A(N1536), .B(N1559), .CI(N1561));
ADDFX1 inst_cellmath__203_0_I781 (.CO(N1570), .S(N1569), .A(N1563), .B(N1538), .CI(N1540));
ADDFX1 inst_cellmath__203_0_I782 (.CO(N1572), .S(N1571), .A(N1567), .B(N1565), .CI(N1542));
ADDFX1 inst_cellmath__203_0_I783 (.CO(inst_cellmath__203_0_out1[16]), .S(inst_cellmath__203_0_out0[15]), .A(N1569), .B(N1544), .CI(N1571));
ADDFX1 inst_cellmath__203_0_I784 (.CO(N1576), .S(N1575), .A(N1548), .B(N1049), .CI(N1238));
ADDFX1 inst_cellmath__203_0_I785 (.CO(N1578), .S(N1577), .A(N1178), .B(N1208), .CI(N1148));
ADDFX1 inst_cellmath__203_0_I786 (.CO(N1580), .S(N1579), .A(N1088), .B(N1118), .CI(N1550));
ADDFX1 inst_cellmath__203_0_I787 (.CO(N1582), .S(N1581), .A(N1575), .B(N1552), .CI(N1577));
ADDFX1 inst_cellmath__203_0_I788 (.CO(N1584), .S(N1583), .A(N1579), .B(N1554), .CI(N548));
ADDFX1 inst_cellmath__203_0_I789 (.CO(N1586), .S(N1585), .A(N1556), .B(N1581), .CI(N1583));
ADDFX1 inst_cellmath__203_0_I790 (.CO(N1588), .S(N1587), .A(N580), .B(N1558), .CI(N781));
ADDFX1 inst_cellmath__203_0_I791 (.CO(N1590), .S(N1589), .A(N608), .B(N692), .CI(N636));
ADDFX1 inst_cellmath__203_0_I792 (.CO(N1592), .S(N1591), .A(N1585), .B(N664), .CI(N720));
ADDFX1 inst_cellmath__203_0_I793 (.CO(N1594), .S(N1593), .A(N1560), .B(N748), .CI(N1562));
ADDFX1 inst_cellmath__203_0_I794 (.CO(N1596), .S(N1595), .A(N1587), .B(N1564), .CI(N1589));
ADDFX1 inst_cellmath__203_0_I795 (.CO(N1598), .S(N1597), .A(N1566), .B(N1591), .CI(N1593));
ADDFX1 inst_cellmath__203_0_I796 (.CO(N1600), .S(N1599), .A(N1595), .B(N1568), .CI(N1570));
ADDFX1 inst_cellmath__203_0_I797 (.CO(inst_cellmath__203_0_out1[17]), .S(inst_cellmath__203_0_out0[16]), .A(N1572), .B(N1597), .CI(N1599));
ADDFX1 inst_cellmath__203_0_I798 (.CO(N1604), .S(N1603), .A(N1051), .B(N1265), .CI(N1269));
ADDFX1 inst_cellmath__203_0_I799 (.CO(N1606), .S(N1605), .A(N1239), .B(N1089), .CI(N1149));
ADDFX1 inst_cellmath__203_0_I800 (.CO(N1608), .S(N1607), .A(N1179), .B(N1209), .CI(N1119));
ADDFX1 inst_cellmath__203_0_I801 (.CO(N1610), .S(N1609), .A(N1603), .B(N1576), .CI(N1578));
ADDFX1 inst_cellmath__203_0_I802 (.CO(N1612), .S(N1611), .A(N1580), .B(N1605), .CI(N1607));
ADDFX1 inst_cellmath__203_0_I803 (.CO(N1614), .S(N1613), .A(N1609), .B(N1582), .CI(N550));
ADDFX1 inst_cellmath__203_0_I804 (.CO(N1616), .S(N1615), .A(N1584), .B(N1611), .CI(N1613));
ADDFX1 inst_cellmath__203_0_I805 (.CO(N1618), .S(N1617), .A(N783), .B(N581), .CI(N693));
ADDFX1 inst_cellmath__203_0_I806 (.CO(N1620), .S(N1619), .A(N609), .B(N1586), .CI(N637));
ADDFX1 inst_cellmath__203_0_I807 (.CO(N1622), .S(N1621), .A(N721), .B(N665), .CI(N1615));
ADDFX1 inst_cellmath__203_0_I808 (.CO(N1624), .S(N1623), .A(N1588), .B(N749), .CI(N1590));
ADDFX1 inst_cellmath__203_0_I809 (.CO(N1626), .S(N1625), .A(N1617), .B(N1592), .CI(N1619));
ADDFX1 inst_cellmath__203_0_I810 (.CO(N1628), .S(N1627), .A(N1621), .B(N1594), .CI(N1623));
ADDFX1 inst_cellmath__203_0_I811 (.CO(N1630), .S(N1629), .A(N1625), .B(N1596), .CI(N1598));
ADDFX1 inst_cellmath__203_0_I812 (.CO(inst_cellmath__203_0_out1[18]), .S(inst_cellmath__203_0_out0[17]), .A(N1600), .B(N1627), .CI(N1629));
ADDFX1 inst_cellmath__203_0_I813 (.CO(N1634), .S(N1633), .A(N1270), .B(N1053), .CI(N1240));
ADDFX1 inst_cellmath__203_0_I814 (.CO(N1636), .S(N1635), .A(N1210), .B(N1090), .CI(N1180));
ADDFX1 inst_cellmath__203_0_I815 (.CO(N1638), .S(N1637), .A(N1120), .B(N1150), .CI(N1604));
ADDFX1 inst_cellmath__203_0_I816 (.CO(N1640), .S(N1639), .A(N1608), .B(N1606), .CI(N1633));
ADDFX1 inst_cellmath__203_0_I817 (.CO(N1642), .S(N1641), .A(N1637), .B(N1635), .CI(N1610));
ADDFX1 inst_cellmath__203_0_I818 (.CO(N1644), .S(N1643), .A(N1639), .B(N552), .CI(N1612));
ADDFX1 inst_cellmath__203_0_I819 (.CO(N1646), .S(N1645), .A(N1614), .B(N1641), .CI(N1643));
ADDFX1 inst_cellmath__203_0_I820 (.CO(N1648), .S(N1647), .A(N785), .B(N582), .CI(N694));
ADDFX1 inst_cellmath__203_0_I821 (.CO(N1650), .S(N1649), .A(N610), .B(N1616), .CI(N638));
ADDFX1 inst_cellmath__203_0_I822 (.CO(N1652), .S(N1651), .A(N722), .B(N666), .CI(N750));
ADDFX1 inst_cellmath__203_0_I823 (.CO(N1654), .S(N1653), .A(N1618), .B(N1645), .CI(N1620));
ADDFX1 inst_cellmath__203_0_I824 (.CO(N1656), .S(N1655), .A(N1622), .B(N1647), .CI(N1649));
ADDFX1 inst_cellmath__203_0_I825 (.CO(N1658), .S(N1657), .A(N1624), .B(N1651), .CI(N1653));
ADDFX1 inst_cellmath__203_0_I826 (.CO(N1660), .S(N1659), .A(N1655), .B(N1626), .CI(N1628));
ADDFX1 inst_cellmath__203_0_I827 (.CO(inst_cellmath__203_0_out1[19]), .S(inst_cellmath__203_0_out0[18]), .A(N1630), .B(N1657), .CI(N1659));
ADDFX1 inst_cellmath__203_0_I828 (.CO(N1664), .S(N1663), .A(N1055), .B(N1297), .CI(N1301));
ADDFX1 inst_cellmath__203_0_I829 (.CO(N1666), .S(N1665), .A(N1271), .B(N1121), .CI(N1181));
ADDFX1 inst_cellmath__203_0_I830 (.CO(N1668), .S(N1667), .A(N1241), .B(N1091), .CI(N1211));
ADDFX1 inst_cellmath__203_0_I831 (.CO(N1670), .S(N1669), .A(N1634), .B(N1151), .CI(N1663));
ADDFX1 inst_cellmath__203_0_I832 (.CO(N1672), .S(N1671), .A(N1665), .B(N1636), .CI(N1638));
ADDFX1 inst_cellmath__203_0_I833 (.CO(N1674), .S(N1673), .A(N1640), .B(N1667), .CI(N1669));
ADDFX1 inst_cellmath__203_0_I834 (.CO(N1676), .S(N1675), .A(N1671), .B(N554), .CI(N1642));
ADDFX1 inst_cellmath__203_0_I835 (.CO(N1678), .S(N1677), .A(N1644), .B(N1673), .CI(N1675));
ADDFX1 inst_cellmath__203_0_I836 (.CO(N1680), .S(N1679), .A(N787), .B(N583), .CI(N695));
ADDFX1 inst_cellmath__203_0_I837 (.CO(N1682), .S(N1681), .A(N1646), .B(N611), .CI(N667));
ADDFX1 inst_cellmath__203_0_I838 (.CO(N1684), .S(N1683), .A(N751), .B(N639), .CI(N723));
ADDFX1 inst_cellmath__203_0_I839 (.CO(N1686), .S(N1685), .A(N1648), .B(N1677), .CI(N1650));
ADDFX1 inst_cellmath__203_0_I840 (.CO(N1688), .S(N1687), .A(N1652), .B(N1679), .CI(N1681));
ADDFX1 inst_cellmath__203_0_I841 (.CO(N1690), .S(N1689), .A(N1654), .B(N1683), .CI(N1685));
ADDFX1 inst_cellmath__203_0_I842 (.CO(N1692), .S(N1691), .A(N1687), .B(N1656), .CI(N1658));
ADDFX1 inst_cellmath__203_0_I843 (.CO(inst_cellmath__203_0_out1[20]), .S(inst_cellmath__203_0_out0[19]), .A(N1660), .B(N1689), .CI(N1691));
INVXL fap1_A_I1795 (.Y(N5395), .A(N1732));
ADDFX1 fap1_A_I1796 (.CO(N1696), .S(N1695), .A(N1092), .B(N1302), .CI(N5395));
ADDFX1 inst_cellmath__203_0_I845 (.CO(N1700), .S(N1699), .A(N1272), .B(N1122), .CI(N1242));
ADDFX1 inst_cellmath__203_0_I846 (.CO(N1702), .S(N1701), .A(N1212), .B(N1182), .CI(N1152));
ADDFX1 inst_cellmath__203_0_I847 (.CO(N1704), .S(N1703), .A(N1666), .B(N1664), .CI(N1668));
ADDFX1 inst_cellmath__203_0_I848 (.CO(N1706), .S(N1705), .A(N1695), .B(N1699), .CI(N1701));
ADDFX1 inst_cellmath__203_0_I849 (.CO(N1708), .S(N1707), .A(N1672), .B(N1670), .CI(N1703));
ADDFX1 inst_cellmath__203_0_I850 (.CO(N1710), .S(N1709), .A(N1705), .B(N5654), .CI(N1674));
ADDFX1 inst_cellmath__203_0_I851 (.CO(N1712), .S(N1711), .A(N1707), .B(N1676), .CI(N584));
ADDFX1 inst_cellmath__203_0_I852 (.CO(N1714), .S(N1713), .A(N789), .B(N1709), .CI(N696));
ADDFX1 inst_cellmath__203_0_I853 (.CO(N1716), .S(N1715), .A(N640), .B(N612), .CI(N668));
ADDFX1 inst_cellmath__203_0_I854 (.CO(N1718), .S(N1717), .A(N724), .B(N1678), .CI(N752));
ADDFX1 inst_cellmath__203_0_I855 (.CO(N1720), .S(N1719), .A(N1711), .B(N1680), .CI(N1682));
ADDFX1 inst_cellmath__203_0_I856 (.CO(N1722), .S(N1721), .A(N1684), .B(N1713), .CI(N1715));
ADDFX1 inst_cellmath__203_0_I857 (.CO(N1724), .S(N1723), .A(N1686), .B(N1717), .CI(N1719));
ADDFX1 inst_cellmath__203_0_I858 (.CO(N1726), .S(N1725), .A(N1721), .B(N1688), .CI(N1690));
ADDFX1 inst_cellmath__203_0_I859 (.CO(inst_cellmath__203_0_out1[21]), .S(inst_cellmath__203_0_out0[20]), .A(N1692), .B(N1723), .CI(N1725));
ADDFX1 inst_cellmath__203_0_I1798 (.CO(N1730), .S(N1729), .A(N1093), .B(N1059), .CI(N5395));
ADDFX1 inst_cellmath__203_0_I861 (.CO(N1734), .S(N1733), .A(N1303), .B(N1153), .CI(N1213));
ADDFX1 inst_cellmath__203_0_I862 (.CO(N1736), .S(N1735), .A(N1273), .B(N1123), .CI(N1243));
ADDFX1 inst_cellmath__203_0_I863 (.CO(N1738), .S(N1737), .A(N1696), .B(N1183), .CI(N1700));
ADDFX1 inst_cellmath__203_0_I864 (.CO(N1740), .S(N1739), .A(N1733), .B(N1702), .CI(N1729));
ADDFX1 inst_cellmath__203_0_I865 (.CO(N1742), .S(N1741), .A(N1704), .B(N1735), .CI(N1737));
ADDFX1 inst_cellmath__203_0_I866 (.CO(N1744), .S(N1743), .A(N1739), .B(N1706), .CI(N1708));
ADDFX1 inst_cellmath__203_0_I867 (.CO(N1746), .S(N1745), .A(N1710), .B(N1741), .CI(N585));
ADDFX1 inst_cellmath__203_0_I868 (.CO(N1748), .S(N1747), .A(N1743), .B(N791), .CI(N697));
ADDFX1 inst_cellmath__203_0_I869 (.CO(N1750), .S(N1749), .A(N641), .B(N613), .CI(N669));
ADDFX1 inst_cellmath__203_0_I870 (.CO(N1752), .S(N1751), .A(N753), .B(N725), .CI(N1712));
ADDFX1 inst_cellmath__203_0_I871 (.CO(N1754), .S(N1753), .A(N1745), .B(N1714), .CI(N1716));
ADDFX1 inst_cellmath__203_0_I872 (.CO(N1756), .S(N1755), .A(N1718), .B(N1747), .CI(N1749));
ADDFX1 inst_cellmath__203_0_I873 (.CO(N1758), .S(N1757), .A(N1751), .B(N1720), .CI(N1753));
ADDFXL inst_cellmath__203_0_I874 (.CO(N1760), .S(N1759), .A(N1755), .B(N1722), .CI(N1724));
ADDFXL inst_cellmath__203_0_I875 (.CO(inst_cellmath__203_0_out1[22]), .S(inst_cellmath__203_0_out0[21]), .A(N1726), .B(N1757), .CI(N1759));
ADDFX1 inst_cellmath__203_0_I876 (.CO(N1764), .S(N1763), .A(N1061), .B(N1732), .CI(N1124));
ADDFX1 inst_cellmath__203_0_I877 (.CO(N1766), .S(N1765), .A(N1304), .B(N1154), .CI(N1274));
ADDFX1 inst_cellmath__203_0_I878 (.CO(N1768), .S(N1767), .A(N1244), .B(N1214), .CI(N1184));
ADDFX1 inst_cellmath__203_0_I879 (.CO(N1770), .S(N1769), .A(N1734), .B(N1094), .CI(N1730));
ADDFX1 inst_cellmath__203_0_I880 (.CO(N1772), .S(N1771), .A(N1763), .B(N1736), .CI(N1765));
ADDFX1 inst_cellmath__203_0_I881 (.CO(N1774), .S(N1773), .A(N1738), .B(N1767), .CI(N1769));
ADDFX1 inst_cellmath__203_0_I882 (.CO(N1776), .S(N1775), .A(N1771), .B(N1740), .CI(N1742));
ADDFX1 inst_cellmath__203_0_I883 (.CO(N1778), .S(N1777), .A(N5670), .B(N1773), .CI(N1744));
ADDFX1 inst_cellmath__203_0_I884 (.CO(N1780), .S(N1779), .A(N793), .B(N1775), .CI(N698));
ADDFX1 inst_cellmath__203_0_I885 (.CO(N1782), .S(N1781), .A(N642), .B(N614), .CI(N670));
ADDFX1 inst_cellmath__203_0_I886 (.CO(N1784), .S(N1783), .A(N754), .B(N726), .CI(N1746));
ADDFX1 inst_cellmath__203_0_I887 (.CO(N1786), .S(N1785), .A(N1748), .B(N1777), .CI(N1750));
ADDFX1 inst_cellmath__203_0_I888 (.CO(N1788), .S(N1787), .A(N1781), .B(N1779), .CI(N1752));
ADDFX1 inst_cellmath__203_0_I889 (.CO(N1790), .S(N1789), .A(N1783), .B(N1754), .CI(N1785));
ADDFX1 inst_cellmath__203_0_I890 (.CO(N1792), .S(N1791), .A(N1787), .B(N1756), .CI(N1758));
ADDFXL inst_cellmath__203_0_I891 (.CO(inst_cellmath__203_0_out1[23]), .S(inst_cellmath__203_0_out0[22]), .A(N1760), .B(N1789), .CI(N1791));
INVXL fap1_A_I1799 (.Y(N5413), .A(N1798));
ADDFX1 fap1_A_I1800 (.CO(N1796), .S(N1795), .A(N1155), .B(N1125), .CI(N5413));
ADDFX1 inst_cellmath__203_0_I893 (.CO(N1800), .S(N1799), .A(N1245), .B(N1185), .CI(N1305));
ADDFX1 inst_cellmath__203_0_I894 (.CO(N1802), .S(N1801), .A(N1275), .B(N1095), .CI(N1215));
ADDFX1 inst_cellmath__203_0_I895 (.CO(N1804), .S(N1803), .A(N1766), .B(N1764), .CI(N1768));
ADDFX1 inst_cellmath__203_0_I896 (.CO(N1806), .S(N1805), .A(N1795), .B(N1799), .CI(N1801));
ADDFX1 inst_cellmath__203_0_I897 (.CO(N1808), .S(N1807), .A(N1772), .B(N1770), .CI(N1803));
ADDFX1 inst_cellmath__203_0_I898 (.CO(N1810), .S(N1809), .A(N1774), .B(N1805), .CI(N1807));
ADDFX1 inst_cellmath__203_0_I899 (.CO(N1812), .S(N1811), .A(N795), .B(N1776), .CI(N699));
ADDFX1 inst_cellmath__203_0_I900 (.CO(N1814), .S(N1813), .A(N643), .B(N615), .CI(N1778));
ADDFX1 inst_cellmath__203_0_I901 (.CO(N1816), .S(N1815), .A(N1809), .B(N671), .CI(N727));
ADDFX1 inst_cellmath__203_0_I902 (.CO(N1818), .S(N1817), .A(N1780), .B(N755), .CI(N1782));
ADDFX1 inst_cellmath__203_0_I903 (.CO(N1820), .S(N1819), .A(N1813), .B(N1811), .CI(N1815));
ADDFX1 inst_cellmath__203_0_I904 (.CO(N1822), .S(N1821), .A(N1786), .B(N1784), .CI(N1817));
ADDFX1 inst_cellmath__203_0_I905 (.CO(N1824), .S(N1823), .A(N1819), .B(N1788), .CI(N1790));
ADDFX1 inst_cellmath__203_0_I906 (.CO(inst_cellmath__203_0_out1[24]), .S(inst_cellmath__203_0_out0[23]), .A(N1792), .B(N1821), .CI(N1823));
INVXL fap1_A_I1801 (.Y(N5422), .A(N1830));
ADDFX1 fap1_A_I1802 (.CO(N1828), .S(N1827), .A(N1156), .B(N1798), .CI(N5422));
ADDFX1 inst_cellmath__203_0_I908 (.CO(N1832), .S(N1831), .A(N1306), .B(N1186), .CI(N1126));
ADDFX1 inst_cellmath__203_0_I909 (.CO(N1834), .S(N1833), .A(N1246), .B(N1096), .CI(N1276));
ADDFX1 inst_cellmath__203_0_I910 (.CO(N1836), .S(N1835), .A(N1796), .B(N1216), .CI(N1800));
ADDFX1 inst_cellmath__203_0_I911 (.CO(N1838), .S(N1837), .A(N1827), .B(N1802), .CI(N1833));
ADDFX1 inst_cellmath__203_0_I912 (.CO(N1840), .S(N1839), .A(N1804), .B(N1831), .CI(N1835));
ADDFX1 inst_cellmath__203_0_I913 (.CO(N1842), .S(N1841), .A(N1837), .B(N1806), .CI(N1808));
ADDFX1 inst_cellmath__203_0_I914 (.CO(N1844), .S(N1843), .A(N5687), .B(N1839), .CI(N797));
ADDFX1 inst_cellmath__203_0_I915 (.CO(N1846), .S(N1845), .A(N1810), .B(N1841), .CI(N700));
ADDFX1 inst_cellmath__203_0_I916 (.CO(N1848), .S(N1847), .A(N672), .B(N644), .CI(N728));
ADDFX1 inst_cellmath__203_0_I917 (.CO(N1850), .S(N1849), .A(N1812), .B(N756), .CI(N1843));
ADDFX1 inst_cellmath__203_0_I918 (.CO(N1852), .S(N1851), .A(N1816), .B(N1814), .CI(N1845));
ADDFX1 inst_cellmath__203_0_I919 (.CO(N1854), .S(N1853), .A(N1818), .B(N1847), .CI(N1849));
ADDFX1 inst_cellmath__203_0_I920 (.CO(N1856), .S(N1855), .A(N1851), .B(N1820), .CI(N1822));
ADDFXL inst_cellmath__203_0_I921 (.CO(inst_cellmath__203_0_out1[25]), .S(inst_cellmath__203_0_out0[24]), .A(N1824), .B(N1853), .CI(N1855));
XNOR2X1 hap1_A_I1803 (.Y(N1859), .A(N1067), .B(N1830));
OR2XL hap1_A_I1804 (.Y(N1860), .A(N1067), .B(N1830));
ADDFX1 inst_cellmath__203_0_I923 (.CO(N1864), .S(N1863), .A(N1157), .B(N1859), .CI(N1277));
ADDFX1 inst_cellmath__203_0_I924 (.CO(N1866), .S(N1865), .A(N1187), .B(N1217), .CI(N1097));
ADDFX1 inst_cellmath__203_0_I925 (.CO(N1868), .S(N1867), .A(N1307), .B(N1127), .CI(N1247));
ADDFX1 inst_cellmath__203_0_I926 (.CO(N1870), .S(N1869), .A(N1832), .B(N1828), .CI(N1834));
ADDFX1 inst_cellmath__203_0_I927 (.CO(N1872), .S(N1871), .A(N1865), .B(N1863), .CI(N1867));
ADDFX1 inst_cellmath__203_0_I928 (.CO(N1874), .S(N1873), .A(N1838), .B(N1836), .CI(N1869));
ADDFX1 inst_cellmath__203_0_I929 (.CO(N1876), .S(N1875), .A(N1840), .B(N1871), .CI(N1873));
ADDFX1 inst_cellmath__203_0_I930 (.CO(N1878), .S(N1877), .A(N799), .B(N1842), .CI(N701));
ADDFX1 inst_cellmath__203_0_I931 (.CO(N1880), .S(N1879), .A(N673), .B(N645), .CI(N729));
ADDFX1 inst_cellmath__203_0_I932 (.CO(N1882), .S(N1881), .A(N757), .B(N1875), .CI(N1844));
ADDFX1 inst_cellmath__203_0_I933 (.CO(N1884), .S(N1883), .A(N1848), .B(N1846), .CI(N1877));
ADDFX1 inst_cellmath__203_0_I934 (.CO(N1886), .S(N1885), .A(N1850), .B(N1879), .CI(N1881));
ADDFX1 inst_cellmath__203_0_I935 (.CO(N1888), .S(N1887), .A(N1883), .B(N1852), .CI(N1854));
ADDFXL inst_cellmath__203_0_I936 (.CO(inst_cellmath__203_0_out1[26]), .S(inst_cellmath__203_0_out0[25]), .A(N1856), .B(N1885), .CI(N1887));
ADDHX1 inst_cellmath__203_0_I937 (.CO(N1892), .S(N1891), .A(N1860), .B(N1098));
ADDFX1 inst_cellmath__203_0_I938 (.CO(N1894), .S(N1893), .A(N1188), .B(N1891), .CI(N1218));
ADDFX1 inst_cellmath__203_0_I939 (.CO(N1896), .S(N1895), .A(N1278), .B(N1128), .CI(N1308));
ADDFX1 inst_cellmath__203_0_I940 (.CO(N1898), .S(N1897), .A(N1248), .B(N1158), .CI(N1864));
ADDFX1 inst_cellmath__203_0_I941 (.CO(N1900), .S(N1899), .A(N1868), .B(N1866), .CI(N1893));
ADDFX1 inst_cellmath__203_0_I942 (.CO(N1902), .S(N1901), .A(N1870), .B(N1895), .CI(N1897));
ADDFX1 inst_cellmath__203_0_I943 (.CO(N1904), .S(N1903), .A(N1899), .B(N1872), .CI(N1874));
ADDFX1 inst_cellmath__203_0_I944 (.CO(N1906), .S(N1905), .A(N5705), .B(N1901), .CI(N801));
ADDFX1 inst_cellmath__203_0_I945 (.CO(N1908), .S(N1907), .A(N1876), .B(N1903), .CI(N702));
ADDFX1 inst_cellmath__203_0_I946 (.CO(N1910), .S(N1909), .A(N730), .B(N674), .CI(N758));
ADDFX1 inst_cellmath__203_0_I947 (.CO(N1912), .S(N1911), .A(N1905), .B(N1878), .CI(N1880));
ADDFX1 inst_cellmath__203_0_I948 (.CO(N1914), .S(N1913), .A(N1882), .B(N1907), .CI(N1909));
ADDFX1 inst_cellmath__203_0_I949 (.CO(N1916), .S(N1915), .A(N1911), .B(N1884), .CI(N1886));
ADDFX1 inst_cellmath__203_0_I950 (.CO(inst_cellmath__203_0_out1[27]), .S(inst_cellmath__203_0_out0[26]), .A(N1888), .B(N1913), .CI(N1915));
XNOR2X1 hap1_A_I1805 (.Y(N1919), .A(N1099), .B(N1892));
OR2XL hap1_A_I1806 (.Y(N1920), .A(N1099), .B(N1892));
ADDFX1 inst_cellmath__203_0_I952 (.CO(N1924), .S(N1923), .A(N1189), .B(N1919), .CI(N1309));
ADDFX1 inst_cellmath__203_0_I953 (.CO(N1926), .S(N1925), .A(N1219), .B(N1249), .CI(N1129));
ADDFX1 inst_cellmath__203_0_I954 (.CO(N1928), .S(N1927), .A(N1279), .B(N1159), .CI(N1894));
ADDFX1 inst_cellmath__203_0_I955 (.CO(N1930), .S(N1929), .A(N1923), .B(N1896), .CI(N1925));
ADDFX1 inst_cellmath__203_0_I956 (.CO(N1932), .S(N1931), .A(N1900), .B(N1898), .CI(N1927));
ADDFX1 inst_cellmath__203_0_I957 (.CO(N1934), .S(N1933), .A(N1902), .B(N1929), .CI(N1931));
ADDFX1 inst_cellmath__203_0_I958 (.CO(N1936), .S(N1935), .A(N803), .B(N1904), .CI(N703));
ADDFX1 inst_cellmath__203_0_I959 (.CO(N1938), .S(N1937), .A(N675), .B(N1933), .CI(N731));
ADDFX1 inst_cellmath__203_0_I960 (.CO(N1940), .S(N1939), .A(N1906), .B(N759), .CI(N1908));
ADDFX1 inst_cellmath__203_0_I961 (.CO(N1942), .S(N1941), .A(N1910), .B(N1935), .CI(N1937));
ADDFX1 inst_cellmath__203_0_I962 (.CO(N1944), .S(N1943), .A(N1939), .B(N1912), .CI(N1914));
ADDFX1 inst_cellmath__203_0_I963 (.CO(inst_cellmath__203_0_out1[28]), .S(inst_cellmath__203_0_out0[27]), .A(N1916), .B(N1941), .CI(N1943));
INVXL fap1_A_I1807 (.Y(N5443), .A(N5820));
ADDFX1 fap1_A_I1808 (.CO(N1948), .S(N1947), .A(N1920), .B(N1130), .CI(N5443));
ADDFX1 inst_cellmath__203_0_I965 (.CO(N1952), .S(N1951), .A(N1250), .B(N1220), .CI(N1160));
ADDFX1 inst_cellmath__203_0_I966 (.CO(N1954), .S(N1953), .A(N1190), .B(N1310), .CI(N1280));
ADDFX1 inst_cellmath__203_0_I967 (.CO(N1956), .S(N1955), .A(N1924), .B(N1947), .CI(N1926));
ADDFX1 inst_cellmath__203_0_I968 (.CO(N1958), .S(N1957), .A(N1953), .B(N1951), .CI(N1928));
ADDFX1 inst_cellmath__203_0_I969 (.CO(N1960), .S(N1959), .A(N1930), .B(N1955), .CI(N1957));
ADDFX1 inst_cellmath__203_0_I970 (.CO(N1962), .S(N1961), .A(N5720), .B(N1932), .CI(N1959));
ADDFX1 inst_cellmath__203_0_I971 (.CO(N1964), .S(N1963), .A(N805), .B(N1934), .CI(N704));
ADDFX1 inst_cellmath__203_0_I972 (.CO(N1966), .S(N1965), .A(N760), .B(N732), .CI(N1961));
ADDFX1 inst_cellmath__203_0_I973 (.CO(N1968), .S(N1967), .A(N1938), .B(N1936), .CI(N1963));
ADDFX1 inst_cellmath__203_0_I974 (.CO(N1970), .S(N1969), .A(N1965), .B(N1940), .CI(N1942));
ADDFXL inst_cellmath__203_0_I975 (.CO(inst_cellmath__203_0_out1[29]), .S(inst_cellmath__203_0_out0[28]), .A(N1944), .B(N1967), .CI(N1969));
ADDFX1 inst_cellmath__203_0_I976 (.CO(N1974), .S(N1973), .A(N1131), .B(N5820), .CI(N1221));
ADDFX1 inst_cellmath__203_0_I977 (.CO(N1976), .S(N1975), .A(N1251), .B(N1281), .CI(N1161));
ADDFX1 inst_cellmath__203_0_I978 (.CO(N1978), .S(N1977), .A(N1311), .B(N1191), .CI(N1948));
ADDFX1 inst_cellmath__203_0_I979 (.CO(N1980), .S(N1979), .A(N1973), .B(N1952), .CI(N1954));
ADDFX1 inst_cellmath__203_0_I980 (.CO(N1982), .S(N1981), .A(N1977), .B(N1975), .CI(N1956));
ADDFX1 inst_cellmath__203_0_I981 (.CO(N1984), .S(N1983), .A(N1958), .B(N1979), .CI(N1981));
ADDFX1 inst_cellmath__203_0_I982 (.CO(N1986), .S(N1985), .A(N1983), .B(N1960), .CI(N807));
ADDFX1 inst_cellmath__203_0_I983 (.CO(N1988), .S(N1987), .A(N733), .B(N705), .CI(N1962));
ADDFXL inst_cellmath__203_0_I984 (.CO(N1990), .S(N1989), .A(N1964), .B(N761), .CI(N1985));
ADDFX1 inst_cellmath__203_0_I985 (.CO(N1992), .S(N1991), .A(N1987), .B(N1966), .CI(N1968));
ADDFX1 inst_cellmath__203_0_I986 (.CO(inst_cellmath__203_0_out1[30]), .S(inst_cellmath__203_0_out0[29]), .A(N1970), .B(N1989), .CI(N1991));
INVXL fap1_A_I1809 (.Y(N5452), .A(N5848));
ADDFX1 fap1_A_I1810 (.CO(N1996), .S(N1995), .A(N1252), .B(N1162), .CI(N5452));
ADDFX1 inst_cellmath__203_0_I988 (.CO(N2000), .S(N1999), .A(N1192), .B(N1282), .CI(N1222));
ADDFX1 inst_cellmath__203_0_I989 (.CO(N2002), .S(N2001), .A(N1974), .B(N1312), .CI(N1976));
ADDFX1 inst_cellmath__203_0_I990 (.CO(N2004), .S(N2003), .A(N1995), .B(N1978), .CI(N1999));
ADDFX1 inst_cellmath__203_0_I991 (.CO(N2006), .S(N2005), .A(N2001), .B(N1980), .CI(N1982));
ADDFX1 inst_cellmath__203_0_I992 (.CO(N2008), .S(N2007), .A(N2005), .B(N2003), .CI(N5736));
ADDFX1 inst_cellmath__203_0_I993 (.CO(N2010), .S(N2009), .A(N809), .B(N1984), .CI(N734));
ADDFX1 inst_cellmath__203_0_I994 (.CO(N2012), .S(N2011), .A(N2007), .B(N762), .CI(N1986));
ADDFXL inst_cellmath__203_0_I995 (.CO(N2014), .S(N2013), .A(N2009), .B(N1988), .CI(N1990));
ADDFXL inst_cellmath__203_0_I996 (.CO(inst_cellmath__203_0_out1[31]), .S(inst_cellmath__203_0_out0[30]), .A(N1992), .B(N2011), .CI(N2013));
ADDFX1 inst_cellmath__203_0_I997 (.CO(N2018), .S(N2017), .A(N1163), .B(N5848), .CI(N1253));
ADDFX1 inst_cellmath__203_0_I998 (.CO(N2020), .S(N2019), .A(N1283), .B(N1313), .CI(N1193));
ADDFX1 inst_cellmath__203_0_I999 (.CO(N2022), .S(N2021), .A(N1996), .B(N1223), .CI(N2000));
ADDFX1 inst_cellmath__203_0_I1000 (.CO(N2024), .S(N2023), .A(N2019), .B(N2017), .CI(N2002));
ADDFX1 inst_cellmath__203_0_I1001 (.CO(N2026), .S(N2025), .A(N2021), .B(N2004), .CI(N2023));
ADDFX1 inst_cellmath__203_0_I1002 (.CO(N2028), .S(N2027), .A(N2025), .B(N2006), .CI(N811));
ADDFX1 inst_cellmath__203_0_I1003 (.CO(N2030), .S(N2029), .A(N735), .B(N2008), .CI(N763));
ADDFX1 inst_cellmath__203_0_I1004 (.CO(N2032), .S(N2031), .A(N2010), .B(N2027), .CI(N2012));
ADDFX1 inst_cellmath__203_0_I1005 (.CO(inst_cellmath__203_0_out1[32]), .S(inst_cellmath__203_0_out0[31]), .A(N2014), .B(N2029), .CI(N2031));
INVXL fap1_A_I1811 (.Y(N5461), .A(N5874));
ADDFX1 fap1_A_I1812 (.CO(N2036), .S(N2035), .A(N1284), .B(N1194), .CI(N5461));
ADDFX1 inst_cellmath__203_0_I1007 (.CO(N2040), .S(N2039), .A(N1224), .B(N1314), .CI(N1254));
ADDFX1 inst_cellmath__203_0_I1008 (.CO(N2042), .S(N2041), .A(N2020), .B(N2018), .CI(N2035));
ADDFX1 inst_cellmath__203_0_I1009 (.CO(N2044), .S(N2043), .A(N2022), .B(N2039), .CI(N2024));
ADDFX1 inst_cellmath__203_0_I1010 (.CO(N2046), .S(N2045), .A(N2026), .B(N2041), .CI(N2043));
ADDFX1 inst_cellmath__203_0_I1011 (.CO(N2048), .S(N2047), .A(N813), .B(N5751), .CI(N764));
ADDFX1 inst_cellmath__203_0_I1012 (.CO(N2050), .S(N2049), .A(N2028), .B(N2045), .CI(N2030));
ADDFX1 inst_cellmath__203_0_I1013 (.CO(inst_cellmath__203_0_out1[33]), .S(inst_cellmath__203_0_out0[32]), .A(N2032), .B(N2047), .CI(N2049));
ADDFX1 inst_cellmath__203_0_I1014 (.CO(N2054), .S(N2053), .A(N1195), .B(N5874), .CI(N1285));
ADDFX1 inst_cellmath__203_0_I1015 (.CO(N2056), .S(N2055), .A(N1225), .B(N1315), .CI(N1255));
ADDFX1 inst_cellmath__203_0_I1016 (.CO(N2058), .S(N2057), .A(N2040), .B(N2036), .CI(N2053));
ADDFX1 inst_cellmath__203_0_I1017 (.CO(N2060), .S(N2059), .A(N2042), .B(N2055), .CI(N2057));
ADDFX1 inst_cellmath__203_0_I1018 (.CO(N2062), .S(N2061), .A(N2059), .B(N2044), .CI(N815));
ADDFX1 inst_cellmath__203_0_I1019 (.CO(N2064), .S(N2063), .A(N765), .B(N2046), .CI(N2061));
ADDFX1 inst_cellmath__203_0_I1020 (.CO(inst_cellmath__203_0_out0[34]), .S(inst_cellmath__203_0_out0[33]), .A(N2050), .B(N2048), .CI(N2063));
INVXL fap1_A_I1813 (.Y(N5470), .A(N5900));
ADDFX1 fap1_A_I1814 (.CO(N2068), .S(N2067), .A(N1316), .B(N1226), .CI(N5470));
ADDFX1 inst_cellmath__203_0_I1022 (.CO(N2072), .S(N2071), .A(N1286), .B(N1256), .CI(N2054));
ADDFX1 inst_cellmath__203_0_I1023 (.CO(N2074), .S(N2073), .A(N2067), .B(N2056), .CI(N2071));
ADDFX1 inst_cellmath__203_0_I1024 (.CO(N2076), .S(N2075), .A(N2073), .B(N2058), .CI(N2060));
ADDFX1 inst_cellmath__203_0_I1025 (.CO(N2078), .S(N2077), .A(N2075), .B(N817), .CI(N5767));
ADDFX1 inst_cellmath__203_0_I1026 (.CO(inst_cellmath__203_0_out0[35]), .S(inst_cellmath__203_0_out1[34]), .A(N2077), .B(N2062), .CI(N2064));
ADDFX1 inst_cellmath__203_0_I1027 (.CO(N2082), .S(N2081), .A(N1227), .B(N5900), .CI(N1317));
ADDFX1 inst_cellmath__203_0_I1028 (.CO(N2084), .S(N2083), .A(N1287), .B(N1257), .CI(N2068));
ADDFX1 inst_cellmath__203_0_I1029 (.CO(N2086), .S(N2085), .A(N2072), .B(N2081), .CI(N2083));
ADDFX1 inst_cellmath__203_0_I1030 (.CO(N2088), .S(N2087), .A(N2085), .B(N2074), .CI(N2076));
ADDFX1 inst_cellmath__203_0_I1031 (.CO(inst_cellmath__203_0_out0[36]), .S(inst_cellmath__203_0_out1[35]), .A(N2087), .B(N819), .CI(N2078));
INVXL fap1_A_I1815 (.Y(N5479), .A(N5926));
ADDFX1 fap1_A_I1816 (.CO(N2092), .S(N2091), .A(N1288), .B(N1258), .CI(N5479));
ADDFX1 inst_cellmath__203_0_I1033 (.CO(N2096), .S(N2095), .A(N2082), .B(N1318), .CI(N2091));
ADDFX1 inst_cellmath__203_0_I1034 (.CO(N2098), .S(N2097), .A(N2095), .B(N2084), .CI(N2086));
ADDFX1 inst_cellmath__203_0_I1035 (.CO(inst_cellmath__203_0_out0[37]), .S(inst_cellmath__203_0_out1[36]), .A(N1366), .B(N2097), .CI(N2088));
ADDFX1 inst_cellmath__203_0_I1036 (.CO(N2102), .S(N2101), .A(N1259), .B(N5926), .CI(N1289));
ADDFX1 inst_cellmath__203_0_I1037 (.CO(N2104), .S(N2103), .A(N2092), .B(N1319), .CI(N2101));
ADDFX1 inst_cellmath__203_0_I1038 (.CO(inst_cellmath__203_0_out0[38]), .S(inst_cellmath__203_0_out1[37]), .A(N2103), .B(N2096), .CI(N2098));
ADDFX1 inst_cellmath__203_0_I1039 (.CO(N2108), .S(N2107), .A(N1290), .B(N5949), .CI(N1320));
ADDFX1 inst_cellmath__203_0_I1040 (.CO(inst_cellmath__203_0_out0[39]), .S(inst_cellmath__203_0_out1[38]), .A(N2107), .B(N2102), .CI(N2104));
INVXL inst_cellmath__203_0_I1041 (.Y(N2111), .A(N2112));
ADDFX1 inst_cellmath__203_0_I1042 (.CO(inst_cellmath__203_0_out0[40]), .S(inst_cellmath__203_0_out1[39]), .A(N1321), .B(N2111), .CI(N2108));
ADDFX1 inst_cellmath__203_0_I1043 (.CO(inst_cellmath__203_0_out0[41]), .S(inst_cellmath__203_0_out1[40]), .A(N2112), .B(N5974), .CI(N1322));
INVXL inst_cellmath__203_0_I1044 (.Y(inst_cellmath__203_0_out1[41]), .A(inst_cellmath__203_0_out0[42]));
assign inst_cellmath__203_0_out0[0] = 1'B0;
assign inst_cellmath__203_0_out0[43] = 1'B0;
assign inst_cellmath__203_0_out0[44] = 1'B0;
assign inst_cellmath__203_0_out0[45] = 1'B0;
assign inst_cellmath__203_0_out0[46] = 1'B0;
assign inst_cellmath__203_0_out1[43] = 1'B1;
assign inst_cellmath__203_0_out1[44] = 1'B1;
assign inst_cellmath__203_0_out1[45] = 1'B1;
assign inst_cellmath__203_0_out1[46] = 1'B1;
endmodule

module cynw_cm_float_cos_inst_cellmath__201_0_bdw1157874770_bdw (
	inst_cellmath__201_0_out0,
	inst_cellmath__201_0_in0,
	inst_cellmath__201_0_in1,
	inst_cellmath__201_0_in2
	); /* architecture "gate_level" */ 
output [49:0] inst_cellmath__201_0_out0;
input [46:0] inst_cellmath__201_0_in0,
	inst_cellmath__201_0_in1;
input [72:43] inst_cellmath__201_0_in2;
wire [46:0] inst_cellmath__203__W1;
wire N989,N991,N992,N993,N994,N995,N996 
	,N997,N998,N999,N1000,N1001,N1002,N1003,N1004 
	,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012 
	,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020 
	,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028 
	,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036 
	,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044 
	,N1045,N1046,N1047,N1048,N1049,N1054,N1055,N1056 
	,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064 
	,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072 
	,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080 
	,N1081,N1082,N1083,N1084,N1085,N1088,N1089,N1096 
	,N1104,N1116,N1136,N1138,N1156,N1174,N1196,N1226 
	,N1228,N1256,N1292,N1294,N1298,N1299,N1330,N1339 
	,N1342,N1345,N1348,N1351,N1354,N1357,N1360,N1363 
	,N1366,N1369,N1372,N1375,N1378,N1381,N1384,N1403 
	,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412 
	,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420 
	,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428 
	,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436 
	,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444 
	,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452 
	,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460 
	,N1461,N1462,N1463,N1464,N1465,N1466,N1470,N1472 
	,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480 
	,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488 
	,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496 
	,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504 
	,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512 
	,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520 
	,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528 
	,N1529,N1530,N1531,N1534,N1539,N1541,N1543,N1544 
	,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552 
	,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560 
	,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568 
	,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576 
	,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584 
	,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592 
	,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600 
	,N1609,N1611,N1613,N1615,N1617,N1618,N1619,N1620 
	,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628 
	,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636 
	,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644 
	,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652 
	,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660 
	,N1661,N1662,N1663,N1664,N1665,N1666,N1683,N1685 
	,N1687,N1689,N1691,N1693,N1695,N1697,N1699,N1700 
	,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708 
	,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716 
	,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724 
	,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732 
	,N1765,N1767,N1769,N1771,N1773,N1775,N1777,N1779 
	,N1781,N1783,N1785,N1787,N1789,N1791,N1793,N1797 
	,N1798,N1870,N1873,N1876,N1879,N1882,N1885,N1888 
	,N1891,N1894,N1897,N1900,N1903,N1906,N1909,N1912 
	,N1915,N1918,N1921,N1924,N1927,N1930,N1933,N1936 
	,N1939,N1942,N1945,N1948,N1951,N1954,N1957,N1960 
	,N2310,N2315,N2316,N2325,N2332,N2333,N2349,N2350 
	,N2364,N2376,N2377,N2396,N2397,N2399,N2413,N2414 
	,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428 
	,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2438 
	,N2456,N2483;
INVXL inst_cellmath__201_0_I102 (.Y(inst_cellmath__203__W1[46]), .A(inst_cellmath__201_0_in0[46]));
INVXL inst_cellmath__201_0_I243 (.Y(N989), .A(inst_cellmath__201_0_in1[46]));
ADDHX1 inst_cellmath__201_0_I245 (.CO(N992), .S(N991), .A(inst_cellmath__201_0_in2[43]), .B(inst_cellmath__201_0_in1[18]));
ADDFX1 inst_cellmath__201_0_I246 (.CO(N994), .S(N993), .A(inst_cellmath__201_0_in1[19]), .B(inst_cellmath__201_0_in2[44]), .CI(inst_cellmath__201_0_in0[19]));
ADDFHX1 inst_cellmath__201_0_I247 (.CO(N996), .S(N995), .A(inst_cellmath__201_0_in1[20]), .B(inst_cellmath__201_0_in2[45]), .CI(inst_cellmath__201_0_in0[20]));
ADDFX1 inst_cellmath__201_0_I248 (.CO(N998), .S(N997), .A(inst_cellmath__201_0_in1[21]), .B(inst_cellmath__201_0_in2[46]), .CI(inst_cellmath__201_0_in0[21]));
ADDFHX1 inst_cellmath__201_0_I249 (.CO(N1000), .S(N999), .A(inst_cellmath__201_0_in1[22]), .B(inst_cellmath__201_0_in2[47]), .CI(inst_cellmath__201_0_in0[22]));
ADDFHX1 inst_cellmath__201_0_I250 (.CO(N1002), .S(N1001), .A(inst_cellmath__201_0_in1[23]), .B(inst_cellmath__201_0_in2[48]), .CI(inst_cellmath__201_0_in0[23]));
ADDFHX1 inst_cellmath__201_0_I251 (.CO(N1004), .S(N1003), .A(inst_cellmath__201_0_in1[24]), .B(inst_cellmath__201_0_in2[49]), .CI(inst_cellmath__201_0_in0[24]));
ADDFX1 inst_cellmath__201_0_I252 (.CO(N1006), .S(N1005), .A(inst_cellmath__201_0_in1[25]), .B(inst_cellmath__201_0_in2[50]), .CI(inst_cellmath__201_0_in0[25]));
ADDFX1 inst_cellmath__201_0_I253 (.CO(N1008), .S(N1007), .A(inst_cellmath__201_0_in1[26]), .B(inst_cellmath__201_0_in2[51]), .CI(inst_cellmath__201_0_in0[26]));
ADDFX1 inst_cellmath__201_0_I254 (.CO(N1010), .S(N1009), .A(inst_cellmath__201_0_in1[27]), .B(inst_cellmath__201_0_in2[52]), .CI(inst_cellmath__201_0_in0[27]));
ADDFX1 inst_cellmath__201_0_I255 (.CO(N1012), .S(N1011), .A(inst_cellmath__201_0_in1[28]), .B(inst_cellmath__201_0_in2[53]), .CI(inst_cellmath__201_0_in0[28]));
ADDFX1 inst_cellmath__201_0_I256 (.CO(N1014), .S(N1013), .A(inst_cellmath__201_0_in1[29]), .B(inst_cellmath__201_0_in2[54]), .CI(inst_cellmath__201_0_in0[29]));
ADDFX1 inst_cellmath__201_0_I257 (.CO(N1016), .S(N1015), .A(inst_cellmath__201_0_in1[30]), .B(inst_cellmath__201_0_in2[55]), .CI(inst_cellmath__201_0_in0[30]));
ADDFX1 inst_cellmath__201_0_I258 (.CO(N1018), .S(N1017), .A(inst_cellmath__201_0_in1[31]), .B(inst_cellmath__201_0_in2[56]), .CI(inst_cellmath__201_0_in0[31]));
ADDFX1 inst_cellmath__201_0_I259 (.CO(N1020), .S(N1019), .A(inst_cellmath__201_0_in1[32]), .B(inst_cellmath__201_0_in2[57]), .CI(inst_cellmath__201_0_in0[32]));
ADDFX1 inst_cellmath__201_0_I260 (.CO(N1022), .S(N1021), .A(inst_cellmath__201_0_in0[33]), .B(inst_cellmath__201_0_in2[58]), .CI(inst_cellmath__201_0_in1[33]));
ADDFX1 inst_cellmath__201_0_I261 (.CO(N1024), .S(N1023), .A(inst_cellmath__201_0_in1[34]), .B(inst_cellmath__201_0_in2[59]), .CI(inst_cellmath__201_0_in0[34]));
ADDFX1 inst_cellmath__201_0_I262 (.CO(N1026), .S(N1025), .A(inst_cellmath__201_0_in0[35]), .B(inst_cellmath__201_0_in2[60]), .CI(inst_cellmath__201_0_in1[35]));
ADDFX1 inst_cellmath__201_0_I263 (.CO(N1028), .S(N1027), .A(inst_cellmath__201_0_in1[36]), .B(inst_cellmath__201_0_in2[61]), .CI(inst_cellmath__201_0_in0[36]));
ADDFX1 inst_cellmath__201_0_I264 (.CO(N1030), .S(N1029), .A(inst_cellmath__201_0_in1[37]), .B(inst_cellmath__201_0_in2[62]), .CI(inst_cellmath__201_0_in0[37]));
ADDFX1 inst_cellmath__201_0_I265 (.CO(N1032), .S(N1031), .A(inst_cellmath__201_0_in1[38]), .B(inst_cellmath__201_0_in2[63]), .CI(inst_cellmath__201_0_in0[38]));
ADDFX1 inst_cellmath__201_0_I266 (.CO(N1034), .S(N1033), .A(inst_cellmath__201_0_in1[39]), .B(inst_cellmath__201_0_in2[64]), .CI(inst_cellmath__201_0_in0[39]));
ADDFX1 inst_cellmath__201_0_I267 (.CO(N1036), .S(N1035), .A(inst_cellmath__201_0_in1[40]), .B(inst_cellmath__201_0_in2[65]), .CI(inst_cellmath__201_0_in0[40]));
ADDFX1 inst_cellmath__201_0_I268 (.CO(N1038), .S(N1037), .A(inst_cellmath__201_0_in2[66]), .B(inst_cellmath__201_0_in1[41]), .CI(inst_cellmath__201_0_in0[41]));
ADDFX1 inst_cellmath__201_0_I269 (.CO(N1040), .S(N1039), .A(inst_cellmath__201_0_in0[42]), .B(inst_cellmath__201_0_in1[42]), .CI(inst_cellmath__201_0_in2[67]));
ADDFX1 inst_cellmath__201_0_I270 (.CO(N1042), .S(N1041), .A(inst_cellmath__201_0_in0[43]), .B(inst_cellmath__201_0_in1[43]), .CI(inst_cellmath__201_0_in2[68]));
ADDFX1 inst_cellmath__201_0_I271 (.CO(N1044), .S(N1043), .A(inst_cellmath__201_0_in0[44]), .B(inst_cellmath__201_0_in1[44]), .CI(inst_cellmath__201_0_in2[69]));
ADDFX1 inst_cellmath__201_0_I272 (.CO(N1046), .S(N1045), .A(inst_cellmath__201_0_in0[45]), .B(inst_cellmath__201_0_in1[45]), .CI(inst_cellmath__201_0_in2[70]));
ADDFX1 inst_cellmath__201_0_I273 (.CO(N1048), .S(N1047), .A(inst_cellmath__203__W1[46]), .B(N989), .CI(inst_cellmath__201_0_in2[71]));
INVXL inst_cellmath__201_0_I274 (.Y(N1049), .A(inst_cellmath__201_0_in2[72]));
NOR2XL inst_cellmath__201_0_I276 (.Y(N1054), .A(inst_cellmath__201_0_in1[1]), .B(inst_cellmath__201_0_in0[1]));
NAND2XL inst_cellmath__201_0_I277 (.Y(N1055), .A(inst_cellmath__201_0_in1[1]), .B(inst_cellmath__201_0_in0[1]));
NOR2XL inst_cellmath__201_0_I278 (.Y(N1056), .A(inst_cellmath__201_0_in1[2]), .B(inst_cellmath__201_0_in0[2]));
NAND2XL inst_cellmath__201_0_I279 (.Y(N1057), .A(inst_cellmath__201_0_in1[2]), .B(inst_cellmath__201_0_in0[2]));
NOR2XL inst_cellmath__201_0_I280 (.Y(N1058), .A(inst_cellmath__201_0_in1[3]), .B(inst_cellmath__201_0_in0[3]));
NAND2XL inst_cellmath__201_0_I281 (.Y(N1059), .A(inst_cellmath__201_0_in1[3]), .B(inst_cellmath__201_0_in0[3]));
NOR2XL inst_cellmath__201_0_I282 (.Y(N1060), .A(inst_cellmath__201_0_in1[4]), .B(inst_cellmath__201_0_in0[4]));
NAND2XL inst_cellmath__201_0_I283 (.Y(N1061), .A(inst_cellmath__201_0_in1[4]), .B(inst_cellmath__201_0_in0[4]));
NOR2XL inst_cellmath__201_0_I284 (.Y(N1062), .A(inst_cellmath__201_0_in1[5]), .B(inst_cellmath__201_0_in0[5]));
NAND2XL inst_cellmath__201_0_I285 (.Y(N1063), .A(inst_cellmath__201_0_in1[5]), .B(inst_cellmath__201_0_in0[5]));
NOR2XL inst_cellmath__201_0_I286 (.Y(N1064), .A(inst_cellmath__201_0_in1[6]), .B(inst_cellmath__201_0_in0[6]));
NAND2XL inst_cellmath__201_0_I287 (.Y(N1065), .A(inst_cellmath__201_0_in1[6]), .B(inst_cellmath__201_0_in0[6]));
NOR2XL inst_cellmath__201_0_I288 (.Y(N1066), .A(inst_cellmath__201_0_in1[7]), .B(inst_cellmath__201_0_in0[7]));
NAND2XL inst_cellmath__201_0_I289 (.Y(N1067), .A(inst_cellmath__201_0_in1[7]), .B(inst_cellmath__201_0_in0[7]));
NOR2XL inst_cellmath__201_0_I290 (.Y(N1068), .A(inst_cellmath__201_0_in1[8]), .B(inst_cellmath__201_0_in0[8]));
NAND2XL inst_cellmath__201_0_I291 (.Y(N1069), .A(inst_cellmath__201_0_in1[8]), .B(inst_cellmath__201_0_in0[8]));
NOR2XL inst_cellmath__201_0_I292 (.Y(N1070), .A(inst_cellmath__201_0_in1[9]), .B(inst_cellmath__201_0_in0[9]));
NAND2XL inst_cellmath__201_0_I293 (.Y(N1071), .A(inst_cellmath__201_0_in1[9]), .B(inst_cellmath__201_0_in0[9]));
NOR2XL inst_cellmath__201_0_I294 (.Y(N1072), .A(inst_cellmath__201_0_in1[10]), .B(inst_cellmath__201_0_in0[10]));
NAND2XL inst_cellmath__201_0_I295 (.Y(N1073), .A(inst_cellmath__201_0_in1[10]), .B(inst_cellmath__201_0_in0[10]));
NOR2XL inst_cellmath__201_0_I296 (.Y(N1074), .A(inst_cellmath__201_0_in1[11]), .B(inst_cellmath__201_0_in0[11]));
NAND2XL inst_cellmath__201_0_I297 (.Y(N1075), .A(inst_cellmath__201_0_in1[11]), .B(inst_cellmath__201_0_in0[11]));
NOR2XL inst_cellmath__201_0_I298 (.Y(N1076), .A(inst_cellmath__201_0_in1[12]), .B(inst_cellmath__201_0_in0[12]));
NAND2XL inst_cellmath__201_0_I299 (.Y(N1077), .A(inst_cellmath__201_0_in1[12]), .B(inst_cellmath__201_0_in0[12]));
NOR2XL inst_cellmath__201_0_I300 (.Y(N1078), .A(inst_cellmath__201_0_in1[13]), .B(inst_cellmath__201_0_in0[13]));
NAND2XL inst_cellmath__201_0_I301 (.Y(N1079), .A(inst_cellmath__201_0_in1[13]), .B(inst_cellmath__201_0_in0[13]));
NOR2XL inst_cellmath__201_0_I302 (.Y(N1080), .A(inst_cellmath__201_0_in1[14]), .B(inst_cellmath__201_0_in0[14]));
NAND2XL inst_cellmath__201_0_I303 (.Y(N1081), .A(inst_cellmath__201_0_in1[14]), .B(inst_cellmath__201_0_in0[14]));
NOR2XL inst_cellmath__201_0_I304 (.Y(N1082), .A(inst_cellmath__201_0_in1[15]), .B(inst_cellmath__201_0_in0[15]));
NAND2XL inst_cellmath__201_0_I305 (.Y(N1083), .A(inst_cellmath__201_0_in1[15]), .B(inst_cellmath__201_0_in0[15]));
NOR2XL inst_cellmath__201_0_I306 (.Y(N1084), .A(inst_cellmath__201_0_in1[16]), .B(inst_cellmath__201_0_in0[16]));
NAND2XL inst_cellmath__201_0_I307 (.Y(N1085), .A(inst_cellmath__201_0_in1[16]), .B(inst_cellmath__201_0_in0[16]));
AOI21XL inst_cellmath__201_0_I310 (.Y(N1088), .A0(N1057), .A1(N1054), .B0(N1056));
NAND2XL inst_cellmath__201_0_I311 (.Y(N1089), .A(N1057), .B(N1055));
AND2XL inst_cellmath__201_0_I1498 (.Y(N2310), .A(inst_cellmath__201_0_in0[0]), .B(inst_cellmath__201_0_in1[0]));
OAI21XL inst_cellmath__201_0_I318 (.Y(N1096), .A0(N1089), .A1(N2310), .B0(N1088));
AOI21XL inst_cellmath__201_0_I326 (.Y(N1104), .A0(N1059), .A1(N1096), .B0(N1058));
INVXL inst_cellmath__201_0_I1349 (.Y(N2315), .A(N1060));
INVXL inst_cellmath__201_0_I1350 (.Y(N2316), .A(N1061));
OAI21XL inst_cellmath__201_0_I338 (.Y(N1116), .A0(N2316), .A1(N1104), .B0(N2315));
AO21XL inst_cellmath__201_0_I1499 (.Y(N2325), .A0(N1062), .A1(N1065), .B0(N1064));
AOI21XL inst_cellmath__201_0_I358 (.Y(N1136), .A0(N1063), .A1(N1116), .B0(N1062));
AOI31X1 inst_cellmath__201_0_I1501 (.Y(N1138), .A0(N1065), .A1(N1063), .A2(N1116), .B0(N2325));
INVXL inst_cellmath__201_0_I1366 (.Y(N2332), .A(N1066));
INVXL inst_cellmath__201_0_I1367 (.Y(N2333), .A(N1067));
OAI21X1 inst_cellmath__201_0_I378 (.Y(N1156), .A0(N2333), .A1(N1138), .B0(N2332));
AOI21X1 inst_cellmath__201_0_I396 (.Y(N1174), .A0(N1069), .A1(N1156), .B0(N1068));
INVXL inst_cellmath__201_0_I1383 (.Y(N2349), .A(N1070));
INVXL inst_cellmath__201_0_I1384 (.Y(N2350), .A(N1071));
OAI21X1 inst_cellmath__201_0_I418 (.Y(N1196), .A0(N2350), .A1(N1174), .B0(N2349));
AO21XL inst_cellmath__201_0_I1502 (.Y(N2364), .A0(N1072), .A1(N1075), .B0(N1074));
AOI21XL inst_cellmath__201_0_I448 (.Y(N1226), .A0(N1073), .A1(N1196), .B0(N1072));
AOI31X2 inst_cellmath__201_0_I1544 (.Y(N1228), .A0(N1075), .A1(N1073), .A2(N1196), .B0(N2364));
INVXL inst_cellmath__201_0_I1410 (.Y(N2376), .A(N1076));
INVXL inst_cellmath__201_0_I1411 (.Y(N2377), .A(N1077));
OAI21X2 inst_cellmath__201_0_I478 (.Y(N1256), .A0(N2377), .A1(N1228), .B0(N2376));
AO21XL inst_cellmath__201_0_I1505 (.Y(N2396), .A0(N1078), .A1(N1081), .B0(N1080));
AND2XL inst_cellmath__201_0_I1506 (.Y(N2397), .A(N1081), .B(N1079));
NOR2BX1 andori2bb1_A_I2723 (.Y(N2483), .AN(N1055), .B(N2310));
NOR2XL andori2bb1_A_I1639 (.Y(N2399), .A(N2483), .B(N1054));
AOI21XL inst_cellmath__201_0_I514 (.Y(N1292), .A0(N1079), .A1(N1256), .B0(N1078));
AOI21X2 inst_cellmath__201_0_I516 (.Y(N1294), .A0(N2397), .A1(N1256), .B0(N2396));
INVXL inst_cellmath__201_0_I1447 (.Y(N2413), .A(N1082));
INVXL inst_cellmath__201_0_I1448 (.Y(N2414), .A(N1083));
AOI21XL inst_cellmath__201_0_I520 (.Y(N1298), .A0(N1085), .A1(N1082), .B0(N1084));
NAND2XL inst_cellmath__201_0_I521 (.Y(N1299), .A(N1085), .B(N1083));
OAI21XL inst_cellmath__201_0_I552 (.Y(N1330), .A0(N2414), .A1(N1294), .B0(N2413));
OAI21X2 inst_cellmath__201_0_I554 (.Y(N1403), .A0(N1299), .A1(N1294), .B0(N1298));
NAND2BXL inst_cellmath__201_0_I561 (.Y(N1339), .AN(N1054), .B(N1055));
NAND2BXL inst_cellmath__201_0_I564 (.Y(N1342), .AN(N1056), .B(N1057));
NAND2BXL inst_cellmath__201_0_I567 (.Y(N1345), .AN(N1058), .B(N1059));
NAND2BXL inst_cellmath__201_0_I570 (.Y(N1348), .AN(N1060), .B(N1061));
NAND2BXL inst_cellmath__201_0_I573 (.Y(N1351), .AN(N1062), .B(N1063));
NAND2BXL inst_cellmath__201_0_I576 (.Y(N1354), .AN(N1064), .B(N1065));
NAND2BXL inst_cellmath__201_0_I579 (.Y(N1357), .AN(N1066), .B(N1067));
NAND2BXL inst_cellmath__201_0_I582 (.Y(N1360), .AN(N1068), .B(N1069));
NAND2BXL inst_cellmath__201_0_I585 (.Y(N1363), .AN(N1070), .B(N1071));
NAND2BXL inst_cellmath__201_0_I588 (.Y(N1366), .AN(N1072), .B(N1073));
NAND2BXL inst_cellmath__201_0_I591 (.Y(N1369), .AN(N1074), .B(N1075));
NAND2BXL inst_cellmath__201_0_I594 (.Y(N1372), .AN(N1076), .B(N1077));
NAND2BXL inst_cellmath__201_0_I597 (.Y(N1375), .AN(N1078), .B(N1079));
NAND2BXL inst_cellmath__201_0_I600 (.Y(N1378), .AN(N1080), .B(N1081));
NAND2BXL inst_cellmath__201_0_I603 (.Y(N1381), .AN(N1082), .B(N1083));
NAND2BXL inst_cellmath__201_0_I606 (.Y(N1384), .AN(N1084), .B(N1085));
XOR2XL inst_cellmath__201_0_I607 (.Y(inst_cellmath__201_0_out0[0]), .A(inst_cellmath__201_0_in0[0]), .B(inst_cellmath__201_0_in1[0]));
XNOR2X1 inst_cellmath__201_0_I608 (.Y(inst_cellmath__201_0_out0[1]), .A(N2310), .B(N1339));
XNOR2X1 inst_cellmath__201_0_I609 (.Y(inst_cellmath__201_0_out0[2]), .A(N2399), .B(N1342));
XOR2XL inst_cellmath__201_0_I1509 (.Y(inst_cellmath__201_0_out0[3]), .A(N1096), .B(N1345));
XNOR2X1 inst_cellmath__201_0_I611 (.Y(inst_cellmath__201_0_out0[4]), .A(N1104), .B(N1348));
XOR2XL inst_cellmath__201_0_I1510 (.Y(inst_cellmath__201_0_out0[5]), .A(N1116), .B(N1351));
XNOR2X1 inst_cellmath__201_0_I613 (.Y(inst_cellmath__201_0_out0[6]), .A(N1136), .B(N1354));
XNOR2X1 inst_cellmath__201_0_I614 (.Y(inst_cellmath__201_0_out0[7]), .A(N1138), .B(N1357));
XOR2XL inst_cellmath__201_0_I1511 (.Y(inst_cellmath__201_0_out0[8]), .A(N1156), .B(N1360));
XNOR2X1 inst_cellmath__201_0_I616 (.Y(inst_cellmath__201_0_out0[9]), .A(N1174), .B(N1363));
XOR2XL inst_cellmath__201_0_I1512 (.Y(inst_cellmath__201_0_out0[10]), .A(N1196), .B(N1366));
XNOR2X1 inst_cellmath__201_0_I618 (.Y(inst_cellmath__201_0_out0[11]), .A(N1226), .B(N1369));
XNOR2X1 inst_cellmath__201_0_I619 (.Y(inst_cellmath__201_0_out0[12]), .A(N1228), .B(N1372));
XOR2XL inst_cellmath__201_0_I1513 (.Y(inst_cellmath__201_0_out0[13]), .A(N1256), .B(N1375));
XNOR2X1 inst_cellmath__201_0_I621 (.Y(inst_cellmath__201_0_out0[14]), .A(N1292), .B(N1378));
XNOR2X1 inst_cellmath__201_0_I622 (.Y(inst_cellmath__201_0_out0[15]), .A(N1294), .B(N1381));
XOR2XL inst_cellmath__201_0_I623 (.Y(inst_cellmath__201_0_out0[16]), .A(N1330), .B(N1384));
NOR2XL inst_cellmath__201_0_I626 (.Y(N1405), .A(inst_cellmath__201_0_in1[17]), .B(inst_cellmath__201_0_in0[17]));
NAND2XL inst_cellmath__201_0_I627 (.Y(N1406), .A(inst_cellmath__201_0_in1[17]), .B(inst_cellmath__201_0_in0[17]));
NOR2XL inst_cellmath__201_0_I628 (.Y(N1407), .A(N991), .B(inst_cellmath__201_0_in0[18]));
NAND2XL inst_cellmath__201_0_I629 (.Y(N1408), .A(N991), .B(inst_cellmath__201_0_in0[18]));
NOR2X2 inst_cellmath__201_0_I630 (.Y(N1409), .A(N992), .B(N993));
NAND2X2 inst_cellmath__201_0_I631 (.Y(N1410), .A(N992), .B(N993));
NOR2X4 inst_cellmath__201_0_I632 (.Y(N1411), .A(N994), .B(N995));
NAND2X6 inst_cellmath__201_0_I633 (.Y(N1412), .A(N994), .B(N995));
NOR2X4 inst_cellmath__201_0_I634 (.Y(N1413), .A(N996), .B(N997));
NAND2X4 inst_cellmath__201_0_I635 (.Y(N1414), .A(N996), .B(N997));
NOR2X4 inst_cellmath__201_0_I636 (.Y(N1415), .A(N998), .B(N999));
NAND2X4 inst_cellmath__201_0_I637 (.Y(N1416), .A(N998), .B(N999));
NOR2X2 inst_cellmath__201_0_I638 (.Y(N1417), .A(N1000), .B(N1001));
NAND2X4 inst_cellmath__201_0_I639 (.Y(N1418), .A(N1000), .B(N1001));
NOR2X2 inst_cellmath__201_0_I640 (.Y(N1419), .A(N1002), .B(N1003));
NAND2X4 inst_cellmath__201_0_I641 (.Y(N1420), .A(N1002), .B(N1003));
NOR2X2 inst_cellmath__201_0_I642 (.Y(N1421), .A(N1004), .B(N1005));
NAND2X4 inst_cellmath__201_0_I643 (.Y(N1422), .A(N1004), .B(N1005));
NOR2X2 inst_cellmath__201_0_I644 (.Y(N1423), .A(N1006), .B(N1007));
NAND2X4 inst_cellmath__201_0_I645 (.Y(N1424), .A(N1006), .B(N1007));
NOR2X1 inst_cellmath__201_0_I646 (.Y(N1425), .A(N1008), .B(N1009));
NAND2X2 inst_cellmath__201_0_I647 (.Y(N1426), .A(N1008), .B(N1009));
NOR2X2 inst_cellmath__201_0_I648 (.Y(N1427), .A(N1010), .B(N1011));
NAND2X2 inst_cellmath__201_0_I649 (.Y(N1428), .A(N1010), .B(N1011));
NOR2X1 inst_cellmath__201_0_I650 (.Y(N1429), .A(N1012), .B(N1013));
NAND2X2 inst_cellmath__201_0_I651 (.Y(N1430), .A(N1012), .B(N1013));
NOR2X1 inst_cellmath__201_0_I652 (.Y(N1431), .A(N1014), .B(N1015));
NAND2X2 inst_cellmath__201_0_I653 (.Y(N1432), .A(N1014), .B(N1015));
NOR2XL inst_cellmath__201_0_I654 (.Y(N1433), .A(N1016), .B(N1017));
NAND2X2 inst_cellmath__201_0_I655 (.Y(N1434), .A(N1016), .B(N1017));
NOR2XL inst_cellmath__201_0_I656 (.Y(N1435), .A(N1018), .B(N1019));
NAND2X1 inst_cellmath__201_0_I657 (.Y(N1436), .A(N1018), .B(N1019));
NOR2XL inst_cellmath__201_0_I658 (.Y(N1437), .A(N1021), .B(N1020));
NAND2XL inst_cellmath__201_0_I659 (.Y(N1438), .A(N1021), .B(N1020));
NOR2XL inst_cellmath__201_0_I660 (.Y(N1439), .A(N1022), .B(N1023));
NAND2XL inst_cellmath__201_0_I661 (.Y(N1440), .A(N1022), .B(N1023));
NOR2XL inst_cellmath__201_0_I662 (.Y(N1441), .A(N1024), .B(N1025));
NAND2XL inst_cellmath__201_0_I663 (.Y(N1442), .A(N1024), .B(N1025));
NOR2XL inst_cellmath__201_0_I664 (.Y(N1443), .A(N1027), .B(N1026));
NAND2XL inst_cellmath__201_0_I665 (.Y(N1444), .A(N1027), .B(N1026));
NOR2XL inst_cellmath__201_0_I666 (.Y(N1445), .A(N1029), .B(N1028));
NAND2XL inst_cellmath__201_0_I667 (.Y(N1446), .A(N1029), .B(N1028));
NOR2XL inst_cellmath__201_0_I668 (.Y(N1447), .A(N1031), .B(N1030));
NAND2XL inst_cellmath__201_0_I669 (.Y(N1448), .A(N1031), .B(N1030));
NOR2XL inst_cellmath__201_0_I670 (.Y(N1449), .A(N1033), .B(N1032));
NAND2XL inst_cellmath__201_0_I671 (.Y(N1450), .A(N1033), .B(N1032));
NOR2XL inst_cellmath__201_0_I672 (.Y(N1451), .A(N1035), .B(N1034));
NAND2XL inst_cellmath__201_0_I673 (.Y(N1452), .A(N1035), .B(N1034));
NOR2XL inst_cellmath__201_0_I674 (.Y(N1453), .A(N1037), .B(N1036));
NAND2XL inst_cellmath__201_0_I675 (.Y(N1454), .A(N1037), .B(N1036));
NOR2XL inst_cellmath__201_0_I676 (.Y(N1455), .A(N1039), .B(N1038));
NAND2XL inst_cellmath__201_0_I677 (.Y(N1456), .A(N1039), .B(N1038));
NOR2XL inst_cellmath__201_0_I678 (.Y(N1457), .A(N1040), .B(N1041));
NAND2XL inst_cellmath__201_0_I679 (.Y(N1458), .A(N1040), .B(N1041));
NOR2XL inst_cellmath__201_0_I680 (.Y(N1459), .A(N1042), .B(N1043));
NAND2XL inst_cellmath__201_0_I681 (.Y(N1460), .A(N1042), .B(N1043));
NOR2XL inst_cellmath__201_0_I682 (.Y(N1461), .A(N1045), .B(N1044));
NAND2XL inst_cellmath__201_0_I683 (.Y(N1462), .A(N1045), .B(N1044));
NOR2XL inst_cellmath__201_0_I684 (.Y(N1463), .A(N1047), .B(N1046));
NAND2XL inst_cellmath__201_0_I685 (.Y(N1464), .A(N1047), .B(N1046));
NOR2XL inst_cellmath__201_0_I686 (.Y(N1465), .A(N1049), .B(N1048));
NAND2XL inst_cellmath__201_0_I687 (.Y(N1466), .A(N1049), .B(N1048));
INVXL inst_cellmath__201_0_I1455 (.Y(N2421), .A(N1403));
AOI21X1 inst_cellmath__201_0_I691 (.Y(N1470), .A0(N1406), .A1(N1403), .B0(N1405));
AOI21XL inst_cellmath__201_0_I693 (.Y(N1472), .A0(N1408), .A1(N1405), .B0(N1407));
NAND2XL inst_cellmath__201_0_I694 (.Y(N1473), .A(N1408), .B(N1406));
AOI21X2 inst_cellmath__201_0_I695 (.Y(N1474), .A0(N1410), .A1(N1407), .B0(N1409));
NAND2X1 inst_cellmath__201_0_I696 (.Y(N1475), .A(N1410), .B(N1408));
AOI21X4 inst_cellmath__201_0_I697 (.Y(N1476), .A0(N1412), .A1(N1409), .B0(N1411));
NAND2X4 inst_cellmath__201_0_I698 (.Y(N1477), .A(N1412), .B(N1410));
AOI21X4 inst_cellmath__201_0_I699 (.Y(N1478), .A0(N1414), .A1(N1411), .B0(N1413));
NAND2X2 inst_cellmath__201_0_I700 (.Y(N1479), .A(N1414), .B(N1412));
AOI21X4 inst_cellmath__201_0_I701 (.Y(N1480), .A0(N1416), .A1(N1413), .B0(N1415));
NAND2X4 inst_cellmath__201_0_I702 (.Y(N1481), .A(N1416), .B(N1414));
AOI21X4 inst_cellmath__201_0_I703 (.Y(N1482), .A0(N1418), .A1(N1415), .B0(N1417));
NAND2X4 inst_cellmath__201_0_I704 (.Y(N1483), .A(N1418), .B(N1416));
AOI21X4 inst_cellmath__201_0_I705 (.Y(N1484), .A0(N1420), .A1(N1417), .B0(N1419));
NAND2X4 inst_cellmath__201_0_I706 (.Y(N1485), .A(N1420), .B(N1418));
AOI21X4 inst_cellmath__201_0_I707 (.Y(N1486), .A0(N1422), .A1(N1419), .B0(N1421));
NAND2X4 inst_cellmath__201_0_I708 (.Y(N1487), .A(N1422), .B(N1420));
AOI21X4 inst_cellmath__201_0_I709 (.Y(N1488), .A0(N1424), .A1(N1421), .B0(N1423));
NAND2X4 inst_cellmath__201_0_I710 (.Y(N1489), .A(N1424), .B(N1422));
AOI21X2 inst_cellmath__201_0_I711 (.Y(N1490), .A0(N1426), .A1(N1423), .B0(N1425));
NAND2X4 inst_cellmath__201_0_I712 (.Y(N1491), .A(N1426), .B(N1424));
AOI21X2 inst_cellmath__201_0_I713 (.Y(N1492), .A0(N1428), .A1(N1425), .B0(N1427));
NAND2X2 inst_cellmath__201_0_I714 (.Y(N1493), .A(N1428), .B(N1426));
AOI21X1 inst_cellmath__201_0_I715 (.Y(N1494), .A0(N1430), .A1(N1427), .B0(N1429));
NAND2X2 inst_cellmath__201_0_I716 (.Y(N1495), .A(N1430), .B(N1428));
AOI21X2 inst_cellmath__201_0_I717 (.Y(N1496), .A0(N1432), .A1(N1429), .B0(N1431));
NAND2X2 inst_cellmath__201_0_I718 (.Y(N1497), .A(N1432), .B(N1430));
AOI21X1 inst_cellmath__201_0_I719 (.Y(N1498), .A0(N1434), .A1(N1431), .B0(N1433));
NAND2X2 inst_cellmath__201_0_I720 (.Y(N1499), .A(N1434), .B(N1432));
AOI21X1 inst_cellmath__201_0_I721 (.Y(N1500), .A0(N1436), .A1(N1433), .B0(N1435));
NAND2X2 inst_cellmath__201_0_I722 (.Y(N1501), .A(N1436), .B(N1434));
AOI21XL inst_cellmath__201_0_I723 (.Y(N1502), .A0(N1438), .A1(N1435), .B0(N1437));
NAND2XL inst_cellmath__201_0_I724 (.Y(N1503), .A(N1438), .B(N1436));
AOI21XL inst_cellmath__201_0_I725 (.Y(N1504), .A0(N1440), .A1(N1437), .B0(N1439));
NAND2XL inst_cellmath__201_0_I726 (.Y(N1505), .A(N1440), .B(N1438));
AOI21XL inst_cellmath__201_0_I727 (.Y(N1506), .A0(N1442), .A1(N1439), .B0(N1441));
NAND2XL inst_cellmath__201_0_I728 (.Y(N1507), .A(N1442), .B(N1440));
AOI21XL inst_cellmath__201_0_I729 (.Y(N1508), .A0(N1444), .A1(N1441), .B0(N1443));
NAND2XL inst_cellmath__201_0_I730 (.Y(N1509), .A(N1444), .B(N1442));
AOI21XL inst_cellmath__201_0_I731 (.Y(N1510), .A0(N1446), .A1(N1443), .B0(N1445));
NAND2XL inst_cellmath__201_0_I732 (.Y(N1511), .A(N1446), .B(N1444));
AOI21XL inst_cellmath__201_0_I733 (.Y(N1512), .A0(N1448), .A1(N1445), .B0(N1447));
NAND2XL inst_cellmath__201_0_I734 (.Y(N1513), .A(N1448), .B(N1446));
AOI21XL inst_cellmath__201_0_I735 (.Y(N1514), .A0(N1450), .A1(N1447), .B0(N1449));
NAND2XL inst_cellmath__201_0_I736 (.Y(N1515), .A(N1450), .B(N1448));
AOI21XL inst_cellmath__201_0_I737 (.Y(N1516), .A0(N1452), .A1(N1449), .B0(N1451));
NAND2XL inst_cellmath__201_0_I738 (.Y(N1517), .A(N1452), .B(N1450));
AOI21XL inst_cellmath__201_0_I739 (.Y(N1518), .A0(N1454), .A1(N1451), .B0(N1453));
NAND2XL inst_cellmath__201_0_I740 (.Y(N1519), .A(N1454), .B(N1452));
AOI21XL inst_cellmath__201_0_I741 (.Y(N1520), .A0(N1456), .A1(N1453), .B0(N1455));
NAND2XL inst_cellmath__201_0_I742 (.Y(N1521), .A(N1456), .B(N1454));
AOI21XL inst_cellmath__201_0_I743 (.Y(N1522), .A0(N1458), .A1(N1455), .B0(N1457));
NAND2XL inst_cellmath__201_0_I744 (.Y(N1523), .A(N1458), .B(N1456));
AOI21XL inst_cellmath__201_0_I745 (.Y(N1524), .A0(N1460), .A1(N1457), .B0(N1459));
NAND2XL inst_cellmath__201_0_I746 (.Y(N1525), .A(N1460), .B(N1458));
AOI21XL inst_cellmath__201_0_I747 (.Y(N1526), .A0(N1462), .A1(N1459), .B0(N1461));
NAND2XL inst_cellmath__201_0_I748 (.Y(N1527), .A(N1462), .B(N1460));
AOI21XL inst_cellmath__201_0_I749 (.Y(N1528), .A0(N1464), .A1(N1461), .B0(N1463));
NAND2XL inst_cellmath__201_0_I750 (.Y(N1529), .A(N1464), .B(N1462));
AOI21XL inst_cellmath__201_0_I751 (.Y(N1530), .A0(N1466), .A1(N1463), .B0(N1465));
NAND2XL inst_cellmath__201_0_I752 (.Y(N1531), .A(N1466), .B(N1464));
NAND2XL inst_cellmath__201_0_I754 (.Y(N1534), .A(N1049), .B(N1466));
INVXL inst_cellmath__201_0_I1456 (.Y(N2422), .A(N2421));
INVXL inst_cellmath__201_0_I1457 (.Y(N2423), .A(N1470));
OAI21X1 inst_cellmath__201_0_I759 (.Y(N1539), .A0(N1473), .A1(N2421), .B0(N1472));
OAI21X1 inst_cellmath__201_0_I761 (.Y(N1541), .A0(N1475), .A1(N1470), .B0(N1474));
OAI21X4 inst_cellmath__201_0_I763 (.Y(N1543), .A0(N1477), .A1(N1472), .B0(N1476));
NOR2X4 inst_cellmath__201_0_I764 (.Y(N1544), .A(N1477), .B(N1473));
OAI21X2 inst_cellmath__201_0_I765 (.Y(N1545), .A0(N1479), .A1(N1474), .B0(N1478));
NOR2X2 inst_cellmath__201_0_I766 (.Y(N1546), .A(N1479), .B(N1475));
OAI21X2 inst_cellmath__201_0_I767 (.Y(N1547), .A0(N1481), .A1(N1476), .B0(N1480));
NOR2X2 inst_cellmath__201_0_I768 (.Y(N1548), .A(N1481), .B(N1477));
OAI21X4 inst_cellmath__201_0_I769 (.Y(N1549), .A0(N1483), .A1(N1478), .B0(N1482));
NOR2X2 inst_cellmath__201_0_I770 (.Y(N1550), .A(N1483), .B(N1479));
OAI21X4 inst_cellmath__201_0_I771 (.Y(N1551), .A0(N1485), .A1(N1480), .B0(N1484));
NOR2X4 inst_cellmath__201_0_I772 (.Y(N1552), .A(N1485), .B(N1481));
OAI21X2 inst_cellmath__201_0_I773 (.Y(N1553), .A0(N1487), .A1(N1482), .B0(N1486));
NOR2X2 inst_cellmath__201_0_I774 (.Y(N1554), .A(N1487), .B(N1483));
OAI21X4 inst_cellmath__201_0_I775 (.Y(N1555), .A0(N1489), .A1(N1484), .B0(N1488));
NOR2X2 inst_cellmath__201_0_I776 (.Y(N1556), .A(N1489), .B(N1485));
OAI21X4 inst_cellmath__201_0_I777 (.Y(N1557), .A0(N1491), .A1(N1486), .B0(N1490));
NOR2X2 inst_cellmath__201_0_I778 (.Y(N1558), .A(N1491), .B(N1487));
OAI21X4 inst_cellmath__201_0_I779 (.Y(N1559), .A0(N1493), .A1(N1488), .B0(N1492));
NOR2X4 inst_cellmath__201_0_I780 (.Y(N1560), .A(N1493), .B(N1489));
OAI21X2 inst_cellmath__201_0_I781 (.Y(N1561), .A0(N1495), .A1(N1490), .B0(N1494));
NOR2X2 inst_cellmath__201_0_I782 (.Y(N1562), .A(N1495), .B(N1491));
OAI21X2 inst_cellmath__201_0_I783 (.Y(N1563), .A0(N1497), .A1(N1492), .B0(N1496));
NOR2X2 inst_cellmath__201_0_I784 (.Y(N1564), .A(N1497), .B(N1493));
OAI21X2 inst_cellmath__201_0_I785 (.Y(N1565), .A0(N1499), .A1(N1494), .B0(N1498));
NOR2X2 inst_cellmath__201_0_I786 (.Y(N1566), .A(N1499), .B(N1495));
OAI21X2 inst_cellmath__201_0_I787 (.Y(N1567), .A0(N1501), .A1(N1496), .B0(N1500));
NOR2X2 inst_cellmath__201_0_I788 (.Y(N1568), .A(N1501), .B(N1497));
OAI21X1 inst_cellmath__201_0_I789 (.Y(N1569), .A0(N1503), .A1(N1498), .B0(N1502));
NOR2X1 inst_cellmath__201_0_I790 (.Y(N1570), .A(N1503), .B(N1499));
OAI21X1 inst_cellmath__201_0_I791 (.Y(N1571), .A0(N1505), .A1(N1500), .B0(N1504));
NOR2X1 inst_cellmath__201_0_I792 (.Y(N1572), .A(N1505), .B(N1501));
OAI21XL inst_cellmath__201_0_I793 (.Y(N1573), .A0(N1507), .A1(N1502), .B0(N1506));
NOR2XL inst_cellmath__201_0_I794 (.Y(N1574), .A(N1507), .B(N1503));
OAI21XL inst_cellmath__201_0_I795 (.Y(N1575), .A0(N1509), .A1(N1504), .B0(N1508));
NOR2XL inst_cellmath__201_0_I796 (.Y(N1576), .A(N1509), .B(N1505));
OAI21XL inst_cellmath__201_0_I797 (.Y(N1577), .A0(N1511), .A1(N1506), .B0(N1510));
NOR2XL inst_cellmath__201_0_I798 (.Y(N1578), .A(N1511), .B(N1507));
OAI21XL inst_cellmath__201_0_I799 (.Y(N1579), .A0(N1513), .A1(N1508), .B0(N1512));
NOR2XL inst_cellmath__201_0_I800 (.Y(N1580), .A(N1513), .B(N1509));
OAI21XL inst_cellmath__201_0_I801 (.Y(N1581), .A0(N1515), .A1(N1510), .B0(N1514));
NOR2XL inst_cellmath__201_0_I802 (.Y(N1582), .A(N1515), .B(N1511));
OAI21XL inst_cellmath__201_0_I803 (.Y(N1583), .A0(N1517), .A1(N1512), .B0(N1516));
NOR2XL inst_cellmath__201_0_I804 (.Y(N1584), .A(N1517), .B(N1513));
OAI21XL inst_cellmath__201_0_I805 (.Y(N1585), .A0(N1519), .A1(N1514), .B0(N1518));
NOR2XL inst_cellmath__201_0_I806 (.Y(N1586), .A(N1519), .B(N1515));
OAI21XL inst_cellmath__201_0_I807 (.Y(N1587), .A0(N1521), .A1(N1516), .B0(N1520));
NOR2XL inst_cellmath__201_0_I808 (.Y(N1588), .A(N1521), .B(N1517));
OAI21XL inst_cellmath__201_0_I809 (.Y(N1589), .A0(N1523), .A1(N1518), .B0(N1522));
NOR2XL inst_cellmath__201_0_I810 (.Y(N1590), .A(N1523), .B(N1519));
OAI21XL inst_cellmath__201_0_I811 (.Y(N1591), .A0(N1525), .A1(N1520), .B0(N1524));
NOR2XL inst_cellmath__201_0_I812 (.Y(N1592), .A(N1525), .B(N1521));
OAI21XL inst_cellmath__201_0_I813 (.Y(N1593), .A0(N1527), .A1(N1522), .B0(N1526));
NOR2XL inst_cellmath__201_0_I814 (.Y(N1594), .A(N1527), .B(N1523));
OAI21XL inst_cellmath__201_0_I815 (.Y(N1595), .A0(N1529), .A1(N1524), .B0(N1528));
NOR2XL inst_cellmath__201_0_I816 (.Y(N1596), .A(N1529), .B(N1525));
OAI21XL inst_cellmath__201_0_I817 (.Y(N1597), .A0(N1531), .A1(N1526), .B0(N1530));
NOR2XL inst_cellmath__201_0_I818 (.Y(N1598), .A(N1531), .B(N1527));
OAI2BB2XL inst_cellmath__201_0_I1295 (.Y(N1599), .A0N(N1049), .A1N(N1465), .B0(N1534), .B1(N1528));
NOR2XL inst_cellmath__201_0_I820 (.Y(N1600), .A(N1534), .B(N1529));
INVXL inst_cellmath__201_0_I1458 (.Y(N2424), .A(N2422));
INVXL inst_cellmath__201_0_I1459 (.Y(N2425), .A(N2423));
INVXL inst_cellmath__201_0_I1460 (.Y(N2426), .A(N1539));
INVX1 inst_cellmath__201_0_I1461 (.Y(N2427), .A(N1541));
AOI21X2 inst_cellmath__201_0_I829 (.Y(N1609), .A0(N1544), .A1(N2422), .B0(N1543));
AOI21X1 inst_cellmath__201_0_I831 (.Y(N1611), .A0(N1546), .A1(N2423), .B0(N1545));
AOI21X1 inst_cellmath__201_0_I833 (.Y(N1613), .A0(N1548), .A1(N1539), .B0(N1547));
AOI21X1 inst_cellmath__201_0_I835 (.Y(N1615), .A0(N1550), .A1(N1541), .B0(N1549));
AOI21X4 inst_cellmath__201_0_I837 (.Y(N1617), .A0(N1552), .A1(N1543), .B0(N1551));
NAND2X2 inst_cellmath__201_0_I838 (.Y(N1618), .A(N1552), .B(N1544));
AOI21X1 inst_cellmath__201_0_I839 (.Y(N1619), .A0(N1554), .A1(N1545), .B0(N1553));
NAND2XL inst_cellmath__201_0_I840 (.Y(N1620), .A(N1554), .B(N1546));
AOI21X1 inst_cellmath__201_0_I841 (.Y(N1621), .A0(N1556), .A1(N1547), .B0(N1555));
NAND2XL inst_cellmath__201_0_I842 (.Y(N1622), .A(N1556), .B(N1548));
AOI21X4 inst_cellmath__201_0_I843 (.Y(N1623), .A0(N1558), .A1(N1549), .B0(N1557));
NAND2X1 inst_cellmath__201_0_I844 (.Y(N1624), .A(N1558), .B(N1550));
AOI21X4 inst_cellmath__201_0_I845 (.Y(N1625), .A0(N1560), .A1(N1551), .B0(N1559));
NAND2X2 inst_cellmath__201_0_I846 (.Y(N1626), .A(N1560), .B(N1552));
AOI21X2 inst_cellmath__201_0_I847 (.Y(N1627), .A0(N1562), .A1(N1553), .B0(N1561));
NAND2X1 inst_cellmath__201_0_I848 (.Y(N1628), .A(N1562), .B(N1554));
AOI21X2 inst_cellmath__201_0_I849 (.Y(N1629), .A0(N1564), .A1(N1555), .B0(N1563));
NAND2X1 inst_cellmath__201_0_I850 (.Y(N1630), .A(N1564), .B(N1556));
AOI21X1 inst_cellmath__201_0_I851 (.Y(N1631), .A0(N1566), .A1(N1557), .B0(N1565));
NAND2XL inst_cellmath__201_0_I852 (.Y(N1632), .A(N1566), .B(N1558));
AOI21X2 inst_cellmath__201_0_I853 (.Y(N1633), .A0(N1568), .A1(N1559), .B0(N1567));
NAND2X2 inst_cellmath__201_0_I854 (.Y(N1634), .A(N1568), .B(N1560));
AOI21XL inst_cellmath__201_0_I855 (.Y(N1635), .A0(N1570), .A1(N1561), .B0(N1569));
NAND2XL inst_cellmath__201_0_I856 (.Y(N1636), .A(N1570), .B(N1562));
AOI21X1 inst_cellmath__201_0_I857 (.Y(N1637), .A0(N1572), .A1(N1563), .B0(N1571));
NAND2X1 inst_cellmath__201_0_I858 (.Y(N1638), .A(N1572), .B(N1564));
AOI21XL inst_cellmath__201_0_I859 (.Y(N1639), .A0(N1574), .A1(N1565), .B0(N1573));
NAND2XL inst_cellmath__201_0_I860 (.Y(N1640), .A(N1574), .B(N1566));
AOI21XL inst_cellmath__201_0_I861 (.Y(N1641), .A0(N1576), .A1(N1567), .B0(N1575));
NAND2XL inst_cellmath__201_0_I862 (.Y(N1642), .A(N1576), .B(N1568));
AOI21XL inst_cellmath__201_0_I863 (.Y(N1643), .A0(N1578), .A1(N1569), .B0(N1577));
NAND2XL inst_cellmath__201_0_I864 (.Y(N1644), .A(N1578), .B(N1570));
AOI21XL inst_cellmath__201_0_I865 (.Y(N1645), .A0(N1580), .A1(N1571), .B0(N1579));
NAND2XL inst_cellmath__201_0_I866 (.Y(N1646), .A(N1580), .B(N1572));
AOI21XL inst_cellmath__201_0_I867 (.Y(N1647), .A0(N1582), .A1(N1573), .B0(N1581));
NAND2XL inst_cellmath__201_0_I868 (.Y(N1648), .A(N1582), .B(N1574));
AOI21XL inst_cellmath__201_0_I869 (.Y(N1649), .A0(N1584), .A1(N1575), .B0(N1583));
NAND2XL inst_cellmath__201_0_I870 (.Y(N1650), .A(N1584), .B(N1576));
AOI21XL inst_cellmath__201_0_I871 (.Y(N1651), .A0(N1586), .A1(N1577), .B0(N1585));
NAND2XL inst_cellmath__201_0_I872 (.Y(N1652), .A(N1586), .B(N1578));
AOI21XL inst_cellmath__201_0_I873 (.Y(N1653), .A0(N1588), .A1(N1579), .B0(N1587));
NAND2XL inst_cellmath__201_0_I874 (.Y(N1654), .A(N1588), .B(N1580));
AOI21XL inst_cellmath__201_0_I875 (.Y(N1655), .A0(N1590), .A1(N1581), .B0(N1589));
NAND2XL inst_cellmath__201_0_I876 (.Y(N1656), .A(N1590), .B(N1582));
AOI21XL inst_cellmath__201_0_I877 (.Y(N1657), .A0(N1592), .A1(N1583), .B0(N1591));
NAND2XL inst_cellmath__201_0_I878 (.Y(N1658), .A(N1592), .B(N1584));
AOI21XL inst_cellmath__201_0_I879 (.Y(N1659), .A0(N1594), .A1(N1585), .B0(N1593));
NAND2XL inst_cellmath__201_0_I880 (.Y(N1660), .A(N1594), .B(N1586));
AOI21XL inst_cellmath__201_0_I881 (.Y(N1661), .A0(N1596), .A1(N1587), .B0(N1595));
NAND2XL inst_cellmath__201_0_I882 (.Y(N1662), .A(N1596), .B(N1588));
AOI21XL inst_cellmath__201_0_I883 (.Y(N1663), .A0(N1598), .A1(N1589), .B0(N1597));
NAND2XL inst_cellmath__201_0_I884 (.Y(N1664), .A(N1598), .B(N1590));
AOI21XL inst_cellmath__201_0_I885 (.Y(N1665), .A0(N1600), .A1(N1591), .B0(N1599));
NAND2XL inst_cellmath__201_0_I886 (.Y(N1666), .A(N1600), .B(N1592));
INVXL inst_cellmath__201_0_I1462 (.Y(N2428), .A(N2424));
INVXL inst_cellmath__201_0_I1463 (.Y(N2429), .A(N2425));
INVXL inst_cellmath__201_0_I1464 (.Y(N2430), .A(N2426));
INVXL inst_cellmath__201_0_I1465 (.Y(N2431), .A(N2427));
INVXL inst_cellmath__201_0_I1466 (.Y(N2432), .A(N1609));
INVXL inst_cellmath__201_0_I1467 (.Y(N2433), .A(N1611));
INVXL inst_cellmath__201_0_I1468 (.Y(N2434), .A(N1613));
INVXL inst_cellmath__201_0_I1469 (.Y(N2435), .A(N1615));
OAI21XL inst_cellmath__201_0_I903 (.Y(N1683), .A0(N1618), .A1(N2424), .B0(N1617));
OAI21XL inst_cellmath__201_0_I905 (.Y(N1685), .A0(N1620), .A1(N2425), .B0(N1619));
OAI21XL inst_cellmath__201_0_I907 (.Y(N1687), .A0(N1622), .A1(N2426), .B0(N1621));
OAI21XL inst_cellmath__201_0_I909 (.Y(N1689), .A0(N1624), .A1(N2427), .B0(N1623));
OAI21X1 inst_cellmath__201_0_I911 (.Y(N1691), .A0(N1626), .A1(N1609), .B0(N1625));
OAI21X1 inst_cellmath__201_0_I913 (.Y(N1693), .A0(N1628), .A1(N1611), .B0(N1627));
OAI21X1 inst_cellmath__201_0_I915 (.Y(N1695), .A0(N1630), .A1(N1613), .B0(N1629));
OAI21XL inst_cellmath__201_0_I917 (.Y(N1697), .A0(N1632), .A1(N1615), .B0(N1631));
OAI21X2 inst_cellmath__201_0_I919 (.Y(N1699), .A0(N1634), .A1(N1617), .B0(N1633));
NOR2X1 inst_cellmath__201_0_I920 (.Y(N1700), .A(N1634), .B(N1618));
OAI21XL inst_cellmath__201_0_I921 (.Y(N1701), .A0(N1636), .A1(N1619), .B0(N1635));
NOR2XL inst_cellmath__201_0_I922 (.Y(N1702), .A(N1636), .B(N1620));
OAI21XL inst_cellmath__201_0_I923 (.Y(N1703), .A0(N1638), .A1(N1621), .B0(N1637));
NOR2XL inst_cellmath__201_0_I924 (.Y(N1704), .A(N1638), .B(N1622));
OAI21XL inst_cellmath__201_0_I925 (.Y(N1705), .A0(N1640), .A1(N1623), .B0(N1639));
NOR2XL inst_cellmath__201_0_I926 (.Y(N1706), .A(N1640), .B(N1624));
OAI21XL inst_cellmath__201_0_I927 (.Y(N1707), .A0(N1642), .A1(N1625), .B0(N1641));
NOR2XL inst_cellmath__201_0_I928 (.Y(N1708), .A(N1642), .B(N1626));
OAI21X1 inst_cellmath__201_0_I929 (.Y(N1709), .A0(N1644), .A1(N1627), .B0(N1643));
NOR2XL inst_cellmath__201_0_I930 (.Y(N1710), .A(N1644), .B(N1628));
OAI21XL inst_cellmath__201_0_I931 (.Y(N1711), .A0(N1646), .A1(N1629), .B0(N1645));
NOR2XL inst_cellmath__201_0_I932 (.Y(N1712), .A(N1646), .B(N1630));
OAI21XL inst_cellmath__201_0_I933 (.Y(N1713), .A0(N1648), .A1(N1631), .B0(N1647));
NOR2XL inst_cellmath__201_0_I934 (.Y(N1714), .A(N1648), .B(N1632));
OAI21XL inst_cellmath__201_0_I935 (.Y(N1715), .A0(N1650), .A1(N1633), .B0(N1649));
NOR2XL inst_cellmath__201_0_I936 (.Y(N1716), .A(N1650), .B(N1634));
OAI21XL inst_cellmath__201_0_I937 (.Y(N1717), .A0(N1652), .A1(N1635), .B0(N1651));
NOR2XL inst_cellmath__201_0_I938 (.Y(N1718), .A(N1652), .B(N1636));
OAI21XL inst_cellmath__201_0_I939 (.Y(N1719), .A0(N1654), .A1(N1637), .B0(N1653));
NOR2XL inst_cellmath__201_0_I940 (.Y(N1720), .A(N1654), .B(N1638));
OAI21XL inst_cellmath__201_0_I941 (.Y(N1721), .A0(N1656), .A1(N1639), .B0(N1655));
NOR2XL inst_cellmath__201_0_I942 (.Y(N1722), .A(N1656), .B(N1640));
OAI21XL inst_cellmath__201_0_I943 (.Y(N1723), .A0(N1658), .A1(N1641), .B0(N1657));
NOR2XL inst_cellmath__201_0_I944 (.Y(N1724), .A(N1658), .B(N1642));
OAI21XL inst_cellmath__201_0_I945 (.Y(N1725), .A0(N1660), .A1(N1643), .B0(N1659));
NOR2XL inst_cellmath__201_0_I946 (.Y(N1726), .A(N1660), .B(N1644));
OAI21XL inst_cellmath__201_0_I947 (.Y(N1727), .A0(N1662), .A1(N1645), .B0(N1661));
NOR2XL inst_cellmath__201_0_I948 (.Y(N1728), .A(N1662), .B(N1646));
OAI21XL inst_cellmath__201_0_I949 (.Y(N1729), .A0(N1664), .A1(N1647), .B0(N1663));
NOR2XL inst_cellmath__201_0_I950 (.Y(N1730), .A(N1664), .B(N1648));
OAI21XL inst_cellmath__201_0_I951 (.Y(N1731), .A0(N1666), .A1(N1649), .B0(N1665));
NOR2XL inst_cellmath__201_0_I952 (.Y(N1732), .A(N1666), .B(N1650));
INVXL inst_cellmath__201_0_I1472 (.Y(N2438), .A(N2428));
AOI21XL inst_cellmath__201_0_I985 (.Y(N1765), .A0(N1700), .A1(N2428), .B0(N1699));
AOI21XL inst_cellmath__201_0_I987 (.Y(N1767), .A0(N1702), .A1(N2429), .B0(N1701));
AOI21XL inst_cellmath__201_0_I989 (.Y(N1769), .A0(N1704), .A1(N2430), .B0(N1703));
AOI21XL inst_cellmath__201_0_I991 (.Y(N1771), .A0(N1706), .A1(N2431), .B0(N1705));
AOI21XL inst_cellmath__201_0_I993 (.Y(N1773), .A0(N1708), .A1(N2432), .B0(N1707));
AOI21X1 inst_cellmath__201_0_I995 (.Y(N1775), .A0(N1710), .A1(N2433), .B0(N1709));
AOI21X1 inst_cellmath__201_0_I997 (.Y(N1777), .A0(N1712), .A1(N2434), .B0(N1711));
AOI21XL inst_cellmath__201_0_I999 (.Y(N1779), .A0(N1714), .A1(N2435), .B0(N1713));
AOI21XL inst_cellmath__201_0_I1001 (.Y(N1781), .A0(N1716), .A1(N1683), .B0(N1715));
AOI21XL inst_cellmath__201_0_I1003 (.Y(N1783), .A0(N1718), .A1(N1685), .B0(N1717));
AOI21XL inst_cellmath__201_0_I1005 (.Y(N1785), .A0(N1720), .A1(N1687), .B0(N1719));
AOI21XL inst_cellmath__201_0_I1007 (.Y(N1787), .A0(N1722), .A1(N1689), .B0(N1721));
AOI21XL inst_cellmath__201_0_I1009 (.Y(N1789), .A0(N1724), .A1(N1691), .B0(N1723));
AOI21XL inst_cellmath__201_0_I1011 (.Y(N1791), .A0(N1726), .A1(N1693), .B0(N1725));
AOI21XL inst_cellmath__201_0_I1013 (.Y(N1793), .A0(N1728), .A1(N1695), .B0(N1727));
AOI21X2 inst_cellmath__201_0_I1017 (.Y(N1797), .A0(N1732), .A1(N1699), .B0(N1731));
NAND2X1 inst_cellmath__201_0_I1018 (.Y(N1798), .A(N1732), .B(N1700));
AO21XL inst_cellmath__201_0_I1516 (.Y(N2456), .A0(N1730), .A1(N1697), .B0(N1729));
OAI21X4 inst_cellmath__201_0_I1083 (.Y(inst_cellmath__201_0_out0[49]), .A0(N1798), .A1(N2438), .B0(N1797));
NAND2BXL inst_cellmath__201_0_I1090 (.Y(N1870), .AN(N1405), .B(N1406));
NAND2BXL inst_cellmath__201_0_I1093 (.Y(N1873), .AN(N1407), .B(N1408));
NAND2BXL inst_cellmath__201_0_I1096 (.Y(N1876), .AN(N1409), .B(N1410));
NAND2BXL inst_cellmath__201_0_I1099 (.Y(N1879), .AN(N1411), .B(N1412));
NAND2BXL inst_cellmath__201_0_I1102 (.Y(N1882), .AN(N1413), .B(N1414));
NAND2BXL inst_cellmath__201_0_I1105 (.Y(N1885), .AN(N1415), .B(N1416));
NAND2BXL inst_cellmath__201_0_I1108 (.Y(N1888), .AN(N1417), .B(N1418));
NAND2BXL inst_cellmath__201_0_I1111 (.Y(N1891), .AN(N1419), .B(N1420));
NAND2BXL inst_cellmath__201_0_I1114 (.Y(N1894), .AN(N1421), .B(N1422));
NAND2BXL inst_cellmath__201_0_I1117 (.Y(N1897), .AN(N1423), .B(N1424));
NAND2BXL inst_cellmath__201_0_I1120 (.Y(N1900), .AN(N1425), .B(N1426));
NAND2BXL inst_cellmath__201_0_I1123 (.Y(N1903), .AN(N1427), .B(N1428));
NAND2BXL inst_cellmath__201_0_I1126 (.Y(N1906), .AN(N1429), .B(N1430));
NAND2BXL inst_cellmath__201_0_I1129 (.Y(N1909), .AN(N1431), .B(N1432));
NAND2BXL inst_cellmath__201_0_I1132 (.Y(N1912), .AN(N1433), .B(N1434));
NAND2BXL inst_cellmath__201_0_I1135 (.Y(N1915), .AN(N1435), .B(N1436));
NAND2BXL inst_cellmath__201_0_I1138 (.Y(N1918), .AN(N1437), .B(N1438));
NAND2BXL inst_cellmath__201_0_I1141 (.Y(N1921), .AN(N1439), .B(N1440));
NAND2BXL inst_cellmath__201_0_I1144 (.Y(N1924), .AN(N1441), .B(N1442));
NAND2BXL inst_cellmath__201_0_I1147 (.Y(N1927), .AN(N1443), .B(N1444));
NAND2BXL inst_cellmath__201_0_I1150 (.Y(N1930), .AN(N1445), .B(N1446));
NAND2BXL inst_cellmath__201_0_I1153 (.Y(N1933), .AN(N1447), .B(N1448));
NAND2BXL inst_cellmath__201_0_I1156 (.Y(N1936), .AN(N1449), .B(N1450));
NAND2BXL inst_cellmath__201_0_I1159 (.Y(N1939), .AN(N1451), .B(N1452));
NAND2BXL inst_cellmath__201_0_I1162 (.Y(N1942), .AN(N1453), .B(N1454));
NAND2BXL inst_cellmath__201_0_I1165 (.Y(N1945), .AN(N1455), .B(N1456));
NAND2BXL inst_cellmath__201_0_I1168 (.Y(N1948), .AN(N1457), .B(N1458));
NAND2BXL inst_cellmath__201_0_I1171 (.Y(N1951), .AN(N1459), .B(N1460));
NAND2BXL inst_cellmath__201_0_I1174 (.Y(N1954), .AN(N1461), .B(N1462));
NAND2BXL inst_cellmath__201_0_I1177 (.Y(N1957), .AN(N1463), .B(N1464));
NAND2BXL inst_cellmath__201_0_I1180 (.Y(N1960), .AN(N1465), .B(N1466));
XNOR2X1 inst_cellmath__201_0_I1185 (.Y(inst_cellmath__201_0_out0[17]), .A(N2438), .B(N1870));
XOR2XL inst_cellmath__201_0_I1517 (.Y(inst_cellmath__201_0_out0[18]), .A(N2429), .B(N1873));
XOR2XL inst_cellmath__201_0_I1518 (.Y(inst_cellmath__201_0_out0[19]), .A(N2430), .B(N1876));
XOR2XL inst_cellmath__201_0_I1519 (.Y(inst_cellmath__201_0_out0[20]), .A(N2431), .B(N1879));
XOR2XL inst_cellmath__201_0_I1520 (.Y(inst_cellmath__201_0_out0[21]), .A(N2432), .B(N1882));
XOR2XL inst_cellmath__201_0_I1521 (.Y(inst_cellmath__201_0_out0[22]), .A(N2433), .B(N1885));
XOR2XL inst_cellmath__201_0_I1522 (.Y(inst_cellmath__201_0_out0[23]), .A(N2434), .B(N1888));
XOR2XL inst_cellmath__201_0_I1523 (.Y(inst_cellmath__201_0_out0[24]), .A(N2435), .B(N1891));
XOR2XL inst_cellmath__201_0_I1524 (.Y(inst_cellmath__201_0_out0[25]), .A(N1683), .B(N1894));
XOR2XL inst_cellmath__201_0_I1598 (.Y(inst_cellmath__201_0_out0[26]), .A(N1685), .B(N1897));
XOR2XL inst_cellmath__201_0_I1526 (.Y(inst_cellmath__201_0_out0[27]), .A(N1687), .B(N1900));
XOR2XL inst_cellmath__201_0_I2744 (.Y(inst_cellmath__201_0_out0[28]), .A(N1689), .B(N1903));
XOR2XL inst_cellmath__201_0_I2745 (.Y(inst_cellmath__201_0_out0[29]), .A(N1691), .B(N1906));
XOR2XL inst_cellmath__201_0_I2727 (.Y(inst_cellmath__201_0_out0[30]), .A(N1693), .B(N1909));
XOR2XL inst_cellmath__201_0_I2746 (.Y(inst_cellmath__201_0_out0[31]), .A(N1695), .B(N1912));
XOR2XL inst_cellmath__201_0_I1602 (.Y(inst_cellmath__201_0_out0[32]), .A(N1697), .B(N1915));
XNOR2X1 inst_cellmath__201_0_I2729 (.Y(inst_cellmath__201_0_out0[33]), .A(N1765), .B(N1918));
XNOR2XL inst_cellmath__201_0_I2730 (.Y(inst_cellmath__201_0_out0[34]), .A(N1767), .B(N1921));
XNOR2X1 inst_cellmath__201_0_I2731 (.Y(inst_cellmath__201_0_out0[35]), .A(N1769), .B(N1924));
XNOR2X1 inst_cellmath__201_0_I2732 (.Y(inst_cellmath__201_0_out0[36]), .A(N1771), .B(N1927));
XNOR2XL inst_cellmath__201_0_I2733 (.Y(inst_cellmath__201_0_out0[37]), .A(N1773), .B(N1930));
XNOR2X1 inst_cellmath__201_0_I2734 (.Y(inst_cellmath__201_0_out0[38]), .A(N1775), .B(N1933));
XNOR2X1 inst_cellmath__201_0_I2735 (.Y(inst_cellmath__201_0_out0[39]), .A(N1777), .B(N1936));
XNOR2X1 inst_cellmath__201_0_I1208 (.Y(inst_cellmath__201_0_out0[40]), .A(N1779), .B(N1939));
XNOR2XL inst_cellmath__201_0_I2736 (.Y(inst_cellmath__201_0_out0[41]), .A(N1781), .B(N1942));
XNOR2X1 inst_cellmath__201_0_I2737 (.Y(inst_cellmath__201_0_out0[42]), .A(N1783), .B(N1945));
XNOR2X1 inst_cellmath__201_0_I2738 (.Y(inst_cellmath__201_0_out0[43]), .A(N1785), .B(N1948));
XNOR2X1 inst_cellmath__201_0_I2739 (.Y(inst_cellmath__201_0_out0[44]), .A(N1787), .B(N1951));
XNOR2X1 inst_cellmath__201_0_I2740 (.Y(inst_cellmath__201_0_out0[45]), .A(N1789), .B(N1954));
XNOR2X1 inst_cellmath__201_0_I2741 (.Y(inst_cellmath__201_0_out0[46]), .A(N1791), .B(N1957));
XNOR2X1 inst_cellmath__201_0_I2742 (.Y(inst_cellmath__201_0_out0[47]), .A(N1793), .B(N1960));
XNOR2X1 inst_cellmath__201_0_I1216 (.Y(inst_cellmath__201_0_out0[48]), .A(N2456), .B(N1049));
assign inst_cellmath__203__W1[0] = inst_cellmath__201_0_in1[0];
assign inst_cellmath__203__W1[1] = inst_cellmath__201_0_in0[1];
assign inst_cellmath__203__W1[2] = inst_cellmath__201_0_in0[2];
assign inst_cellmath__203__W1[3] = inst_cellmath__201_0_in0[3];
assign inst_cellmath__203__W1[4] = inst_cellmath__201_0_in0[4];
assign inst_cellmath__203__W1[5] = inst_cellmath__201_0_in0[5];
assign inst_cellmath__203__W1[6] = inst_cellmath__201_0_in0[6];
assign inst_cellmath__203__W1[7] = inst_cellmath__201_0_in0[7];
assign inst_cellmath__203__W1[8] = inst_cellmath__201_0_in0[8];
assign inst_cellmath__203__W1[9] = inst_cellmath__201_0_in0[9];
assign inst_cellmath__203__W1[10] = inst_cellmath__201_0_in0[10];
assign inst_cellmath__203__W1[11] = inst_cellmath__201_0_in0[11];
assign inst_cellmath__203__W1[12] = inst_cellmath__201_0_in0[12];
assign inst_cellmath__203__W1[13] = inst_cellmath__201_0_in0[13];
assign inst_cellmath__203__W1[14] = inst_cellmath__201_0_in0[14];
assign inst_cellmath__203__W1[15] = inst_cellmath__201_0_in0[15];
assign inst_cellmath__203__W1[16] = inst_cellmath__201_0_in0[16];
assign inst_cellmath__203__W1[17] = inst_cellmath__201_0_in0[17];
assign inst_cellmath__203__W1[18] = inst_cellmath__201_0_in0[18];
assign inst_cellmath__203__W1[19] = inst_cellmath__201_0_in0[19];
assign inst_cellmath__203__W1[20] = inst_cellmath__201_0_in0[20];
assign inst_cellmath__203__W1[21] = inst_cellmath__201_0_in0[21];
assign inst_cellmath__203__W1[22] = inst_cellmath__201_0_in0[22];
assign inst_cellmath__203__W1[23] = inst_cellmath__201_0_in0[23];
assign inst_cellmath__203__W1[24] = inst_cellmath__201_0_in0[24];
assign inst_cellmath__203__W1[25] = inst_cellmath__201_0_in0[25];
assign inst_cellmath__203__W1[26] = inst_cellmath__201_0_in0[26];
assign inst_cellmath__203__W1[27] = inst_cellmath__201_0_in0[27];
assign inst_cellmath__203__W1[28] = inst_cellmath__201_0_in0[28];
assign inst_cellmath__203__W1[29] = inst_cellmath__201_0_in0[29];
assign inst_cellmath__203__W1[30] = inst_cellmath__201_0_in0[30];
assign inst_cellmath__203__W1[31] = inst_cellmath__201_0_in0[31];
assign inst_cellmath__203__W1[32] = inst_cellmath__201_0_in0[32];
assign inst_cellmath__203__W1[33] = inst_cellmath__201_0_in1[33];
assign inst_cellmath__203__W1[34] = inst_cellmath__201_0_in0[34];
assign inst_cellmath__203__W1[35] = inst_cellmath__201_0_in1[35];
assign inst_cellmath__203__W1[36] = inst_cellmath__201_0_in0[36];
assign inst_cellmath__203__W1[37] = inst_cellmath__201_0_in0[37];
assign inst_cellmath__203__W1[38] = inst_cellmath__201_0_in0[38];
assign inst_cellmath__203__W1[39] = inst_cellmath__201_0_in0[39];
assign inst_cellmath__203__W1[40] = inst_cellmath__201_0_in0[40];
assign inst_cellmath__203__W1[41] = inst_cellmath__201_0_in0[41];
assign inst_cellmath__203__W1[42] = inst_cellmath__201_0_in0[42];
assign inst_cellmath__203__W1[43] = inst_cellmath__201_0_in0[43];
assign inst_cellmath__203__W1[44] = inst_cellmath__201_0_in0[44];
assign inst_cellmath__203__W1[45] = inst_cellmath__201_0_in0[45];
endmodule

module cynw_cm_float_cos_inst_cellmath__200_0_bdw1157874770_bdw (
	inst_cellmath__200_0_out0,
	inst_cellmath__200_0_in0
	); /* architecture "gate_level" */ 
output [48:0] inst_cellmath__200_0_out0;
input [49:0] inst_cellmath__200_0_in0;
wire N398;
CLKINVX6 inst_cellmath__200_0_I99 (.Y(N398), .A(inst_cellmath__200_0_in0[49]));
AND2XL inst_cellmath__200_0_I49 (.Y(inst_cellmath__200_0_out0[0]), .A(inst_cellmath__200_0_in0[0]), .B(N398));
AND2XL inst_cellmath__200_0_I50 (.Y(inst_cellmath__200_0_out0[1]), .A(inst_cellmath__200_0_in0[1]), .B(N398));
AND2XL inst_cellmath__200_0_I51 (.Y(inst_cellmath__200_0_out0[2]), .A(inst_cellmath__200_0_in0[2]), .B(N398));
AND2XL inst_cellmath__200_0_I52 (.Y(inst_cellmath__200_0_out0[3]), .A(inst_cellmath__200_0_in0[3]), .B(N398));
AND2XL inst_cellmath__200_0_I53 (.Y(inst_cellmath__200_0_out0[4]), .A(inst_cellmath__200_0_in0[4]), .B(N398));
AND2XL inst_cellmath__200_0_I54 (.Y(inst_cellmath__200_0_out0[5]), .A(inst_cellmath__200_0_in0[5]), .B(N398));
AND2XL inst_cellmath__200_0_I55 (.Y(inst_cellmath__200_0_out0[6]), .A(inst_cellmath__200_0_in0[6]), .B(N398));
AND2XL inst_cellmath__200_0_I56 (.Y(inst_cellmath__200_0_out0[7]), .A(inst_cellmath__200_0_in0[7]), .B(N398));
AND2XL inst_cellmath__200_0_I57 (.Y(inst_cellmath__200_0_out0[8]), .A(inst_cellmath__200_0_in0[8]), .B(N398));
AND2XL inst_cellmath__200_0_I58 (.Y(inst_cellmath__200_0_out0[9]), .A(inst_cellmath__200_0_in0[9]), .B(N398));
AND2XL inst_cellmath__200_0_I59 (.Y(inst_cellmath__200_0_out0[10]), .A(inst_cellmath__200_0_in0[10]), .B(N398));
AND2XL inst_cellmath__200_0_I60 (.Y(inst_cellmath__200_0_out0[11]), .A(inst_cellmath__200_0_in0[11]), .B(N398));
AND2XL inst_cellmath__200_0_I61 (.Y(inst_cellmath__200_0_out0[12]), .A(inst_cellmath__200_0_in0[12]), .B(N398));
AND2XL inst_cellmath__200_0_I62 (.Y(inst_cellmath__200_0_out0[13]), .A(inst_cellmath__200_0_in0[13]), .B(N398));
AND2XL inst_cellmath__200_0_I63 (.Y(inst_cellmath__200_0_out0[14]), .A(inst_cellmath__200_0_in0[14]), .B(N398));
AND2XL inst_cellmath__200_0_I64 (.Y(inst_cellmath__200_0_out0[15]), .A(inst_cellmath__200_0_in0[15]), .B(N398));
AND2XL inst_cellmath__200_0_I65 (.Y(inst_cellmath__200_0_out0[16]), .A(inst_cellmath__200_0_in0[16]), .B(N398));
AND2XL inst_cellmath__200_0_I66 (.Y(inst_cellmath__200_0_out0[17]), .A(inst_cellmath__200_0_in0[17]), .B(N398));
AND2XL inst_cellmath__200_0_I67 (.Y(inst_cellmath__200_0_out0[18]), .A(inst_cellmath__200_0_in0[18]), .B(N398));
AND2XL inst_cellmath__200_0_I68 (.Y(inst_cellmath__200_0_out0[19]), .A(inst_cellmath__200_0_in0[19]), .B(N398));
AND2XL inst_cellmath__200_0_I69 (.Y(inst_cellmath__200_0_out0[20]), .A(inst_cellmath__200_0_in0[20]), .B(N398));
AND2XL inst_cellmath__200_0_I70 (.Y(inst_cellmath__200_0_out0[21]), .A(inst_cellmath__200_0_in0[21]), .B(N398));
AND2XL inst_cellmath__200_0_I71 (.Y(inst_cellmath__200_0_out0[22]), .A(inst_cellmath__200_0_in0[22]), .B(N398));
AND2XL inst_cellmath__200_0_I72 (.Y(inst_cellmath__200_0_out0[23]), .A(inst_cellmath__200_0_in0[23]), .B(N398));
AND2XL inst_cellmath__200_0_I73 (.Y(inst_cellmath__200_0_out0[24]), .A(inst_cellmath__200_0_in0[24]), .B(N398));
AND2XL inst_cellmath__200_0_I74 (.Y(inst_cellmath__200_0_out0[25]), .A(inst_cellmath__200_0_in0[25]), .B(N398));
AND2X1 inst_cellmath__200_0_I75 (.Y(inst_cellmath__200_0_out0[26]), .A(N398), .B(inst_cellmath__200_0_in0[26]));
AND2XL inst_cellmath__200_0_I76 (.Y(inst_cellmath__200_0_out0[27]), .A(inst_cellmath__200_0_in0[27]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I77 (.Y(inst_cellmath__200_0_out0[28]), .A(inst_cellmath__200_0_in0[28]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I78 (.Y(inst_cellmath__200_0_out0[29]), .A(inst_cellmath__200_0_in0[29]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I79 (.Y(inst_cellmath__200_0_out0[30]), .A(inst_cellmath__200_0_in0[30]), .B(N398));
AND2X1 inst_cellmath__200_0_I80 (.Y(inst_cellmath__200_0_out0[31]), .A(N398), .B(inst_cellmath__200_0_in0[31]));
CLKAND2X2 inst_cellmath__200_0_I81 (.Y(inst_cellmath__200_0_out0[32]), .A(inst_cellmath__200_0_in0[32]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I82 (.Y(inst_cellmath__200_0_out0[33]), .A(inst_cellmath__200_0_in0[33]), .B(N398));
AND2X1 inst_cellmath__200_0_I83 (.Y(inst_cellmath__200_0_out0[34]), .A(N398), .B(inst_cellmath__200_0_in0[34]));
AND2X1 inst_cellmath__200_0_I84 (.Y(inst_cellmath__200_0_out0[35]), .A(N398), .B(inst_cellmath__200_0_in0[35]));
AND2X1 inst_cellmath__200_0_I85 (.Y(inst_cellmath__200_0_out0[36]), .A(N398), .B(inst_cellmath__200_0_in0[36]));
CLKAND2X2 inst_cellmath__200_0_I86 (.Y(inst_cellmath__200_0_out0[37]), .A(inst_cellmath__200_0_in0[37]), .B(N398));
AND2X4 inst_cellmath__200_0_I87 (.Y(inst_cellmath__200_0_out0[38]), .A(inst_cellmath__200_0_in0[38]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I88 (.Y(inst_cellmath__200_0_out0[39]), .A(inst_cellmath__200_0_in0[39]), .B(N398));
AND2XL inst_cellmath__200_0_I89 (.Y(inst_cellmath__200_0_out0[40]), .A(inst_cellmath__200_0_in0[40]), .B(N398));
AND2XL inst_cellmath__200_0_I90 (.Y(inst_cellmath__200_0_out0[41]), .A(inst_cellmath__200_0_in0[41]), .B(N398));
AND2X1 inst_cellmath__200_0_I91 (.Y(inst_cellmath__200_0_out0[42]), .A(N398), .B(inst_cellmath__200_0_in0[42]));
AND2X1 inst_cellmath__200_0_I92 (.Y(inst_cellmath__200_0_out0[43]), .A(N398), .B(inst_cellmath__200_0_in0[43]));
AND2X6 inst_cellmath__200_0_I93 (.Y(inst_cellmath__200_0_out0[44]), .A(inst_cellmath__200_0_in0[44]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I94 (.Y(inst_cellmath__200_0_out0[45]), .A(inst_cellmath__200_0_in0[45]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I95 (.Y(inst_cellmath__200_0_out0[46]), .A(inst_cellmath__200_0_in0[46]), .B(N398));
CLKAND2X2 inst_cellmath__200_0_I96 (.Y(inst_cellmath__200_0_out0[47]), .A(inst_cellmath__200_0_in0[47]), .B(N398));
AND2XL inst_cellmath__200_0_I97 (.Y(inst_cellmath__200_0_out0[48]), .A(inst_cellmath__200_0_in0[48]), .B(N398));
endmodule

module cynw_cm_float_cos_inst_cellmath__17_0_bdw1157874770_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NOR2X1 inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[0]));
NOR2X1 inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[6]), .B(inst_cellmath__17_0_in0[5]));
NOR2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[4]), .B(inst_cellmath__17_0_in0[3]));
NOR2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[2]), .B(inst_cellmath__17_0_in0[1]));
NAND2X1 inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_cos_inst_cellmath__46__15__bdw1157874770_bdw (
	inst_cellmath__46__15__out0,
	inst_cellmath__46__15__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__46__15__out0;
input [7:6] inst_cellmath__46__15__in0;
OR2XL inst_cellmath__46__15__I0 (.Y(inst_cellmath__46__15__out0[0]), .A(inst_cellmath__46__15__in0[7]), .B(inst_cellmath__46__15__in0[6]));
endmodule

module cynw_cm_float_cos_inst_cellmath__46_0_bdw1157874770_bdw (
	inst_cellmath__46_0_out0,
	inst_cellmath__46_0_in0,
	inst_cellmath__46_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__46_0_out0;
input [0:0] inst_cellmath__46_0_in0;
input [8:8] inst_cellmath__46_0_in1;
wire N5;
INVXL inst_cellmath__46_0_I0 (.Y(N5), .A(inst_cellmath__46_0_in1[8]));
AND2XL inst_cellmath__46_0_I1 (.Y(inst_cellmath__46_0_out0), .A(N5), .B(inst_cellmath__46_0_in0[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__21_0_bdw1157874770_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__21_0_out0;
input [7:0] inst_cellmath__21_0_in0;
wire N62,N64,N68,N70;
NAND2X1 inst_cellmath__21_0_I29 (.Y(N62), .A(inst_cellmath__21_0_in0[2]), .B(inst_cellmath__21_0_in0[1]));
NOR2XL inst_cellmath__21_0_I30 (.Y(N64), .A(inst_cellmath__21_0_in0[3]), .B(inst_cellmath__21_0_in0[4]));
NAND2X1 inst_cellmath__21_0_I32 (.Y(N68), .A(inst_cellmath__21_0_in0[5]), .B(inst_cellmath__21_0_in0[6]));
AOI21X1 inst_cellmath__21_0_I37 (.Y(N70), .A0(N62), .A1(N64), .B0(N68));
NOR2X1 inst_cellmath__21_0_I34 (.Y(inst_cellmath__21_0_out0), .A(inst_cellmath__21_0_in0[7]), .B(N70));
endmodule

module cynw_cm_float_cos_inst_cellmath__83__62__bdw1157874770_bdw (
	inst_cellmath__83__62__out0,
	inst_cellmath__83__62__in0,
	inst_cellmath__83__62__in1,
	inst_cellmath__83__62__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__83__62__out0;
input  inst_cellmath__83__62__in0,
	inst_cellmath__83__62__in1,
	inst_cellmath__83__62__in2;
wire N7,N25;
OR2XL inst_cellmath__83__62__I0 (.Y(N7), .A(inst_cellmath__83__62__in2), .B(inst_cellmath__83__62__in1));
NOR2X2 or2_A_I10 (.Y(N25), .A(N7), .B(inst_cellmath__83__62__in0));
INVXL or2_A_I11 (.Y(inst_cellmath__83__62__out0[0]), .A(N25));
endmodule

module cynw_cm_float_cos_inst_cellmath__19_0_bdw1157874770_bdw (
	inst_cellmath__19_0_out0,
	inst_cellmath__19_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19_0_out0;
input [7:0] inst_cellmath__19_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2X1 inst_cellmath__19_0_I0 (.Y(N11), .A(inst_cellmath__19_0_in0[7]), .B(inst_cellmath__19_0_in0[0]));
NAND2XL inst_cellmath__19_0_I1 (.Y(N12), .A(inst_cellmath__19_0_in0[6]), .B(inst_cellmath__19_0_in0[5]));
NAND2X1 inst_cellmath__19_0_I2 (.Y(N13), .A(inst_cellmath__19_0_in0[4]), .B(inst_cellmath__19_0_in0[3]));
NAND2XL inst_cellmath__19_0_I3 (.Y(N14), .A(inst_cellmath__19_0_in0[2]), .B(inst_cellmath__19_0_in0[1]));
NOR2XL inst_cellmath__19_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__19_0_I5 (.Y(N16), .A(N13), .B(N14));
CLKAND2X2 inst_cellmath__19_0_I6 (.Y(inst_cellmath__19_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_cos_inst_cellmath__24_0_bdw1157874770_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__24_0_out0;
input [22:0] inst_cellmath__24_0_in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N37,N38,N39,N40 
	,N41,N42,N43,N44,N45,N47,N48;
NOR2XL inst_cellmath__24_0_I0 (.Y(N26), .A(inst_cellmath__24_0_in0[0]), .B(inst_cellmath__24_0_in0[1]));
NOR2XL inst_cellmath__24_0_I1 (.Y(N27), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
NOR2XL inst_cellmath__24_0_I2 (.Y(N28), .A(inst_cellmath__24_0_in0[20]), .B(inst_cellmath__24_0_in0[19]));
NOR2XL inst_cellmath__24_0_I3 (.Y(N29), .A(inst_cellmath__24_0_in0[18]), .B(inst_cellmath__24_0_in0[17]));
NOR2XL inst_cellmath__24_0_I4 (.Y(N30), .A(inst_cellmath__24_0_in0[16]), .B(inst_cellmath__24_0_in0[15]));
NOR2XL inst_cellmath__24_0_I5 (.Y(N31), .A(inst_cellmath__24_0_in0[14]), .B(inst_cellmath__24_0_in0[13]));
NOR2XL inst_cellmath__24_0_I6 (.Y(N32), .A(inst_cellmath__24_0_in0[12]), .B(inst_cellmath__24_0_in0[11]));
NOR2XL inst_cellmath__24_0_I7 (.Y(N33), .A(inst_cellmath__24_0_in0[10]), .B(inst_cellmath__24_0_in0[9]));
NOR2X6 inst_cellmath__24_0_I8 (.Y(N34), .A(inst_cellmath__24_0_in0[8]), .B(inst_cellmath__24_0_in0[7]));
NOR2XL inst_cellmath__24_0_I9 (.Y(N35), .A(inst_cellmath__24_0_in0[6]), .B(inst_cellmath__24_0_in0[5]));
NOR2XL inst_cellmath__24_0_I10 (.Y(N36), .A(inst_cellmath__24_0_in0[4]), .B(inst_cellmath__24_0_in0[3]));
INVXL inst_cellmath__24_0_I11 (.Y(N37), .A(inst_cellmath__24_0_in0[2]));
NAND2XL inst_cellmath__24_0_I12 (.Y(N38), .A(N37), .B(N26));
NAND2XL inst_cellmath__24_0_I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__24_0_I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__24_0_I15 (.Y(N41), .A(N31), .B(N32));
NAND2XL inst_cellmath__24_0_I16 (.Y(N42), .A(N33), .B(N34));
NAND2XL inst_cellmath__24_0_I17 (.Y(N43), .A(N35), .B(N36));
NOR2XL inst_cellmath__24_0_I18 (.Y(N44), .A(N38), .B(N39));
NOR2XL inst_cellmath__24_0_I19 (.Y(N45), .A(N40), .B(N41));
NAND2XL inst_cellmath__24_0_I21 (.Y(N47), .A(N44), .B(N45));
OR2XL inst_cellmath__24_0_I169 (.Y(N48), .A(N42), .B(N43));
NOR2XL inst_cellmath__24_0_I23 (.Y(inst_cellmath__24_0_out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_cos_inst_cellmath__69_0_bdw1157874770_bdw (
	inst_cellmath__69_0_out0,
	inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__69_0_out0;
input  inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1;
wire N5;
INVXL inst_cellmath__69_0_I0 (.Y(N5), .A(inst_cellmath__69_0_in1));
NOR2X2 inst_cellmath__69_0_I1 (.Y(inst_cellmath__69_0_out0), .A(N5), .B(inst_cellmath__69_0_in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__82_0_bdw1157874770_bdw (
	inst_cellmath__82_0_out0,
	inst_cellmath__82_0_in0,
	inst_cellmath__82_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__82_0_out0;
input  inst_cellmath__82_0_in0,
	inst_cellmath__82_0_in1;
wire N19;
NOR2X1 inst_cellmath__82_0_I4 (.Y(N19), .A(inst_cellmath__82_0_in1), .B(inst_cellmath__82_0_in0));
INVX1 inst_cellmath__82_0_I5 (.Y(inst_cellmath__82_0_out0), .A(N19));
endmodule

module cynw_cm_float_cos_inst_cellmath__66_0_bdw1157874770_bdw (
	inst_cellmath__66_0_out0,
	inst_cellmath__66_0_in0,
	inst_cellmath__66_0_in1,
	inst_cellmath__66_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__66_0_out0;
input  inst_cellmath__66_0_in0,
	inst_cellmath__66_0_in1,
	inst_cellmath__66_0_in2;
wire N6,N8;
INVXL inst_cellmath__66_0_I0 (.Y(N6), .A(inst_cellmath__66_0_in2));
CLKAND2X3 inst_cellmath__66_0_I1 (.Y(N8), .A(N6), .B(inst_cellmath__66_0_in1));
CLKAND2X3 inst_cellmath__66_0_I3 (.Y(inst_cellmath__66_0_out0), .A(N8), .B(inst_cellmath__66_0_in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__67_0_bdw1157874770_bdw (
	inst_cellmath__67_0_out0,
	inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1,
	inst_cellmath__67_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__67_0_out0;
input  inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1,
	inst_cellmath__67_0_in2;
wire N7;
CLKAND2X3 inst_cellmath__67_0_I0 (.Y(N7), .A(inst_cellmath__67_0_in2), .B(inst_cellmath__67_0_in1));
CLKAND2X3 inst_cellmath__67_0_I2 (.Y(inst_cellmath__67_0_out0), .A(N7), .B(inst_cellmath__67_0_in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__68_0_bdw1157874770_bdw (
	inst_cellmath__68_0_out0,
	inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__68_0_out0;
input  inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1;
OR2XL inst_cellmath__68_0_I0 (.Y(inst_cellmath__68_0_out0), .A(inst_cellmath__68_0_in0), .B(inst_cellmath__68_0_in1));
endmodule

module cynw_cm_float_cos_inst_cellmath__228__231__bdw1157874770_bdw (
	inst_cellmath__228__231__out0,
	inst_cellmath__228__231__in0,
	inst_cellmath__228__231__in1,
	inst_cellmath__228__231__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__228__231__out0;
input [0:0] inst_cellmath__228__231__in0;
input  inst_cellmath__228__231__in1,
	inst_cellmath__228__231__in2;
wire N7,N25;
OR2XL inst_cellmath__228__231__I0 (.Y(N7), .A(inst_cellmath__228__231__in1), .B(inst_cellmath__228__231__in2));
NOR2X2 or2_A_I10 (.Y(N25), .A(N7), .B(inst_cellmath__228__231__in0[0]));
INVX1 or2_A_I11 (.Y(inst_cellmath__228__231__out0[0]), .A(N25));
endmodule

module cynw_cm_float_cos_inst_cellmath__219_0_bdw1157874770_bdw (
	inst_cellmath__219_0_out0,
	inst_cellmath__219_0_in0,
	inst_cellmath__219_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__219_0_out0;
input [22:22] inst_cellmath__219_0_in0;
input [48:48] inst_cellmath__219_0_in1;
AND2XL inst_cellmath__219_0_I0 (.Y(inst_cellmath__219_0_out0), .A(inst_cellmath__219_0_in0[22]), .B(inst_cellmath__219_0_in1[48]));
endmodule

module cynw_cm_float_cos_inst_cellmath__211__182__bdw1157874770_bdw (
	inst_cellmath__211__182__out0,
	inst_cellmath__211__182__in0
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__211__182__out0;
input [47:25] inst_cellmath__211__182__in0;
wire N100,N106,N108,N109,N112,N113,N114 
	,N115,N116,N117,N118,N119,N120,N121,N122 
	,N123,N124,N125,N126,N127,N128,N129,N131 
	,N132,N133,N134,N135,N137,N139,N140,N141 
	,N155,N157,N158,N160,N162,N163,N164,N165 
	,N166,N168,N169,N170,N171,N172,N180,N182 
	,N183,N185,N189,N191,N216,N218,N232,N234 
	,N240,N242,N248;
INVXL inst_cellmath__211__182__I7 (.Y(N100), .A(inst_cellmath__211__182__in0[47]));
INVX2 inst_cellmath__211__182__I11 (.Y(N106), .A(inst_cellmath__211__182__in0[25]));
INVX1 inst_cellmath__211__182__I12 (.Y(N108), .A(inst_cellmath__211__182__in0[27]));
OAI21X4 inst_cellmath__211__182__I13 (.Y(N109), .A0(inst_cellmath__211__182__in0[26]), .A1(N106), .B0(N108));
INVX2 inst_cellmath__211__182__I16 (.Y(N112), .A(inst_cellmath__211__182__in0[28]));
NOR2X4 inst_cellmath__211__182__I17 (.Y(N113), .A(inst_cellmath__211__182__in0[29]), .B(N112));
INVX1 inst_cellmath__211__182__I18 (.Y(N114), .A(inst_cellmath__211__182__in0[31]));
OAI21X4 inst_cellmath__211__182__I19 (.Y(N115), .A0(inst_cellmath__211__182__in0[30]), .A1(N113), .B0(N114));
NOR2X2 inst_cellmath__211__182__I20 (.Y(N116), .A(inst_cellmath__211__182__in0[29]), .B(inst_cellmath__211__182__in0[28]));
NOR2X2 inst_cellmath__211__182__I21 (.Y(N117), .A(inst_cellmath__211__182__in0[31]), .B(inst_cellmath__211__182__in0[30]));
INVXL inst_cellmath__211__182__I22 (.Y(N118), .A(inst_cellmath__211__182__in0[32]));
NOR2X1 inst_cellmath__211__182__I23 (.Y(N119), .A(inst_cellmath__211__182__in0[33]), .B(N118));
INVXL inst_cellmath__211__182__I24 (.Y(N120), .A(inst_cellmath__211__182__in0[35]));
OAI21X2 inst_cellmath__211__182__I25 (.Y(N121), .A0(inst_cellmath__211__182__in0[34]), .A1(N119), .B0(N120));
NOR2X2 inst_cellmath__211__182__I26 (.Y(N122), .A(inst_cellmath__211__182__in0[33]), .B(inst_cellmath__211__182__in0[32]));
NOR2X2 inst_cellmath__211__182__I27 (.Y(N123), .A(inst_cellmath__211__182__in0[35]), .B(inst_cellmath__211__182__in0[34]));
INVX1 inst_cellmath__211__182__I28 (.Y(N124), .A(inst_cellmath__211__182__in0[36]));
NOR2X1 inst_cellmath__211__182__I29 (.Y(N125), .A(inst_cellmath__211__182__in0[37]), .B(N124));
INVXL inst_cellmath__211__182__I30 (.Y(N126), .A(inst_cellmath__211__182__in0[39]));
OAI21X2 inst_cellmath__211__182__I31 (.Y(N127), .A0(inst_cellmath__211__182__in0[38]), .A1(N125), .B0(N126));
NOR2X2 inst_cellmath__211__182__I32 (.Y(N128), .A(inst_cellmath__211__182__in0[37]), .B(inst_cellmath__211__182__in0[36]));
NOR2X4 inst_cellmath__211__182__I33 (.Y(N129), .A(inst_cellmath__211__182__in0[39]), .B(inst_cellmath__211__182__in0[38]));
NOR2BX1 inst_cellmath__211__182__I576 (.Y(N131), .AN(inst_cellmath__211__182__in0[40]), .B(inst_cellmath__211__182__in0[41]));
INVXL inst_cellmath__211__182__I36 (.Y(N132), .A(inst_cellmath__211__182__in0[43]));
OAI21X2 inst_cellmath__211__182__I37 (.Y(N133), .A0(inst_cellmath__211__182__in0[42]), .A1(N131), .B0(N132));
NOR2XL inst_cellmath__211__182__I38 (.Y(N134), .A(inst_cellmath__211__182__in0[41]), .B(inst_cellmath__211__182__in0[40]));
NOR2X2 inst_cellmath__211__182__I39 (.Y(N135), .A(inst_cellmath__211__182__in0[43]), .B(inst_cellmath__211__182__in0[42]));
NOR2BX1 inst_cellmath__211__182__I577 (.Y(N137), .AN(inst_cellmath__211__182__in0[44]), .B(inst_cellmath__211__182__in0[45]));
OAI21X1 inst_cellmath__211__182__I43 (.Y(N139), .A0(inst_cellmath__211__182__in0[46]), .A1(N137), .B0(N100));
NOR2X2 inst_cellmath__211__182__I44 (.Y(N140), .A(inst_cellmath__211__182__in0[45]), .B(inst_cellmath__211__182__in0[44]));
NOR2X2 inst_cellmath__211__182__I45 (.Y(N141), .A(inst_cellmath__211__182__in0[47]), .B(inst_cellmath__211__182__in0[46]));
OR2XL inst_cellmath__211__182__I578 (.Y(N155), .A(inst_cellmath__211__182__in0[27]), .B(inst_cellmath__211__182__in0[26]));
INVXL inst_cellmath__211__182__I60 (.Y(N157), .A(N117));
AOI21XL inst_cellmath__211__182__I61 (.Y(N158), .A0(N116), .A1(N155), .B0(N157));
NAND2X2 inst_cellmath__211__182__I63 (.Y(N160), .A(N117), .B(N116));
NAND2BXL inst_cellmath__211__182__I579 (.Y(N162), .AN(N122), .B(N123));
INVXL inst_cellmath__211__182__I66 (.Y(N163), .A(N129));
AOI21XL inst_cellmath__211__182__I67 (.Y(N164), .A0(N128), .A1(N162), .B0(N163));
NAND2X2 inst_cellmath__211__182__I68 (.Y(N165), .A(N123), .B(N122));
NAND2X4 inst_cellmath__211__182__I69 (.Y(N166), .A(N129), .B(N128));
NAND2BXL inst_cellmath__211__182__I580 (.Y(N168), .AN(N134), .B(N135));
INVXL inst_cellmath__211__182__I72 (.Y(N169), .A(N141));
AOI21XL inst_cellmath__211__182__I73 (.Y(N170), .A0(N140), .A1(N168), .B0(N169));
NAND2X1 inst_cellmath__211__182__I74 (.Y(N171), .A(N135), .B(N134));
NAND2X2 inst_cellmath__211__182__I75 (.Y(N172), .A(N141), .B(N140));
INVXL inst_cellmath__211__182__I83 (.Y(N180), .A(N160));
INVXL inst_cellmath__211__182__I84 (.Y(N182), .A(N166));
OAI21XL inst_cellmath__211__182__I85 (.Y(N183), .A0(N165), .A1(N180), .B0(N182));
NOR2X4 inst_cellmath__211__182__I87 (.Y(N185), .A(N166), .B(N165));
NAND2BXL inst_cellmath__211__182__I582 (.Y(N189), .AN(N172), .B(N171));
NOR2X2 inst_cellmath__211__182__I92 (.Y(N191), .A(N172), .B(N171));
NAND2BXL inst_cellmath__211__182__I583 (.Y(inst_cellmath__211__182__out0[3]), .AN(N185), .B(N191));
INVX2 inst_cellmath__211__182__I140 (.Y(N248), .A(N191));
INVXL inst_cellmath__211__182__I101 (.Y(inst_cellmath__211__182__out0[4]), .A(N248));
OAI21XL inst_cellmath__211__182__I106 (.Y(inst_cellmath__211__182__out0[2]), .A0(N248), .A1(N183), .B0(N189));
AOI21XL inst_cellmath__211__182__I112 (.Y(N216), .A0(N185), .A1(N158), .B0(N164));
INVXL inst_cellmath__211__182__I114 (.Y(N218), .A(N170));
OAI21X1 inst_cellmath__211__182__I116 (.Y(inst_cellmath__211__182__out0[1]), .A0(N248), .A1(N216), .B0(N218));
OAI21X2 inst_cellmath__211__182__I126 (.Y(N232), .A0(N160), .A1(N109), .B0(N115));
OAI21X2 inst_cellmath__211__182__I128 (.Y(N234), .A0(N166), .A1(N121), .B0(N127));
AOI21X2 inst_cellmath__211__182__I134 (.Y(N240), .A0(N185), .A1(N232), .B0(N234));
OA21X1 inst_cellmath__211__182__I584 (.Y(N242), .A0(N172), .A1(N133), .B0(N139));
OAI21X2 inst_cellmath__211__182__I138 (.Y(inst_cellmath__211__182__out0[0]), .A0(N248), .A1(N240), .B0(N242));
endmodule

module cynw_cm_float_cos_inst_cellmath__215_0_bdw1157874770_bdw (
	inst_cellmath__215_0_out0,
	inst_cellmath__215_0_in0
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__215_0_out0;
input [4:0] inst_cellmath__215_0_in0;
wire N47,N67,N72,N145,N155,N168;
INVXL inst_cellmath__215_0_I81 (.Y(N155), .A(inst_cellmath__215_0_in0[0]));
AND2XL inst_cellmath__215_0_I21 (.Y(N47), .A(inst_cellmath__215_0_in0[1]), .B(inst_cellmath__215_0_in0[0]));
NAND2XL hyperpropagate_3_1_A_I102 (.Y(N168), .A(inst_cellmath__215_0_in0[2]), .B(inst_cellmath__215_0_in0[1]));
NOR2XL hyperpropagate_3_1_A_I103 (.Y(N67), .A(N155), .B(N168));
AO21XL inst_cellmath__215_0_I35 (.Y(N72), .A0(inst_cellmath__215_0_in0[2]), .A1(N47), .B0(inst_cellmath__215_0_in0[3]));
INVXL inst_cellmath__215_0_I64 (.Y(inst_cellmath__215_0_out0[0]), .A(inst_cellmath__215_0_in0[0]));
XNOR2X1 inst_cellmath__215_0_I98 (.Y(inst_cellmath__215_0_out0[1]), .A(N155), .B(inst_cellmath__215_0_in0[1]));
XOR2XL inst_cellmath__215_0_I96 (.Y(inst_cellmath__215_0_out0[2]), .A(N47), .B(inst_cellmath__215_0_in0[2]));
XNOR2X1 inst_cellmath__215_0_I67 (.Y(inst_cellmath__215_0_out0[3]), .A(N67), .B(inst_cellmath__215_0_in0[3]));
INVXL xnor2_A_I75 (.Y(N145), .A(N72));
MXI2XL xnor2_A_I76 (.Y(inst_cellmath__215_0_out0[4]), .A(N72), .B(N145), .S0(inst_cellmath__215_0_in0[4]));
endmodule

module cynw_cm_float_cos_inst_cellmath__220__188__bdw1157874770_bdw (
	inst_cellmath__220__188__out0,
	inst_cellmath__220__188__in0,
	inst_cellmath__220__188__in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__220__188__out0;
input [4:0] inst_cellmath__220__188__in0;
input [47:25] inst_cellmath__220__188__in1;
wire N55,N57,N58,N59,N60,N61,N62 
	,N63,N64,N65,N66,N67,N68,N69,N70 
	,N71,N72,N73,N74,N75,N76,N77,N78 
	,N106,N108,N110,N111,N112,N113,N114,N115 
	,N116,N117,N118,N119,N120,N121,N122,N123 
	,N124,N125,N126,N127,N128,N129,N130,N158 
	,N160,N162,N164,N166,N168,N170,N172,N174 
	,N175,N176,N177,N178,N179,N180,N181,N182 
	,N183,N184,N185,N186,N187,N188,N216,N218 
	,N220,N222,N224,N226,N228,N230,N232,N234 
	,N236,N238,N240,N242,N244,N246,N248,N249 
	,N250,N251,N252,N253,N254,N335,N340,N341 
	,N342,N343,N345,N346,N347,N348,N349,N350 
	,N351,N352,N353,N355,N357,N358,N360,N364 
	;
BUFX2 inst_cellmath__220__188__I281 (.Y(N335), .A(inst_cellmath__220__188__in0[0]));
INVXL inst_cellmath__220__188__I257 (.Y(N341), .A(N335));
INVX2 inst_cellmath__220__188__I256 (.Y(N340), .A(N335));
AND2XL inst_cellmath__220__188__I2 (.Y(N55), .A(N341), .B(inst_cellmath__220__188__in1[25]));
MX2XL inst_cellmath__220__188__I3 (.Y(N57), .A(inst_cellmath__220__188__in1[25]), .B(inst_cellmath__220__188__in1[26]), .S0(N341));
MX2XL inst_cellmath__220__188__I4 (.Y(N58), .A(inst_cellmath__220__188__in1[26]), .B(inst_cellmath__220__188__in1[27]), .S0(N341));
MX2XL inst_cellmath__220__188__I5 (.Y(N59), .A(inst_cellmath__220__188__in1[27]), .B(inst_cellmath__220__188__in1[28]), .S0(N340));
MX2XL inst_cellmath__220__188__I6 (.Y(N60), .A(inst_cellmath__220__188__in1[28]), .B(inst_cellmath__220__188__in1[29]), .S0(N340));
MX2XL inst_cellmath__220__188__I7 (.Y(N61), .A(inst_cellmath__220__188__in1[29]), .B(inst_cellmath__220__188__in1[30]), .S0(N340));
MX2XL inst_cellmath__220__188__I8 (.Y(N62), .A(inst_cellmath__220__188__in1[30]), .B(inst_cellmath__220__188__in1[31]), .S0(N340));
MX2XL inst_cellmath__220__188__I9 (.Y(N63), .A(inst_cellmath__220__188__in1[31]), .B(inst_cellmath__220__188__in1[32]), .S0(N340));
MX2XL inst_cellmath__220__188__I10 (.Y(N64), .A(inst_cellmath__220__188__in1[32]), .B(inst_cellmath__220__188__in1[33]), .S0(N340));
MX2XL inst_cellmath__220__188__I11 (.Y(N65), .A(inst_cellmath__220__188__in1[33]), .B(inst_cellmath__220__188__in1[34]), .S0(N340));
MX2XL inst_cellmath__220__188__I12 (.Y(N66), .A(inst_cellmath__220__188__in1[34]), .B(inst_cellmath__220__188__in1[35]), .S0(N340));
MX2XL inst_cellmath__220__188__I13 (.Y(N67), .A(inst_cellmath__220__188__in1[35]), .B(inst_cellmath__220__188__in1[36]), .S0(N340));
MX2XL inst_cellmath__220__188__I14 (.Y(N68), .A(inst_cellmath__220__188__in1[36]), .B(inst_cellmath__220__188__in1[37]), .S0(N340));
MX2XL inst_cellmath__220__188__I15 (.Y(N69), .A(inst_cellmath__220__188__in1[37]), .B(inst_cellmath__220__188__in1[38]), .S0(N340));
MX2XL inst_cellmath__220__188__I16 (.Y(N70), .A(inst_cellmath__220__188__in1[38]), .B(inst_cellmath__220__188__in1[39]), .S0(N340));
MX2XL inst_cellmath__220__188__I17 (.Y(N71), .A(inst_cellmath__220__188__in1[39]), .B(inst_cellmath__220__188__in1[40]), .S0(N340));
MX2XL inst_cellmath__220__188__I18 (.Y(N72), .A(inst_cellmath__220__188__in1[40]), .B(inst_cellmath__220__188__in1[41]), .S0(N340));
MX2XL inst_cellmath__220__188__I19 (.Y(N73), .A(inst_cellmath__220__188__in1[41]), .B(inst_cellmath__220__188__in1[42]), .S0(N340));
MX2XL inst_cellmath__220__188__I20 (.Y(N74), .A(inst_cellmath__220__188__in1[42]), .B(inst_cellmath__220__188__in1[43]), .S0(N340));
MX2XL inst_cellmath__220__188__I21 (.Y(N75), .A(inst_cellmath__220__188__in1[43]), .B(inst_cellmath__220__188__in1[44]), .S0(N341));
MX2XL inst_cellmath__220__188__I22 (.Y(N76), .A(inst_cellmath__220__188__in1[44]), .B(inst_cellmath__220__188__in1[45]), .S0(N341));
MX2XL inst_cellmath__220__188__I23 (.Y(N77), .A(inst_cellmath__220__188__in1[45]), .B(inst_cellmath__220__188__in1[46]), .S0(N341));
MX2XL inst_cellmath__220__188__I24 (.Y(N78), .A(inst_cellmath__220__188__in1[46]), .B(inst_cellmath__220__188__in1[47]), .S0(N341));
CLKINVX6 inst_cellmath__220__188__I258 (.Y(N342), .A(inst_cellmath__220__188__in0[1]));
NAND2XL inst_cellmath__220__188__I52 (.Y(N106), .A(N55), .B(N342));
NAND2XL inst_cellmath__220__188__I53 (.Y(N108), .A(N57), .B(N342));
MXI2XL inst_cellmath__220__188__I54 (.Y(N110), .A(N55), .B(N58), .S0(N342));
MXI2XL inst_cellmath__220__188__I55 (.Y(N111), .A(N57), .B(N59), .S0(N342));
MXI2XL inst_cellmath__220__188__I56 (.Y(N112), .A(N58), .B(N60), .S0(N342));
MXI2XL inst_cellmath__220__188__I57 (.Y(N113), .A(N59), .B(N61), .S0(N342));
MXI2XL inst_cellmath__220__188__I58 (.Y(N114), .A(N60), .B(N62), .S0(N342));
MXI2XL inst_cellmath__220__188__I59 (.Y(N115), .A(N61), .B(N63), .S0(N342));
MXI2X1 inst_cellmath__220__188__I60 (.Y(N116), .A(N62), .B(N64), .S0(N342));
MXI2XL inst_cellmath__220__188__I61 (.Y(N117), .A(N63), .B(N65), .S0(N342));
MXI2XL inst_cellmath__220__188__I62 (.Y(N118), .A(N64), .B(N66), .S0(N342));
MXI2XL inst_cellmath__220__188__I63 (.Y(N119), .A(N65), .B(N67), .S0(N342));
MXI2XL inst_cellmath__220__188__I64 (.Y(N120), .A(N66), .B(N68), .S0(N342));
MXI2XL inst_cellmath__220__188__I65 (.Y(N121), .A(N67), .B(N69), .S0(N342));
MXI2XL inst_cellmath__220__188__I66 (.Y(N122), .A(N68), .B(N70), .S0(N342));
MXI2XL inst_cellmath__220__188__I67 (.Y(N123), .A(N69), .B(N71), .S0(N342));
MXI2XL inst_cellmath__220__188__I68 (.Y(N124), .A(N70), .B(N72), .S0(N342));
MXI2XL inst_cellmath__220__188__I69 (.Y(N125), .A(N71), .B(N73), .S0(N342));
MXI2XL inst_cellmath__220__188__I70 (.Y(N126), .A(N72), .B(N74), .S0(N342));
MXI2XL inst_cellmath__220__188__I71 (.Y(N127), .A(N73), .B(N75), .S0(N342));
MXI2X2 inst_cellmath__220__188__I72 (.Y(N128), .A(N74), .B(N76), .S0(N342));
MXI2X2 inst_cellmath__220__188__I73 (.Y(N129), .A(N75), .B(N77), .S0(N342));
MXI2X2 inst_cellmath__220__188__I74 (.Y(N130), .A(N76), .B(N78), .S0(N342));
INVX3 inst_cellmath__220__188__I259 (.Y(N343), .A(inst_cellmath__220__188__in0[3]));
INVXL inst_cellmath__220__188__I265 (.Y(N349), .A(N343));
INVXL inst_cellmath__220__188__I264 (.Y(N348), .A(N343));
INVXL inst_cellmath__220__188__I263 (.Y(N347), .A(N343));
INVXL inst_cellmath__220__188__I262 (.Y(N346), .A(N343));
INVX1 inst_cellmath__220__188__I261 (.Y(N345), .A(N343));
NOR2XL inst_cellmath__220__188__I102 (.Y(N158), .A(N106), .B(N349));
NOR2XL inst_cellmath__220__188__I103 (.Y(N160), .A(N108), .B(N349));
NOR2XL inst_cellmath__220__188__I104 (.Y(N162), .A(N110), .B(N349));
NOR2XL inst_cellmath__220__188__I105 (.Y(N164), .A(N111), .B(N348));
NOR2XL inst_cellmath__220__188__I106 (.Y(N166), .A(N112), .B(N348));
NOR2XL inst_cellmath__220__188__I107 (.Y(N168), .A(N113), .B(N348));
NOR2XL inst_cellmath__220__188__I108 (.Y(N170), .A(N114), .B(N348));
NOR2XL inst_cellmath__220__188__I109 (.Y(N172), .A(N115), .B(N347));
MXI2XL inst_cellmath__220__188__I110 (.Y(N174), .A(N116), .B(N106), .S0(N347));
MXI2XL inst_cellmath__220__188__I111 (.Y(N175), .A(N117), .B(N108), .S0(N347));
MXI2XL inst_cellmath__220__188__I112 (.Y(N176), .A(N118), .B(N110), .S0(N347));
MXI2XL inst_cellmath__220__188__I113 (.Y(N177), .A(N119), .B(N111), .S0(N346));
MXI2XL inst_cellmath__220__188__I114 (.Y(N178), .A(N120), .B(N112), .S0(N346));
MXI2XL inst_cellmath__220__188__I115 (.Y(N179), .A(N121), .B(N113), .S0(N346));
MXI2XL inst_cellmath__220__188__I116 (.Y(N180), .A(N122), .B(N114), .S0(N346));
MXI2XL inst_cellmath__220__188__I117 (.Y(N181), .A(N123), .B(N115), .S0(N345));
MXI2X1 inst_cellmath__220__188__I118 (.Y(N182), .A(N124), .B(N116), .S0(N345));
MXI2XL inst_cellmath__220__188__I119 (.Y(N183), .A(N125), .B(N117), .S0(N345));
MXI2XL inst_cellmath__220__188__I120 (.Y(N184), .A(N126), .B(N118), .S0(N345));
MXI2XL inst_cellmath__220__188__I121 (.Y(N185), .A(N127), .B(N119), .S0(N348));
MXI2XL inst_cellmath__220__188__I122 (.Y(N186), .A(N128), .B(N120), .S0(N348));
MXI2XL inst_cellmath__220__188__I123 (.Y(N187), .A(N129), .B(N121), .S0(N348));
MXI2XL inst_cellmath__220__188__I124 (.Y(N188), .A(N130), .B(N122), .S0(N348));
INVX1 inst_cellmath__220__188__I266 (.Y(N350), .A(inst_cellmath__220__188__in0[4]));
INVX2 inst_cellmath__220__188__I267 (.Y(N351), .A(N350));
INVX2 inst_cellmath__220__188__I273 (.Y(N357), .A(N351));
INVXL inst_cellmath__220__188__I271 (.Y(N355), .A(N351));
INVXL inst_cellmath__220__188__I269 (.Y(N353), .A(N351));
INVXL inst_cellmath__220__188__I268 (.Y(N352), .A(N351));
NAND2XL inst_cellmath__220__188__I152 (.Y(N216), .A(N158), .B(N357));
NAND2XL inst_cellmath__220__188__I153 (.Y(N218), .A(N160), .B(N357));
NAND2XL inst_cellmath__220__188__I154 (.Y(N220), .A(N162), .B(N357));
NAND2XL inst_cellmath__220__188__I155 (.Y(N222), .A(N164), .B(N357));
NAND2XL inst_cellmath__220__188__I156 (.Y(N224), .A(N166), .B(N357));
NAND2XL inst_cellmath__220__188__I157 (.Y(N226), .A(N168), .B(N357));
NAND2XL inst_cellmath__220__188__I158 (.Y(N228), .A(N170), .B(N357));
NAND2XL inst_cellmath__220__188__I159 (.Y(N230), .A(N172), .B(N355));
NAND2XL inst_cellmath__220__188__I160 (.Y(N232), .A(N174), .B(N355));
NAND2XL inst_cellmath__220__188__I161 (.Y(N234), .A(N175), .B(N355));
NAND2XL inst_cellmath__220__188__I162 (.Y(N236), .A(N176), .B(N355));
NAND2XL inst_cellmath__220__188__I163 (.Y(N238), .A(N177), .B(N355));
NAND2XL inst_cellmath__220__188__I164 (.Y(N240), .A(N178), .B(N355));
NAND2XL inst_cellmath__220__188__I165 (.Y(N242), .A(N179), .B(N355));
NAND2XL inst_cellmath__220__188__I166 (.Y(N244), .A(N180), .B(N355));
NAND2XL inst_cellmath__220__188__I167 (.Y(N246), .A(N181), .B(N353));
MXI2X1 inst_cellmath__220__188__I168 (.Y(N248), .A(N158), .B(N182), .S0(N353));
MXI2XL inst_cellmath__220__188__I169 (.Y(N249), .A(N160), .B(N183), .S0(N353));
MXI2XL inst_cellmath__220__188__I170 (.Y(N250), .A(N162), .B(N184), .S0(N353));
MXI2XL inst_cellmath__220__188__I171 (.Y(N251), .A(N164), .B(N185), .S0(N352));
MXI2XL inst_cellmath__220__188__I172 (.Y(N252), .A(N166), .B(N186), .S0(N352));
MXI2XL inst_cellmath__220__188__I173 (.Y(N253), .A(N168), .B(N187), .S0(N352));
MXI2XL inst_cellmath__220__188__I174 (.Y(N254), .A(N170), .B(N188), .S0(N352));
INVX3 inst_cellmath__220__188__I274 (.Y(N358), .A(inst_cellmath__220__188__in0[2]));
INVX2 inst_cellmath__220__188__I280 (.Y(N364), .A(N358));
INVXL inst_cellmath__220__188__I276 (.Y(N360), .A(N358));
NOR2XL inst_cellmath__220__188__I202 (.Y(inst_cellmath__220__188__out0[0]), .A(N216), .B(N364));
NOR2XL inst_cellmath__220__188__I203 (.Y(inst_cellmath__220__188__out0[1]), .A(N218), .B(N364));
NOR2XL inst_cellmath__220__188__I204 (.Y(inst_cellmath__220__188__out0[2]), .A(N220), .B(N364));
NOR2XL inst_cellmath__220__188__I205 (.Y(inst_cellmath__220__188__out0[3]), .A(N222), .B(N364));
MXI2X1 inst_cellmath__220__188__I206 (.Y(inst_cellmath__220__188__out0[4]), .A(N224), .B(N216), .S0(N364));
MXI2X1 inst_cellmath__220__188__I207 (.Y(inst_cellmath__220__188__out0[5]), .A(N226), .B(N218), .S0(N364));
MXI2X1 inst_cellmath__220__188__I208 (.Y(inst_cellmath__220__188__out0[6]), .A(N228), .B(N220), .S0(N364));
MXI2X1 inst_cellmath__220__188__I209 (.Y(inst_cellmath__220__188__out0[7]), .A(N230), .B(N222), .S0(N364));
MXI2X1 inst_cellmath__220__188__I210 (.Y(inst_cellmath__220__188__out0[8]), .A(N232), .B(N224), .S0(N364));
MXI2XL inst_cellmath__220__188__I211 (.Y(inst_cellmath__220__188__out0[9]), .A(N234), .B(N226), .S0(N364));
MXI2X1 inst_cellmath__220__188__I212 (.Y(inst_cellmath__220__188__out0[10]), .A(N236), .B(N228), .S0(N364));
MXI2X1 inst_cellmath__220__188__I213 (.Y(inst_cellmath__220__188__out0[11]), .A(N238), .B(N230), .S0(N364));
MXI2X1 inst_cellmath__220__188__I214 (.Y(inst_cellmath__220__188__out0[12]), .A(N240), .B(N232), .S0(N364));
MXI2X1 inst_cellmath__220__188__I215 (.Y(inst_cellmath__220__188__out0[13]), .A(N242), .B(N234), .S0(N364));
MXI2X1 inst_cellmath__220__188__I216 (.Y(inst_cellmath__220__188__out0[14]), .A(N244), .B(N236), .S0(N364));
MXI2X1 inst_cellmath__220__188__I217 (.Y(inst_cellmath__220__188__out0[15]), .A(N246), .B(N238), .S0(N360));
MXI2X1 inst_cellmath__220__188__I218 (.Y(inst_cellmath__220__188__out0[16]), .A(N248), .B(N240), .S0(N360));
MXI2XL inst_cellmath__220__188__I219 (.Y(inst_cellmath__220__188__out0[17]), .A(N249), .B(N242), .S0(N360));
MXI2X1 inst_cellmath__220__188__I220 (.Y(inst_cellmath__220__188__out0[18]), .A(N250), .B(N244), .S0(N360));
MXI2XL inst_cellmath__220__188__I221 (.Y(inst_cellmath__220__188__out0[19]), .A(N251), .B(N246), .S0(N360));
MXI2XL inst_cellmath__220__188__I222 (.Y(inst_cellmath__220__188__out0[20]), .A(N252), .B(N248), .S0(N360));
MXI2XL inst_cellmath__220__188__I223 (.Y(inst_cellmath__220__188__out0[21]), .A(N253), .B(N249), .S0(N360));
MXI2XL inst_cellmath__220__188__I224 (.Y(inst_cellmath__220__188__out0[22]), .A(N254), .B(N250), .S0(N360));
endmodule

module cynw_cm_float_cos_inst_cellmath__221__195__bdw1157874770_bdw (
	inst_cellmath__221__195__out0,
	inst_cellmath__221__195__in0
	); /* architecture "gate_level" */ 
output [6:0] inst_cellmath__221__195__out0;
input [4:0] inst_cellmath__221__195__in0;
INVXL inst_cellmath__221__195__I5 (.Y(inst_cellmath__221__195__out0[0]), .A(inst_cellmath__221__195__in0[0]));
INVXL inst_cellmath__221__195__I8 (.Y(inst_cellmath__221__195__out0[3]), .A(inst_cellmath__221__195__in0[3]));
INVXL inst_cellmath__221__195__I9 (.Y(inst_cellmath__221__195__out0[4]), .A(inst_cellmath__221__195__in0[4]));
INVXL inst_cellmath__221__195__I25 (.Y(inst_cellmath__221__195__out0[1]), .A(inst_cellmath__221__195__in0[1]));
INVXL inst_cellmath__221__195__I26 (.Y(inst_cellmath__221__195__out0[2]), .A(inst_cellmath__221__195__in0[2]));
assign inst_cellmath__221__195__out0[5] = 1'B1;
assign inst_cellmath__221__195__out0[6] = 1'B1;
endmodule

module cynw_cm_float_cos_inst_cellmath__220_2WWMM_bdw1157874770_bdw (
	inst_cellmath__220_2WWMM_out0,
	inst_cellmath__220_2WWMM_in0,
	inst_cellmath__220_2WWMM_in1,
	inst_cellmath__220_2WWMM_in2
	); /* architecture "gate_level" */ 
output [30:0] inst_cellmath__220_2WWMM_out0;
input [6:0] inst_cellmath__220_2WWMM_in0;
input [22:0] inst_cellmath__220_2WWMM_in1;
input  inst_cellmath__220_2WWMM_in2;
wire N249;
BUFX2 inst_cellmath__220_2WWMM_I144 (.Y(N249), .A(inst_cellmath__220_2WWMM_in2));
OR2XL inst_cellmath__220_2WWMM_I114 (.Y(inst_cellmath__220_2WWMM_out0[0]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[0]));
OR2XL inst_cellmath__220_2WWMM_I263 (.Y(inst_cellmath__220_2WWMM_out0[1]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[1]));
OR2XL inst_cellmath__220_2WWMM_I264 (.Y(inst_cellmath__220_2WWMM_out0[2]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[2]));
OR2XL inst_cellmath__220_2WWMM_I265 (.Y(inst_cellmath__220_2WWMM_out0[3]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[3]));
OR2XL inst_cellmath__220_2WWMM_I266 (.Y(inst_cellmath__220_2WWMM_out0[4]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[4]));
OR2XL inst_cellmath__220_2WWMM_I119 (.Y(inst_cellmath__220_2WWMM_out0[5]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[5]));
OR2XL inst_cellmath__220_2WWMM_I120 (.Y(inst_cellmath__220_2WWMM_out0[6]), .A(N249), .B(inst_cellmath__220_2WWMM_in0[6]));
NOR2BX1 inst_cellmath__220_2WWMM_I267 (.Y(inst_cellmath__220_2WWMM_out0[8]), .AN(inst_cellmath__220_2WWMM_in1[0]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I171 (.Y(inst_cellmath__220_2WWMM_out0[9]), .AN(inst_cellmath__220_2WWMM_in1[1]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I123 (.Y(inst_cellmath__220_2WWMM_out0[10]), .AN(inst_cellmath__220_2WWMM_in1[2]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I124 (.Y(inst_cellmath__220_2WWMM_out0[11]), .AN(inst_cellmath__220_2WWMM_in1[3]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I125 (.Y(inst_cellmath__220_2WWMM_out0[12]), .AN(inst_cellmath__220_2WWMM_in1[4]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I126 (.Y(inst_cellmath__220_2WWMM_out0[13]), .AN(inst_cellmath__220_2WWMM_in1[5]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I127 (.Y(inst_cellmath__220_2WWMM_out0[14]), .AN(inst_cellmath__220_2WWMM_in1[6]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I128 (.Y(inst_cellmath__220_2WWMM_out0[15]), .AN(inst_cellmath__220_2WWMM_in1[7]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I129 (.Y(inst_cellmath__220_2WWMM_out0[16]), .AN(inst_cellmath__220_2WWMM_in1[8]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I151 (.Y(inst_cellmath__220_2WWMM_out0[17]), .AN(inst_cellmath__220_2WWMM_in1[9]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I131 (.Y(inst_cellmath__220_2WWMM_out0[18]), .AN(inst_cellmath__220_2WWMM_in1[10]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I132 (.Y(inst_cellmath__220_2WWMM_out0[19]), .AN(inst_cellmath__220_2WWMM_in1[11]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I133 (.Y(inst_cellmath__220_2WWMM_out0[20]), .AN(inst_cellmath__220_2WWMM_in1[12]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I134 (.Y(inst_cellmath__220_2WWMM_out0[21]), .AN(inst_cellmath__220_2WWMM_in1[13]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I135 (.Y(inst_cellmath__220_2WWMM_out0[22]), .AN(inst_cellmath__220_2WWMM_in1[14]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I136 (.Y(inst_cellmath__220_2WWMM_out0[23]), .AN(inst_cellmath__220_2WWMM_in1[15]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I268 (.Y(inst_cellmath__220_2WWMM_out0[24]), .AN(inst_cellmath__220_2WWMM_in1[16]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I138 (.Y(inst_cellmath__220_2WWMM_out0[25]), .AN(inst_cellmath__220_2WWMM_in1[17]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I269 (.Y(inst_cellmath__220_2WWMM_out0[26]), .AN(inst_cellmath__220_2WWMM_in1[18]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I270 (.Y(inst_cellmath__220_2WWMM_out0[27]), .AN(inst_cellmath__220_2WWMM_in1[19]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I175 (.Y(inst_cellmath__220_2WWMM_out0[28]), .AN(inst_cellmath__220_2WWMM_in1[20]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I142 (.Y(inst_cellmath__220_2WWMM_out0[29]), .AN(inst_cellmath__220_2WWMM_in1[21]), .B(N249));
NOR2BX1 inst_cellmath__220_2WWMM_I143 (.Y(inst_cellmath__220_2WWMM_out0[30]), .AN(inst_cellmath__220_2WWMM_in1[22]), .B(N249));
assign inst_cellmath__220_2WWMM_out0[7] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__223__208__bdw1157874770_bdw (
	inst_cellmath__223__208__out0,
	inst_cellmath__223__208__in0,
	inst_cellmath__223__208__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__208__out0;
input [6:0] inst_cellmath__223__208__in0;
input [29:8] inst_cellmath__223__208__in1;
wire N35,N38,N39,N40,N44,N46,N47 
	,N49,N50,N51,N52,N54,N55,N56,N57 
	,N58,N59,N60,N61,N63,N65;
OR3XL inst_cellmath__223__208__I41 (.Y(N35), .A(inst_cellmath__223__208__in0[6]), .B(inst_cellmath__223__208__in0[5]), .C(inst_cellmath__223__208__in0[0]));
NOR3XL inst_cellmath__223__208__I43 (.Y(N38), .A(N35), .B(inst_cellmath__223__208__in0[1]), .C(inst_cellmath__223__208__in0[3]));
NOR2XL inst_cellmath__223__208__I7 (.Y(N39), .A(inst_cellmath__223__208__in0[4]), .B(inst_cellmath__223__208__in0[2]));
NAND2XL inst_cellmath__223__208__I8 (.Y(N40), .A(N38), .B(N39));
NOR3XL inst_cellmath__223__208__I45 (.Y(N44), .A(N40), .B(inst_cellmath__223__208__in1[8]), .C(inst_cellmath__223__208__in1[11]));
NOR3XL inst_cellmath__223__208__I46 (.Y(N46), .A(inst_cellmath__223__208__in1[9]), .B(inst_cellmath__223__208__in1[15]), .C(inst_cellmath__223__208__in1[10]));
NOR2X2 inst_cellmath__223__208__I15 (.Y(N47), .A(inst_cellmath__223__208__in1[23]), .B(inst_cellmath__223__208__in1[20]));
NOR2XL inst_cellmath__223__208__I17 (.Y(N49), .A(inst_cellmath__223__208__in1[22]), .B(inst_cellmath__223__208__in1[17]));
NOR2XL inst_cellmath__223__208__I18 (.Y(N50), .A(inst_cellmath__223__208__in1[21]), .B(inst_cellmath__223__208__in1[13]));
NOR2XL inst_cellmath__223__208__I19 (.Y(N51), .A(inst_cellmath__223__208__in1[24]), .B(inst_cellmath__223__208__in1[14]));
NAND2X1 inst_cellmath__223__208__I20 (.Y(N52), .A(N44), .B(N47));
OR3XL inst_cellmath__223__208__I47 (.Y(N54), .A(inst_cellmath__223__208__in1[16]), .B(inst_cellmath__223__208__in1[12]), .C(inst_cellmath__223__208__in1[19]));
NAND2XL inst_cellmath__223__208__I23 (.Y(N55), .A(N49), .B(N46));
NAND2XL inst_cellmath__223__208__I24 (.Y(N56), .A(N50), .B(N51));
NOR2XL inst_cellmath__223__208__I25 (.Y(N57), .A(inst_cellmath__223__208__in1[29]), .B(inst_cellmath__223__208__in1[28]));
NOR2XL inst_cellmath__223__208__I26 (.Y(N58), .A(N52), .B(inst_cellmath__223__208__in1[25]));
NOR2XL inst_cellmath__223__208__I27 (.Y(N59), .A(inst_cellmath__223__208__in1[27]), .B(inst_cellmath__223__208__in1[18]));
NOR2XL inst_cellmath__223__208__I28 (.Y(N60), .A(N55), .B(inst_cellmath__223__208__in1[26]));
NOR2XL inst_cellmath__223__208__I29 (.Y(N61), .A(N56), .B(N54));
NAND2XL inst_cellmath__223__208__I31 (.Y(N63), .A(N59), .B(N60));
NAND3X1 inst_cellmath__223__208__I115 (.Y(N65), .A(N57), .B(N58), .C(N61));
OR2XL inst_cellmath__223__208__I34 (.Y(inst_cellmath__223__208__out0[0]), .A(N63), .B(N65));
endmodule

module cynw_cm_float_cos_inst_cellmath__223__199__bdw1157874770_bdw (
	inst_cellmath__223__199__out0,
	inst_cellmath__223__199__in0,
	inst_cellmath__223__199__in1,
	inst_cellmath__223__199__in2,
	inst_cellmath__223__199__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__199__out0;
input  inst_cellmath__223__199__in0;
input [1:1] inst_cellmath__223__199__in1;
input [8:6] inst_cellmath__223__199__in2;
input [0:0] inst_cellmath__223__199__in3;
wire N2,N9,N10,N14;
NOR2XL inst_cellmath__223__199__I0 (.Y(N9), .A(inst_cellmath__223__199__in2[8]), .B(inst_cellmath__223__199__in2[7]));
NOR2XL inst_cellmath__223__199__I1 (.Y(N10), .A(inst_cellmath__223__199__in2[6]), .B(inst_cellmath__223__199__in0));
AND3XL inst_cellmath__223__199__I17 (.Y(N14), .A(N9), .B(N10), .C(inst_cellmath__223__199__in1[1]));
NAND2X2 inst_cellmath__223__199__I6 (.Y(N2), .A(N14), .B(inst_cellmath__223__199__in3[0]));
INVXL inst_cellmath__223__199__I12 (.Y(inst_cellmath__223__199__out0[0]), .A(N2));
endmodule

module cynw_cm_float_cos_inst_cellmath__224__213__bdw1157874770_bdw (
	inst_cellmath__224__213__out0,
	inst_cellmath__224__213__in0,
	inst_cellmath__224__213__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__224__213__out0;
input [0:0] inst_cellmath__224__213__in0;
input  inst_cellmath__224__213__in1;
OR2XL inst_cellmath__224__213__I0 (.Y(inst_cellmath__224__213__out0[0]), .A(inst_cellmath__224__213__in1), .B(inst_cellmath__224__213__in0[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__224__212__bdw1157874770_bdw (
	inst_cellmath__224__212__out0,
	inst_cellmath__224__212__in0,
	inst_cellmath__224__212__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__224__212__out0;
input  inst_cellmath__224__212__in0;
input [0:0] inst_cellmath__224__212__in1;
NAND2BX2 inst_cellmath__224__212__I2 (.Y(inst_cellmath__224__212__out0[0]), .AN(inst_cellmath__224__212__in0), .B(inst_cellmath__224__212__in1[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__225__215__bdw1157874770_bdw (
	inst_cellmath__225__215__out0,
	inst_cellmath__225__215__in0,
	inst_cellmath__225__215__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__225__215__out0;
input  inst_cellmath__225__215__in0,
	inst_cellmath__225__215__in1;
wire N5;
INVX1 inst_cellmath__225__215__I0 (.Y(N5), .A(inst_cellmath__225__215__in0));
NAND2X1 inst_cellmath__225__215__I1 (.Y(inst_cellmath__225__215__out0[0]), .A(N5), .B(inst_cellmath__225__215__in1));
endmodule

module cynw_cm_float_cos_inst_cellmath__228_0_bdw1157874770_bdw (
	inst_cellmath__228_0_out0,
	inst_cellmath__228_0_in0,
	inst_cellmath__228_0_in1,
	inst_cellmath__228_0_in2,
	inst_cellmath__228_0_in3
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__228_0_out0;
input [0:0] inst_cellmath__228_0_in0,
	inst_cellmath__228_0_in1,
	inst_cellmath__228_0_in2;
input [6:0] inst_cellmath__228_0_in3;
wire N99;
INVXL inst_cellmath__228_0_I28 (.Y(N99), .A(inst_cellmath__228_0_in0[0]));
AO22XL inst_cellmath__228_0_I4 (.Y(inst_cellmath__228_0_out0[0]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[0]));
AO22XL inst_cellmath__228_0_I5 (.Y(inst_cellmath__228_0_out0[1]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[1]));
AO22XL inst_cellmath__228_0_I6 (.Y(inst_cellmath__228_0_out0[2]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[2]));
AO22XL inst_cellmath__228_0_I7 (.Y(inst_cellmath__228_0_out0[3]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[3]));
AO22XL inst_cellmath__228_0_I8 (.Y(inst_cellmath__228_0_out0[4]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[4]));
AO22XL inst_cellmath__228_0_I9 (.Y(inst_cellmath__228_0_out0[5]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[5]));
AO22XL inst_cellmath__228_0_I10 (.Y(inst_cellmath__228_0_out0[6]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N99), .B1(inst_cellmath__228_0_in3[6]));
AND2XL inst_cellmath__228_0_I11 (.Y(inst_cellmath__228_0_out0[7]), .A(inst_cellmath__228_0_in2[0]), .B(inst_cellmath__228_0_in0[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__231_0_bdw1157874770_bdw (
	inst_cellmath__231_0_out0,
	inst_cellmath__231_0_in0,
	inst_cellmath__231_0_in1,
	inst_cellmath__231_0_in2,
	inst_cellmath__231_0_in3
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__231_0_out0;
input  inst_cellmath__231_0_in0;
input [0:0] inst_cellmath__231_0_in1;
input [30:8] inst_cellmath__231_0_in2;
input [46:46] inst_cellmath__231_0_in3;
wire N76,N77,N78,N79,N80,N81,N82 
	,N83,N84,N85,N86,N87,N88,N89,N90 
	,N91,N92,N93,N94,N95,N96,N97,N98 
	,N130;
INVXL inst_cellmath__231_0_I76 (.Y(N130), .A(inst_cellmath__231_0_in0));
INVXL inst_cellmath__231_0_I23 (.Y(N76), .A(inst_cellmath__231_0_in2[8]));
INVXL inst_cellmath__231_0_I24 (.Y(N77), .A(inst_cellmath__231_0_in2[9]));
INVXL inst_cellmath__231_0_I25 (.Y(N78), .A(inst_cellmath__231_0_in2[10]));
INVXL inst_cellmath__231_0_I26 (.Y(N79), .A(inst_cellmath__231_0_in2[11]));
INVXL inst_cellmath__231_0_I27 (.Y(N80), .A(inst_cellmath__231_0_in2[12]));
INVXL inst_cellmath__231_0_I28 (.Y(N81), .A(inst_cellmath__231_0_in2[13]));
INVXL inst_cellmath__231_0_I29 (.Y(N82), .A(inst_cellmath__231_0_in2[14]));
INVXL inst_cellmath__231_0_I30 (.Y(N83), .A(inst_cellmath__231_0_in2[15]));
INVXL inst_cellmath__231_0_I31 (.Y(N84), .A(inst_cellmath__231_0_in2[16]));
INVXL inst_cellmath__231_0_I32 (.Y(N85), .A(inst_cellmath__231_0_in2[17]));
INVXL inst_cellmath__231_0_I33 (.Y(N86), .A(inst_cellmath__231_0_in2[18]));
INVXL inst_cellmath__231_0_I34 (.Y(N87), .A(inst_cellmath__231_0_in2[19]));
INVXL inst_cellmath__231_0_I35 (.Y(N88), .A(inst_cellmath__231_0_in2[20]));
INVXL inst_cellmath__231_0_I36 (.Y(N89), .A(inst_cellmath__231_0_in2[21]));
INVXL inst_cellmath__231_0_I37 (.Y(N90), .A(inst_cellmath__231_0_in2[22]));
INVXL inst_cellmath__231_0_I38 (.Y(N91), .A(inst_cellmath__231_0_in2[23]));
INVXL inst_cellmath__231_0_I39 (.Y(N92), .A(inst_cellmath__231_0_in2[24]));
INVXL inst_cellmath__231_0_I40 (.Y(N93), .A(inst_cellmath__231_0_in2[25]));
INVX3 inst_cellmath__231_0_I41 (.Y(N94), .A(inst_cellmath__231_0_in2[26]));
INVXL inst_cellmath__231_0_I42 (.Y(N95), .A(inst_cellmath__231_0_in2[27]));
INVXL inst_cellmath__231_0_I43 (.Y(N96), .A(inst_cellmath__231_0_in2[28]));
INVXL inst_cellmath__231_0_I44 (.Y(N97), .A(inst_cellmath__231_0_in2[29]));
INVXL inst_cellmath__231_0_I45 (.Y(N98), .A(inst_cellmath__231_0_in2[30]));
MXI2XL inst_cellmath__231_0_I46 (.Y(inst_cellmath__231_0_out0[0]), .A(N76), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I47 (.Y(inst_cellmath__231_0_out0[1]), .A(N77), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I48 (.Y(inst_cellmath__231_0_out0[2]), .A(N78), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I49 (.Y(inst_cellmath__231_0_out0[3]), .A(N79), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I50 (.Y(inst_cellmath__231_0_out0[4]), .A(N80), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I51 (.Y(inst_cellmath__231_0_out0[5]), .A(N81), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I52 (.Y(inst_cellmath__231_0_out0[6]), .A(N82), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I53 (.Y(inst_cellmath__231_0_out0[7]), .A(N83), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I54 (.Y(inst_cellmath__231_0_out0[8]), .A(N84), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I55 (.Y(inst_cellmath__231_0_out0[9]), .A(N85), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I56 (.Y(inst_cellmath__231_0_out0[10]), .A(N86), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I57 (.Y(inst_cellmath__231_0_out0[11]), .A(N87), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I58 (.Y(inst_cellmath__231_0_out0[12]), .A(N88), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I59 (.Y(inst_cellmath__231_0_out0[13]), .A(N89), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I60 (.Y(inst_cellmath__231_0_out0[14]), .A(N90), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I61 (.Y(inst_cellmath__231_0_out0[15]), .A(N91), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I62 (.Y(inst_cellmath__231_0_out0[16]), .A(N92), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I63 (.Y(inst_cellmath__231_0_out0[17]), .A(N93), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I64 (.Y(inst_cellmath__231_0_out0[18]), .A(N94), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I65 (.Y(inst_cellmath__231_0_out0[19]), .A(N95), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I66 (.Y(inst_cellmath__231_0_out0[20]), .A(N96), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I67 (.Y(inst_cellmath__231_0_out0[21]), .A(N97), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
MXI2XL inst_cellmath__231_0_I68 (.Y(inst_cellmath__231_0_out0[22]), .A(N98), .B(N130), .S0(inst_cellmath__231_0_in1[0]));
endmodule

/* CADENCE  vrfzTA3fqBE= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



