/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:44 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_add2_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__20,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__23,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39;
wire [7:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40;
wire [8:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44;
wire [7:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49;
wire [25:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51;
wire  DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__52;
wire [5:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55;
wire [25:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56;
wire  DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__62;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63;
wire [7:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66;
wire  DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__69,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__73,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N417,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N418,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N420,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N421,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N422,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N423,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N424,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N425,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N426,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N427,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N428,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N429,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N430,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N431,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N432,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N433,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N434,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N435,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N436,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N437,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N438,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N439,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N440,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N441,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N442,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N443,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N444,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N469,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N470,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N471,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N473,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N474,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N475,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N477,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N478,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N479,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N482,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N483,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N485,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N488,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N493,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N495,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N496,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N498,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N499,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N509,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N510,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N513,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N514,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N515,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N516,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N522,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N539,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N575,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N576,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N577,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N578,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N579,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N580,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N581,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N582,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N583,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N584,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N585,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N586,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N587,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N588,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N589,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N590,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N591,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N592,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N593,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N594,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N595,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N596,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N597,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2804,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2806,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2809,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2811,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2815,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2817,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2822,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2827,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2838,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2844,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2851,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2988,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2992,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3010,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3014,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3131,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3133,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3154,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3162,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3165,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3167,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3171,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3173,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3176,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3182,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3186,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3220,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3222,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3243,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3251,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3254,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3256,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3260,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3262,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3265,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3271,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3275,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3328,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3337,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3341,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3345,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3353,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3379,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3385,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3394,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3400,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3405,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3413,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3418,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3425,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3429,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3435,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3438,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3448,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3458,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3462,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3468,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3472,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3482,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3488,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3494,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3495,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3498,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3504,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3507,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3513,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3518,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3535,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3900,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3905,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3908,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3911,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3913,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3917,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3919,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3924,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3927,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3930,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3932,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3938,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3941,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3944,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3947,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3951,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3954,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3957,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3959,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3963,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3966,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3971,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3974,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3977,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3980,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3983,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3985,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3990,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3993,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3996,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3999,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4002,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4004,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4009,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4012,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4015,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4017,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4023,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4026,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4029,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4032,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4035,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4037,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4040,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4043,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4046,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4049,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4159,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4164,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4177,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4180,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4184,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4188,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4193,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4197,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4200,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4206,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4210,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4216,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4220,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4224,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4230,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4234,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4239,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4242,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4247,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4252,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4256,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4259,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4263,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4267,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4271,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4276,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4280,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4339,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4341,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4342,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4347,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4348,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4349,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4354,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4355,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4360,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4362,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4367,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4368,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4370,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4374,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4376,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4378,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4382,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4383,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4384,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4389,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4390,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4392,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4393,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4398,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4400,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4404,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4408,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4414,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4415,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4420,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4421,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4423,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4428,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4552,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4554,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4557,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4561,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4567,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4570,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4571,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4573,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4575,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4578,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4593,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4603,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4632,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4636,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4639,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4641,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4644,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4646,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4650,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4652,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4653,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4654,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4655,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4657,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4660,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4662,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4668,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4670,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4741,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4742,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4746,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4755,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4759,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4763,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4775,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4779,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4784,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4796,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4799,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4803,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4807,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4818,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4822,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4836,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4842,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4852,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4853,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4855,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4859,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4875,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4876,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4881,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4893,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4895,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6143,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6144,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6145,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6146,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6147,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6149,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6150,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6152,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6165,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6173,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6178,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6187,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6195,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6205,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6212,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6216,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10018,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10124,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10128,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10133,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10141,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10144,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10152,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10157,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10162,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10208,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10211,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10216,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10217,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10220,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10221,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10223,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10290,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10297,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10324,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10327,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10339,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10347,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10363,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10367,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10369,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10374,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10377,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10417,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10423;
wire N3881,N4038,N4247,N4249,N4293,N4572,N4578 
	,N4892,N4894,N4901,N4903,N5139,N5145,N5154,N5398 
	,N5409,N5467,N5475,N5508,N5977,N5979,N5981,N5984 
	,N5986,N5988,N6007,N6009,N6073,N6075,N6077,N6083 
	,N6087,N6089,N6097,N6101,N6107,N6109,N6113,N6122 
	,N6124,N6129,N6133,N6135,N6143,N6147,N6156,N6158 
	,N6173,N6175,N6185,N6192,N6194,N6201,N6203,N6210 
	,N6212,N6217,N6221,N6228,N6230,N6235,N6239,N6246 
	,N6248,N6253,N6257,N6262,N6266,N6271,N6275,N6280 
	,N6284,N6289,N6295,N6298,N6304,N6331,N6341,N6349 
	,N6355,N6364,N6370,N6654,N6657,N6663,N6666,N6675 
	,N6677,N6853,N6854,N6856,N6863,N6870,N6918;
reg x_reg_23__retimed_I3276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3276_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N469;
	end
assign N6677 = x_reg_23__retimed_I3276_QOUT;
reg x_reg_23__retimed_I3275_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3275_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
	end
assign N6675 = x_reg_23__retimed_I3275_QOUT;
reg x_reg_29__retimed_I3271_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__retimed_I3271_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[6];
	end
assign N6666 = x_reg_29__retimed_I3271_QOUT;
reg x_reg_27__retimed_I3270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__retimed_I3270_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4632;
	end
assign N6663 = x_reg_27__retimed_I3270_QOUT;
reg x_reg_30__retimed_I3268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3268_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[4];
	end
assign N6657 = x_reg_30__retimed_I3268_QOUT;
reg x_reg_31__retimed_I3267_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3267_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142;
	end
assign N6654 = x_reg_31__retimed_I3267_QOUT;
reg x_reg_23__retimed_I3144_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3144_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N433;
	end
assign N6304 = x_reg_23__retimed_I3144_QOUT;
reg x_reg_23__retimed_I3141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3141_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4267;
	end
assign N6298 = x_reg_23__retimed_I3141_QOUT;
reg x_reg_23__retimed_I3140_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3140_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N441;
	end
assign N6295 = x_reg_23__retimed_I3140_QOUT;
reg x_reg_23__retimed_I3137_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3137_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4239;
	end
assign N6289 = x_reg_23__retimed_I3137_QOUT;
reg x_reg_23__retimed_I3135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3135_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4234;
	end
assign N6284 = x_reg_23__retimed_I3135_QOUT;
reg x_reg_23__retimed_I3133_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3133_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N427;
	end
assign N6280 = x_reg_23__retimed_I3133_QOUT;
reg x_reg_23__retimed_I3131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3131_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4210;
	end
assign N6275 = x_reg_23__retimed_I3131_QOUT;
reg x_reg_23__retimed_I3129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3129_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N426;
	end
assign N6271 = x_reg_23__retimed_I3129_QOUT;
reg x_reg_23__retimed_I3127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3127_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4256;
	end
assign N6266 = x_reg_23__retimed_I3127_QOUT;
reg x_reg_23__retimed_I3125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3125_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N428;
	end
assign N6262 = x_reg_23__retimed_I3125_QOUT;
reg x_reg_23__retimed_I3123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3123_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4263;
	end
assign N6257 = x_reg_23__retimed_I3123_QOUT;
reg x_reg_23__retimed_I3121_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3121_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N442;
	end
assign N6253 = x_reg_23__retimed_I3121_QOUT;
reg x_reg_23__retimed_I3119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3119_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4271;
	end
assign N6248 = x_reg_23__retimed_I3119_QOUT;
reg x_reg_23__retimed_I3118_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3118_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N424;
	end
assign N6246 = x_reg_23__retimed_I3118_QOUT;
reg x_reg_23__retimed_I3115_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3115_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4224;
	end
assign N6239 = x_reg_23__retimed_I3115_QOUT;
reg x_reg_23__retimed_I3113_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3113_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N422;
	end
assign N6235 = x_reg_23__retimed_I3113_QOUT;
reg x_reg_23__retimed_I3111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3111_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4242;
	end
assign N6230 = x_reg_23__retimed_I3111_QOUT;
reg x_reg_23__retimed_I3110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3110_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N432;
	end
assign N6228 = x_reg_23__retimed_I3110_QOUT;
reg x_reg_23__retimed_I3107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3107_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4184;
	end
assign N6221 = x_reg_23__retimed_I3107_QOUT;
reg x_reg_23__retimed_I3105_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3105_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N434;
	end
assign N6217 = x_reg_23__retimed_I3105_QOUT;
reg x_reg_30__retimed_I3103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3103_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4252;
	end
assign N6212 = x_reg_30__retimed_I3103_QOUT;
reg x_reg_30__retimed_I3102_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3102_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N437;
	end
assign N6210 = x_reg_30__retimed_I3102_QOUT;
reg x_reg_23__retimed_I3099_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3099_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4247;
	end
assign N6203 = x_reg_23__retimed_I3099_QOUT;
reg x_reg_23__retimed_I3098_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3098_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N423;
	end
assign N6201 = x_reg_23__retimed_I3098_QOUT;
reg x_reg_30__retimed_I3095_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3095_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4220;
	end
assign N6194 = x_reg_30__retimed_I3095_QOUT;
reg x_reg_30__retimed_I3094_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3094_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N431;
	end
assign N6192 = x_reg_30__retimed_I3094_QOUT;
reg x_reg_23__retimed_I3091_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3091_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0];
	end
assign N6185 = x_reg_23__retimed_I3091_QOUT;
reg x_reg_30__retimed_I3089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3089_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4276;
	end
assign N6175 = x_reg_30__retimed_I3089_QOUT;
reg x_reg_30__retimed_I3088_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3088_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N438;
	end
assign N6173 = x_reg_30__retimed_I3088_QOUT;
reg x_reg_23__retimed_I3084_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3084_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4216;
	end
assign N6158 = x_reg_23__retimed_I3084_QOUT;
reg x_reg_23__retimed_I3083_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3083_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N440;
	end
assign N6156 = x_reg_23__retimed_I3083_QOUT;
reg x_reg_30__retimed_I3080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3080_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4280;
	end
assign N6147 = x_reg_30__retimed_I3080_QOUT;
reg x_reg_30__retimed_I3078_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3078_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N429;
	end
assign N6143 = x_reg_30__retimed_I3078_QOUT;
reg x_reg_30__retimed_I3076_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3076_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4193;
	end
assign N6135 = x_reg_30__retimed_I3076_QOUT;
reg x_reg_30__retimed_I3075_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3075_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N439;
	end
assign N6133 = x_reg_30__retimed_I3075_QOUT;
reg x_reg_30__retimed_I3073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3073_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6145;
	end
assign N6129 = x_reg_30__retimed_I3073_QOUT;
reg x_reg_23__retimed_I3072_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3072_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4230;
	end
assign N6124 = x_reg_23__retimed_I3072_QOUT;
reg x_reg_23__retimed_I3071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3071_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N436;
	end
assign N6122 = x_reg_23__retimed_I3071_QOUT;
reg x_reg_23__retimed_I3068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3068_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4188;
	end
assign N6113 = x_reg_23__retimed_I3068_QOUT;
reg x_reg_23__retimed_I3066_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3066_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N425;
	end
assign N6109 = x_reg_23__retimed_I3066_QOUT;
reg x_reg_23__retimed_I3065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3065_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6146;
	end
assign N6107 = x_reg_23__retimed_I3065_QOUT;
reg x_reg_30__retimed_I3064_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3064_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4197;
	end
assign N6101 = x_reg_30__retimed_I3064_QOUT;
reg x_reg_30__retimed_I3062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3062_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N430;
	end
assign N6097 = x_reg_30__retimed_I3062_QOUT;
reg x_reg_23__retimed_I3060_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3060_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4200;
	end
assign N6089 = x_reg_23__retimed_I3060_QOUT;
reg x_reg_23__retimed_I3059_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3059_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N421;
	end
assign N6087 = x_reg_23__retimed_I3059_QOUT;
reg x_reg_23__retimed_I3057_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3057_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6143;
	end
assign N6083 = x_reg_23__retimed_I3057_QOUT;
reg x_reg_30__retimed_I3056_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3056_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4206;
	end
assign N6077 = x_reg_30__retimed_I3056_QOUT;
reg x_reg_30__retimed_I3055_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3055_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N435;
	end
assign N6075 = x_reg_30__retimed_I3055_QOUT;
reg x_reg_30__retimed_I3054_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3054_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6150;
	end
assign N6073 = x_reg_30__retimed_I3054_QOUT;
reg x_reg_30__retimed_I3041_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3041_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N443;
	end
assign N6009 = x_reg_30__retimed_I3041_QOUT;
reg x_reg_30__retimed_I3040_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I3040_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6144;
	end
assign N6007 = x_reg_30__retimed_I3040_QOUT;
reg x_reg_23__retimed_I3036_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3036_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4177;
	end
assign N5988 = x_reg_23__retimed_I3036_QOUT;
reg x_reg_23__retimed_I3035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3035_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N420;
	end
assign N5986 = x_reg_23__retimed_I3035_QOUT;
reg x_reg_23__retimed_I3034_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3034_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6152;
	end
assign N5984 = x_reg_23__retimed_I3034_QOUT;
reg x_reg_23__retimed_I3033_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3033_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6147;
	end
assign N5981 = x_reg_23__retimed_I3033_QOUT;
reg x_reg_23__retimed_I3032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3032_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4259;
	end
assign N5979 = x_reg_23__retimed_I3032_QOUT;
reg x_reg_23__retimed_I3031_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3031_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[0];
	end
assign N5977 = x_reg_23__retimed_I3031_QOUT;
reg x_reg_23__retimed_I2872_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I2872_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[0];
	end
assign N5508 = x_reg_23__retimed_I2872_QOUT;
reg x_reg_24__retimed_I2861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I2861_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4652;
	end
assign N5475 = x_reg_24__retimed_I2861_QOUT;
reg x_reg_30__retimed_I2858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2858_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1];
	end
assign N5467 = x_reg_30__retimed_I2858_QOUT;
reg x_reg_30__retimed_I2849_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2849_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4571;
	end
assign N5409 = x_reg_30__retimed_I2849_QOUT;
reg x_reg_25__retimed_I2844_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__retimed_I2844_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4644;
	end
assign N5398 = x_reg_25__retimed_I2844_QOUT;
reg x_reg_30__retimed_I2767_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2767_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3];
	end
assign N5154 = x_reg_30__retimed_I2767_QOUT;
reg x_reg_26__retimed_I2763_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__retimed_I2763_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4668;
	end
assign N5145 = x_reg_26__retimed_I2763_QOUT;
reg x_reg_30__retimed_I2761_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2761_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4593;
	end
assign N5139 = x_reg_30__retimed_I2761_QOUT;
reg x_reg_31__retimed_I2682_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I2682_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4159;
	end
assign N4903 = x_reg_31__retimed_I2682_QOUT;
reg x_reg_31__retimed_I2681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I2681_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4164;
	end
assign N4901 = x_reg_31__retimed_I2681_QOUT;
reg x_reg_30__retimed_I2678_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2678_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21;
	end
assign N4894 = x_reg_30__retimed_I2678_QOUT;
reg x_reg_30__retimed_I2677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2677_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24;
	end
assign N4892 = x_reg_30__retimed_I2677_QOUT;
reg x_reg_28__retimed_I2572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__retimed_I2572_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4660;
	end
assign N4578 = x_reg_28__retimed_I2572_QOUT;
reg x_reg_30__retimed_I2570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2570_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[5];
	end
assign N4572 = x_reg_30__retimed_I2570_QOUT;
reg x_reg_30__retimed_I2465_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2465_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N498;
	end
assign N4293 = x_reg_30__retimed_I2465_QOUT;
reg x_reg_31__retimed_I2460_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I2460_QOUT <= b_sign;
	end
assign N4249 = x_reg_31__retimed_I2460_QOUT;
reg x_reg_31__retimed_I2459_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I2459_QOUT <= a_sign;
	end
assign N4247 = x_reg_31__retimed_I2459_QOUT;
reg x_reg_30__retimed_I2367_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I2367_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[7];
	end
assign N4038 = x_reg_30__retimed_I2367_QOUT;
reg x_reg_21__retimed_I2300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I2300_QOUT <= DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__62;
	end
assign N3881 = x_reg_21__retimed_I2300_QOUT;
assign N6853 = !N3881;
assign N6854 = !N6853;
assign bdw_enable = !astall;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3131 = !(b_exp[0] & b_exp[1]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3133 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6187 = !((b_exp[7] & b_exp[6]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3133);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3131 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6187);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3167 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3171 = !(((b_man[0] | b_man[1]) | b_man[2]) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3167);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3154 = !(b_man[10] | b_man[9]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3173 = !(b_man[6] | b_man[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3162 = !(b_man[8] | b_man[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3182 = !(b_man[4] | b_man[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3165 = !(((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3154 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3173) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3162) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3182);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3176 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3186 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32 = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3171) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3165) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3176) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3186);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__23 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10018 = !a_exp[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10018;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3220 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019 & a_exp[1]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3222 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6195 = !((a_exp[7] & a_exp[6]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3222);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3220 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6195);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3256 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3260 = !(((a_man[0] | a_man[1]) | a_man[2]) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3256);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3243 = !(a_man[10] | a_man[9]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3262 = !(a_man[6] | a_man[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3251 = !(a_man[8] | a_man[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3271 = !(a_man[4] | a_man[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3254 = !(((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3243 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3262) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3251) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3271);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3265 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3275 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29 = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3260) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3254) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3265) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3275);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__20 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0] = a_sign ^ b_sign;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N495 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__62 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__23 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__20) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N495;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3010 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3014 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3010 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3014);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2988 = ((a_exp[7] | a_exp[1]) | a_exp[6]) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2992 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2988 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2992);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504 = !a_exp[4];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362 = !a_exp[3];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502 = !a_exp[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501 = !a_exp[1];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500 = !a_exp[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6178 = !(b_exp[0] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2806 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6178;
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2851, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[1]} = {1'B0, b_exp[1]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2806};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2822, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[2]} = {1'B0, b_exp[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2851};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2844, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10367} = {1'B0, b_exp[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2822};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2815, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[4]} = {1'B0, b_exp[4]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2844};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3328 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[4];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507 = !a_exp[7];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506 = !a_exp[6];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505 = !a_exp[5];
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2838, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[5]} = {1'B0, b_exp[5]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2815};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2809, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[6]} = {1'B0, b_exp[6]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2838};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10347, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[7]} = {1'B0, b_exp[7]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2809};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10347;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8];
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2817, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N509} = {1'B0, b_exp[0]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2811, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N510} = {1'B0, b_exp[1]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2817};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10327, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10377} = {1'B0, b_exp[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2811};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2804, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10339} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362} + {1'B0, b_exp[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10327};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2827, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N513} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504} + {1'B0, b_exp[4]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2804};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3328) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N513 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10324 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10367;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10339 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10324 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350);
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10290, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N514} = {1'B0, b_exp[5]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2827};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10297, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N515} = {1'B0, b_exp[6]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10290};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3345 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[6];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10141 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N515 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3345));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3337 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[5];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10128 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N514 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3337));
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N516} = {1'B0, b_exp[7]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10297};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3353 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[7];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10152 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N516 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3353));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10141 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10128) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10152);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10374 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10377 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10374 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3341 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[1];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[1] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3341) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N510 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[1];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[20] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[19]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[19]);
assign N6856 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[18]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[18]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[19] = !N6856;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[0] = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500 ^ b_exp[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[0] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8] & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N509) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[0] & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[19]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[20]);
assign N6863 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[17]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[17]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[18] = !N6863;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[17] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[16]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[16]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[17]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[18]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[23] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[22]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[22]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[23]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[22] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[21]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[21]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[21] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[20]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[20]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[21]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[22]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10423 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N539 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10423);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[17] = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N539;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N591 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[16]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[16]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[17] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N591) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[18]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[19]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[16] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[15]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[15]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[16]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[17]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[22]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[23]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[20]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[21]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[16] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N590 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[15]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[15]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[16] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N590) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[15] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[14]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[14]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[15]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[16]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3535 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[15] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3535);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N589 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[14]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[14]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[15] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N589) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[14] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[13]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[13]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[14]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[15]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3498 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[14] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3498);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N588 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[13]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[13]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[14] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N588) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[13] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[12]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[12]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[13]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[14]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3462 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[13] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3462);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N587 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[12]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[12]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[13] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N587) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[12] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[11]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[11]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[12]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[13]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3429 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[12] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3429);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N586 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[11]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[11]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[12] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N586) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[11] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842 & a_man[10]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842) & b_man[10]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[11]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[12]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3394 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[11] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3394);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N585 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[10]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[10]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[11] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N585) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign N6870 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[9]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[9]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[10] = !N6870;
assign N6355 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[10]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[11]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420 = !N6355;
assign N6364 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487 = !N6364;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3518 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[10] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3518);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N584 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[9]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[9]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[10] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N584) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[9] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[8]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[8]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[9]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[10]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3482 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[9] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3482);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N583 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[8]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[8]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[9] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N583) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[8] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[7]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[8]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[9]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3448 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[8] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3448 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[8] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[8]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N582 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[7]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[8] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N582) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[7] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[6]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[7]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[8]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3418 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3413 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3418 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[7] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3413 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[7] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[7]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N581 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[6]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[7] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N581) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[6] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[5]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[6]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3385 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3379 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3385 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[6] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3379 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[6] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[6]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N580 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[5]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[6] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N580) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[5] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[4]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[4]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[5]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3507 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3504 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3507 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[5] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3504 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[5] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[5]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N579 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[4]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[4]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[5] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N579) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[4] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[3]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[4]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3472 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3468 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3472 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[4] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3468 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[4] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[4];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N578 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[3]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[4] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N578) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[3] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[2]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[2]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[3]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[4]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3405 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3438 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3405 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3435 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3438 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[3] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3435 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[3] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[3];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N577 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[2]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[2]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[3] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N577) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign N6370 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[1]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[1]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[2] = !N6370;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[2]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10363 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10369 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10363 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3400 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10369 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[2] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3400 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[2] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N576 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[1]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[1]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[2] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N576) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10133 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10124 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[1] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & a_man[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & b_man[0]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3425 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[1]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[2]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3495 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3425 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10162 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3495 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10157 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10144 = !(((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10162 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10157);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[1] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10133 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10124) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10144);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N575 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[0]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[1] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N575) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N522 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3513 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[1]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3458 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3513 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3494 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3458 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3488 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3494 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[0] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3488 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[0] = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[0] & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N522;
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4035, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[0]};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4015, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[1]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[1]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4035};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3930, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4015};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3996, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3930};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3911, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[4]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[4]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3996};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3977, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[5]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[5]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3911};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4043, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[6]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[6]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3977};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3957, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[7]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[7]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4043};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4023, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[8]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[8]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3957};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3938, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[9]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[9]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4023};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4004, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[10]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[10]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3938};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3919, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[11]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[11]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4004};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3985, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[12]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[12]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3919};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3900, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[13]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[13]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3985};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3966, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[14]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[14]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3900};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4032, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[15]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[15]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3966};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3947, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[16]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[16]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4032};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4012, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[17]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[17]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3947};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4230 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[24] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[23] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N597 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[22]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[22]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[23] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N597) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[22] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N596 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[21]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[21]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[22] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N596) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[21] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N595 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[20]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[20]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[21] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N595) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[20] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N594 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[19]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[19]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[20] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N594) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[19] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N593 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[18]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[18]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[19] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N593) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[18] = !((((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772)) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N592 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_man[17]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_man[17]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[18] = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N592) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24];
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4002, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N420} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[1]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[1]};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3917, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N421} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4002};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3983, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N422} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3917};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4049, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N423} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[4]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[4]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3983};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3963, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N424} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[5]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[5]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4049};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4029, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N425} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[6]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[6]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3963};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3944, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N426} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[7]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[7]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4029};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4009, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N427} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[8]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[8]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3944};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3924, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N428} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[9]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[9]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4009};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3990, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N429} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[10]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[10]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3924};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3905, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N430} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[11]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[11]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3990};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3971, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N431} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[12]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[12]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3905};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4037, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N432} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[13]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[13]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3971};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3951, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N433} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[14]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[14]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4037};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4017, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N434} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[15]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[15]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3951};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3932, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N435} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[16]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[16]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4017};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3999, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N436} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[17]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[17]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3932};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3913, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N437} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[18]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[18]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3999};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3980, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N438} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[19]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[19]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3913};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4046, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N439} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[20]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[20]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3980};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3959, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N440} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[21]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[21]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4046};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4026, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N441} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[22]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[22]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3959};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3941, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N442} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[23]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[23]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4026};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N444, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N443} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[24]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3941};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[25] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N444;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[25];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6144 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[25];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6149 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6150 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6149;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17] = (N6124 & N6007) | (N6073 & N6122);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4206 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16] = (N6077 & N6007) | (N6073 & N6075);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4267 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6143 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6165 = !((N6083 & N6298) | (N6073 & N6304));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6165;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4184 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6145 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N485 = !((N6073 & N6217) | (N6221 & N6129));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N485;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4197 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign N6918 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6152 = !N6918;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11] = (N6101 & N6083) | (N6097 & N5984);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4280 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6146 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10] = (N6147 & N6107) | (N6143 & N5984);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4242 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N483 = !((N6228 & N5984) | (N6230 & N6129));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N483;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4220 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N482 = !((N6192 & N5984) | (N6194 & N6129));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N482;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148 = !N6654;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25] = !(N6185 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148);
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3927, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[18]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[18]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4012};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3993, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[19]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[19]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3927};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3908, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[20]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[20]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3993};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3974, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[21]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[21]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3908};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4040, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[22]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[22]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3974};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3954, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[23]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[23]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4040};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N469 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24] ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[24]) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3954;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4180 = !((N6677 & N6185) | ((!N6677) & N6675));
assign N6331 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4180 & N6007) | (N6009 & N6073));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24] = !N6331;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4263 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N493 = !((N6073 & N6253) | (N6257 & N6007));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N493;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4239 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6173 = !((N6083 & N6289) | (N6073 & N6295));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6173;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4216 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21] = (N6158 & N6083) | (N6073 & N6156);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4193 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20] = (N6135 & N6129) | (N5984 & N6133);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4276 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19] = (N6175 & N6007) | (N6073 & N6173);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4252 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N488 = !((N6210 & N5984) | (N6212 & N6129));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N488;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4256 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N479 = !((N6262 & N6073) | (N6266 & N6107));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N479;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4234 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N478 = !((N6073 & N6280) | (N6284 & N6107));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N478;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4210 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N477 = !((N6073 & N6271) | (N6275 & N6107));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N477;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4188 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign N6341 = !((N6107 & N6113) | (N6109 & N5984));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6] = !N6341;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4271 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6147 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N475 = !((N6246 & N5984) | (N6248 & N5981));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N475;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4247 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N474 = !((N6201 & N5984) | (N6203 & N5981));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N474;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4224 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N473 = !((N5984 & N6235) | (N6239 & N5981));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N473;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4200 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign N6349 = !((N6083 & N6089) | (N5984 & N6087));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2] = !N6349;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4420 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352 & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4354 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4374 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4393 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4354) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4374);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2] = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4420) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4393);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6212 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6212;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4384 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336 & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4376 = (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4384);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4415 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395 & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4339 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4360 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4415 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4339);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4348 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359 & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4367 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4389 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4348 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4367);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4342 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4360 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4389);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569 = !(((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4376)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4342));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4370 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4392 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4414 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4370) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20])) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4392);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4400 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4423 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4347 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4400) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24])) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4423);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4414) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4347);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10223 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4408 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4428 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4355 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4408) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12])) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4428);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4341 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4362 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4383 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4341) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16])) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4362);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4355)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4383);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10211 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10221 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10223 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10211);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4259 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N470 = !((N5977 & N5984) | (N5979 & N5981));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N470;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4177 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N471 = !((N5986 & N5984) | (N5988 & N5981));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1] = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N471;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10217 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4349 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4368 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4390 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4349) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4])) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4368);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4378 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4398 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4421 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4378) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8])) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4398);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10220 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4390) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4421);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10217) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10220);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10208 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10221 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10208);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4775 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4775;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1] | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4] = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4382 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407 & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4404 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[3] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4382 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4404);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[3];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4779 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4779 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4741 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4741 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4852 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4803 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4852 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4818 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4818 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4742 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4803 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4796 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4742 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4799 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4799 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4763 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4763 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4875 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4875 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4836 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4836 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[24] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4796 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N498 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[7] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[7]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[4] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[4]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[4]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[2]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[2]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[3]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4603 = ((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[7] & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[4]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2]) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[6] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[6]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4593 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4603 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[5] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[5]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[1]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & a_exp[1]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6205 = !((N4572 & N5467) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N499 = !(N5139 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6205);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77 = ((N4892 | N4894) | N3881) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N499;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[5] = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[3];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4570 = N5154 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4573 = N5467 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[0] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914 & b_exp[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10216 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[0] = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417)) | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10216);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4578 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[0] & (!N5508));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4561 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4573) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4578)) | ((!N5467) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4571 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4557 = N5409 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4567 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4557 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4561) | (N5409 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4575 = ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4570) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4567)) | ((!N5154) & (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566 = !N6657;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4554 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4552 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4554 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4575) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__73 = !(((N4038 | N6666) | N4572) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4552);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 = !(((N4293 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[5]) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__73);
assign x[22] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[24]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4876 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4759 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4876 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856 = DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4895 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4895 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[23] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4759 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[21] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[23]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4893 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4859 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4859 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[22] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4893 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[20] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[22]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4855 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4822 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4822 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[21] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4855 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[19] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[21]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4784 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4784 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[20] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[18] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[20]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4746 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4746 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[19] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[17] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[19]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4881 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4881 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[18] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[16] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[18]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4842 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4842 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[17] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[15] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[17]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4807 = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1]);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4807 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[16] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[14] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[16]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[15] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[13] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[15]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[14] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[12] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[14]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[13] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[11] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[13]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[12] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[10] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[12]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[11] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[9] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[11]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[10] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[8] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[10]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[9] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[7] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[9]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[8] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[6] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[8]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[7] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[5] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[7]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[6] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[4] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[6]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4755 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[5] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4755 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[3] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[5]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4853 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[4] = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4853 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
assign x[2] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[4]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[3] = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871);
assign x[1] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[3]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[2] = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758 | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831);
assign x[0] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[2]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & N6854);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6216 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4654 = !N6666;
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4657, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4644} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1]};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4632, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4668} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3]} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4657};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4650, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4639} = {1'B0, N6657} + {1'B0, N6663};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4660 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[5];
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4652 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1];
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4653, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[0]} = {1'B0, N5508} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4646, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[1]} = {1'B0, N5475} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4653};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4670, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[2]} = {1'B0, N5398} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4646};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4641, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[3]} = {1'B0, N5145} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4670};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4662, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[4]} = {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4639} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4641};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4636, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[5]} = {1'B0, N4578} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4650} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4662};
assign {DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4655, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[6]} = {1'B0, N4572} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4654} + {1'B0, DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4636};
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[7] = ((!N4038) ^ N6666) ^ DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4655;
assign x[30] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6216) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[7] & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72);
assign x[29] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[6]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign x[28] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[5]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign x[27] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[4]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign x[26] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[3]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign x[25] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[2]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign x[24] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[1]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign x[23] = (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[0]) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72) & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77);
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10417 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888 = !DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10417;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4159 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888 & b_sign) | (a_sign & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N418 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28 | (!a_sign));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N417 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31 | (!b_sign));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4164 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N418) | (DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N417 & DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__52 = !((DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148 & N4901) | ((!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148) & N4903));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N496 = !(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[5] | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__52));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__69 = (N4249 & N4247) | DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N496;
assign x[31] = !(N6854 | (!DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__69));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[3] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[2] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[3] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[4] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[5] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[6] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[7] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[0] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[24] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[1] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[9] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[10] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[11] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[12] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[13] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[14] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[15] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[16] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[17] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[18] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[19] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[20] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[21] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[22] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[23] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[24] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[1] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[0] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[1] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[2] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[3] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[4] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[5] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[6] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[7] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[8] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[9] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[10] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[11] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[12] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[13] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[14] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[15] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[16] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[17] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[18] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[19] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[20] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[21] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[22] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[23] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[24] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[0] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[1] = 1'B0;
endmodule

/* CADENCE  ubb0TAvcqx0= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



