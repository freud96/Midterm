/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:19:40 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_add2_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
wire  inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__23,
	inst_cellmath__24,
	inst_cellmath__27,
	inst_cellmath__28,
	inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__32;
wire [24:0] inst_cellmath__39;
wire [7:0] inst_cellmath__40;
wire [8:0] inst_cellmath__44;
wire [7:0] inst_cellmath__47;
wire [24:0] inst_cellmath__48,
	inst_cellmath__49;
wire [25:0] inst_cellmath__51;
wire  inst_cellmath__52;
wire [5:0] inst_delta;
wire [24:0] inst_cellmath__55;
wire [25:0] inst_cellmath__56;
wire  inst_cellmath__62;
wire [24:0] inst_cellmath__63;
wire [7:0] inst_cellmath__66;
wire  inst_cellmath__73,
	inst_cellmath__77;
wire N417,N418,N419,N420,N423,N424,N425 
	,N426,N427,N428,N429,N430,N431,N432,N433 
	,N434,N435,N436,N437,N438,N439,N440,N441 
	,N442,N443,N444,N445,N446,N447,N448,N449 
	,N450,N451,N452,N453,N454,N455,N456,N457 
	,N458,N459,N460,N461,N462,N463,N464,N465 
	,N466,N467,N468,N469,N474,N475,N476,N477 
	,N478,N479,N482,N483,N484,N487,N489,N490 
	,N491,N494,N496,N498,N499,N500,N501,N502 
	,N503,N504,N505,N506,N507,N511,N512,N513 
	,N514,N515,N516,N517,N522,N575,N576,N577 
	,N578,N579,N580,N581,N582,N583,N584,N585 
	,N586,N587,N588,N589,N590,N591,N592,N593 
	,N594,N595,N596,N597,N2396,N2397,N3782,N3783 
	,N3786,N3787,N3788,N3790,N3791,N3792,N3793,N3794 
	,N3796,N3797,N3798,N3800,N3801,N3802,N3806,N3807 
	,N3808,N3810,N3811,N3812,N3815,N3816,N3817,N3820 
	,N3821,N3823,N3824,N3825,N3826,N3829,N3832,N3833 
	,N3835,N3837,N3841,N3842,N3845,N3846,N3847,N3851 
	,N3852,N3854,N3857,N3858,N3859,N3860,N3863,N3867 
	,N3868,N3870,N3873,N3874,N3876,N3877,N3879,N3880 
	,N3883,N3884,N3885,N3888,N4022,N4085,N4090,N4094 
	,N4097,N4107,N4112,N4116,N4119,N4170,N4237,N4241 
	,N4262,N4272,N4279,N4283,N4289,N4291,N4301,N4338 
	,N4340,N4361,N4371,N4378,N4382,N4388,N4390,N4400 
	,N4450,N4474,N4509,N4511,N4513,N4514,N4516,N4518 
	,N4519,N4520,N4522,N4523,N4526,N4527,N4528,N4530 
	,N4532,N4533,N4534,N4536,N4538,N4539,N4540,N4542 
	,N4543,N4545,N4547,N4548,N4550,N4552,N4553,N4554 
	,N4556,N4558,N4559,N4561,N4562,N4563,N4566,N4567 
	,N4568,N4570,N4571,N4572,N4574,N4575,N4577,N4578 
	,N4579,N4580,N4582,N4583,N4584,N4587,N4588,N4589 
	,N4591,N4592,N4594,N4596,N4597,N4600,N4601,N4602 
	,N4603,N4605,N4606,N4607,N4609,N4610,N4611,N4613 
	,N4614,N4615,N4617,N4618,N4619,N4621,N4622,N4624 
	,N4626,N4627,N4628,N4630,N4631,N4632,N4633,N4636 
	,N4637,N4638,N4640,N4643,N4644,N4645,N4647,N4648 
	,N4650,N4651,N4653,N4654,N4655,N4657,N4659,N4660 
	,N4662,N4663,N4665,N4666,N4668,N4836,N4897,N5032 
	,N5033,N5034,N5035,N5037,N5039,N5040,N5041,N5044 
	,N5045,N5046,N5047,N5049,N5051,N5053,N5054,N5057 
	,N5058,N5059,N5060,N5062,N5064,N5065,N5066,N5067 
	,N5069,N5070,N5072,N5073,N5074,N5075,N5076,N5078 
	,N5079,N5080,N5081,N5084,N5085,N5086,N5087,N5088 
	,N5090,N5093,N5094,N5095,N5096,N5097,N5099,N5101 
	,N5102,N5103,N5104,N5105,N5106,N5108,N5110,N5111 
	,N5112,N5114,N5115,N5117,N5118,N5119,N5120,N5122 
	,N5123,N5124,N5126,N5129,N5130,N5131,N5132,N5133 
	,N5134,N5136,N5137,N5139,N5141,N5143,N5144,N5146 
	,N5147,N5148,N5149,N5150,N5151,N5152,N5154,N5155 
	,N5157,N5158,N5159,N5160,N5161,N5163,N5165,N5166 
	,N5167,N5168,N5169,N5170,N5171,N5172,N5174,N5176 
	,N5177,N5178,N5179,N5180,N5183,N5184,N5187,N5189 
	,N5190,N5191,N5192,N5193,N5194,N5196,N5198,N5199 
	,N5200,N5201,N5203,N5205,N5206,N5207,N5208,N5209 
	,N5210,N5211,N5214,N5215,N5216,N5217,N5218,N5220 
	,N5222,N5223,N5225,N5228,N5229,N5230,N5231,N5233 
	,N5235,N5236,N5237,N5239,N5241,N5242,N5243,N5246 
	,N5247,N5248,N5250,N5253,N5254,N5255,N5257,N5258 
	,N5259,N5260,N5262,N5263,N5265,N5267,N5269,N5270 
	,N5271,N5272,N5273,N5274,N5276,N5277,N5279,N5280 
	,N5281,N5282,N5283,N5286,N5287,N5288,N5289,N5290 
	,N5291,N5293,N5294,N5296,N5297,N5298,N5299,N5300 
	,N5301,N5303,N5305,N5306,N5307,N5308,N5310,N5311 
	,N5313,N5314,N5315,N5316,N5317,N5318,N5319,N5321 
	,N5323,N5324,N5325,N5326,N5328,N5330,N5331,N5332 
	,N5333,N5334,N5336,N5338,N5339,N5340,N5342,N5344 
	,N5346,N5347,N5348,N5349,N5350,N5352,N5353,N5354 
	,N5355,N5358,N5359,N5360,N5361,N5362,N5364,N5365 
	,N5368,N5369,N5370,N5371,N5373,N5375,N5376,N5377 
	,N5379,N5380,N5381,N5383,N5384,N5385,N5387,N5388 
	,N5390,N5391,N5392,N5394,N5395,N5397,N5398,N5399 
	,N5400,N5402,N5403,N5404,N5405,N5406,N5408,N5410 
	,N5411,N5412,N5415,N5416,N5417,N5418,N5419,N5420 
	,N5421,N5423,N5425,N5426,N5430,N5431,N5432,N5433 
	,N5434,N5435,N5436,N5437,N5438,N5439,N5814,N5817 
	,N5829,N5832,N5836,N5840,N5845,N5849,N5850,N5858 
	,N5863,N5869,N5873,N5883,N5887,N5892,N5895,N5901 
	,N5906,N5911,N5914,N5918,N5922,N5927,N5932,N5936 
	,N5997,N5998,N6000,N6001,N6003,N6005,N6007,N6009 
	,N6010,N6011,N6013,N6014,N6016,N6017,N6019,N6021 
	,N6022,N6024,N6026,N6028,N6029,N6030,N6032,N6033 
	,N6034,N6036,N6037,N6040,N6042,N6044,N6045,N6046 
	,N6047,N6050,N6051,N6052,N6054,N6055,N6057,N6059 
	,N6060,N6062,N6063,N6064,N6066,N6067,N6069,N6070 
	,N6072,N6073,N6074,N6076,N6077,N6079,N6080,N6082 
	,N6083,N6085,N6086,N6088,N6090,N6171,N6186,N6189 
	,N6192,N6198,N6201,N6207,N6211,N6217,N6223,N6227 
	,N6256,N6257,N6259,N6260,N6264,N6265,N6266,N6270 
	,N6272,N6273,N6274,N6275,N6277,N6279,N6280,N6284 
	,N6286,N6288,N6290,N6315,N6325,N6348,N6354,N6361 
	,N6362,N6363,N6365,N6367,N6369,N6370,N6371,N6372 
	,N6374,N6375,N6376,N6377,N6380,N6381,N6382,N6384 
	,N6385,N6386,N6387,N6388,N6389,N6391,N6392,N6394 
	,N6395,N6396,N6398,N6399,N6400,N6402,N6404,N6405 
	,N6407,N6408,N6409,N6411,N6412,N6413,N6414,N6415 
	,N6417,N6418,N6419,N6421,N6422,N6423,N6424,N6425 
	,N6429,N6430,N6431,N6434,N6436,N6437,N6439,N6511 
	,N6512,N6518,N6552,N6554,N6555,N6557,N6559,N6561 
	,N6563,N6564,N6565,N6569,N6570,N6572,N6573,N6575 
	,N6576,N6577,N6579,N6581,N6583,N6585,N6587,N6588 
	,N6589,N6591,N6592,N6593,N6596,N6598,N6600,N6602 
	,N6603,N6606,N6607,N6608,N6610,N6611,N6613,N6614 
	,N6616,N6618,N6621,N6623,N6625,N6627,N6629,N6630 
	,N6631,N6632,N6634,N6635,N6637,N6639,N6641,N6642 
	,N6646,N6647,N6648,N6650,N6652,N6653,N6655,N6658 
	,N6660,N6661,N6662,N6663,N6666,N6667,N6669,N6670 
	,N6672,N6673,N6676,N6677,N6679,N6681,N6683,N6684 
	,N6686,N6688,N6689,N6691,N6693,N6695,N6696,N6699 
	,N6700,N6704,N6705,N6706,N6708,N6709,N6711,N6712 
	,N6713,N6715,N6716,N6720,N6722,N6888,N6906,N6921 
	,N6922,N8709,N8716,N8754,N8755,N8756,N8758,N8759 
	,N8760,N8764,N8772,N8777,N8783,N8789,N8813,N14148 
	,N14157,N14169,N14173,N14181,N14209,N14214,N14222,N14225 
	,N14232,N14264,N14270,N14271,N14283,N14301,N14303,N14309 
	,N14317,N14319,N14334,N14357,N14358,N14360,N14362,N14365 
	,N14367,N14368,N14373,N14377,N14394,N14397,N14401,N14406 
	,N14418,N14434,N14435,N14440,N14446,N14451,N14455,N14496 
	,N14499,N14504,N14508,N14511,N14514,N14533,N14535,N14539 
	,N14550,N14560,N14570,N14573,N14619,N14623,N14630,N14636 
	,N14642,N14648,N14654,N14662;
CLKINVX12 cynw_cm_float_add2_I1 (.Y(N501), .A(a_exp[1]));
CLKINVX6 cynw_cm_float_add2_I4 (.Y(N504), .A(a_exp[4]));
CLKINVX8 cynw_cm_float_add2_I5 (.Y(N505), .A(a_exp[5]));
CLKINVX6 cynw_cm_float_add2_I6 (.Y(N506), .A(a_exp[6]));
INVX1 cynw_cm_float_add2_I7 (.Y(N507), .A(a_exp[7]));
CLKINVX8 inst_cellmath__43_1_I8634 (.Y(N502), .A(a_exp[2]));
NAND2X8 inst_cellmath__43_1_I590 (.Y(N3883), .A(b_exp[2]), .B(N502));
NOR2X2 inst_cellmath__43_1_I593 (.Y(N3845), .A(b_exp[4]), .B(N504));
NAND2X4 inst_cellmath__43_1_I594 (.Y(N3867), .A(b_exp[4]), .B(N504));
NOR2X2 inst_cellmath__43_1_I595 (.Y(N3786), .A(b_exp[5]), .B(N505));
NAND2X6 inst_cellmath__43_1_I596 (.Y(N3810), .A(b_exp[5]), .B(N505));
NOR2X1 inst_cellmath__43_1_I597 (.Y(N3833), .A(b_exp[6]), .B(N506));
NAND2X8 inst_cellmath__43_1_I598 (.Y(N3854), .A(b_exp[6]), .B(N506));
NAND2X4 inst_cellmath__43_1_I8446 (.Y(N3835), .A(b_exp[1]), .B(N501));
CLKINVX6 inst_cellmath__43_1_I8440 (.Y(N500), .A(a_exp[0]));
NAND2XL inst_cellmath__43_1_I8444 (.Y(N3790), .A(b_exp[0]), .B(N500));
NOR2X8 inst_cellmath__43_1_I8445 (.Y(N3815), .A(b_exp[1]), .B(N501));
AOI21X1 inst_cellmath__43_1_I601 (.Y(N3888), .A0(N3790), .A1(N3835), .B0(N3815));
CLKINVX12 inst_cellmath__43_1_I8635 (.Y(N503), .A(a_exp[3]));
NOR2X2 inst_cellmath__43_1_I8636 (.Y(N3857), .A(b_exp[2]), .B(N502));
NOR2X6 inst_cellmath__43_1_I8637 (.Y(N3801), .A(b_exp[3]), .B(N503));
NAND2X4 inst_cellmath__43_1_I8638 (.Y(N3823), .A(b_exp[3]), .B(N503));
AOI21X1 inst_cellmath__43_1_I8639 (.Y(N3874), .A0(N3823), .A1(N3857), .B0(N3801));
NAND2XL inst_cellmath__43_1_I603 (.Y(N3793), .A(N3823), .B(N3883));
AOI21XL inst_cellmath__43_1_I604 (.Y(N3859), .A0(N3845), .A1(N3810), .B0(N3786));
NAND2XL inst_cellmath__43_1_I605 (.Y(N3884), .A(N3867), .B(N3810));
NAND2X2 inst_cellmath__43_1_I8448 (.Y(N3798), .A(b_exp[7]), .B(N507));
NOR2XL inst_cellmath__43_1_I8447 (.Y(N3879), .A(b_exp[7]), .B(N507));
AOI21XL inst_cellmath__43_1_I606 (.Y(N3846), .A0(N3798), .A1(N3833), .B0(N3879));
NAND2XL inst_cellmath__43_1_I607 (.Y(N3868), .A(N3798), .B(N3854));
INVXL inst_cellmath__43_1_I608 (.Y(N3800), .A(N3888));
OAI21XL inst_cellmath__43_1_I610 (.Y(N3821), .A0(N3884), .A1(N3874), .B0(N3859));
NOR2XL inst_cellmath__43_1_I611 (.Y(N3842), .A(N3884), .B(N3793));
AOI21XL inst_cellmath__43_1_I616 (.Y(N3796), .A0(N3842), .A1(N3800), .B0(N3821));
NAND2BXL inst_cellmath__43_1_I619 (.Y(N3832), .AN(N3857), .B(N3883));
NAND2BXL inst_cellmath__43_1_I620 (.Y(N3797), .AN(N3801), .B(N3823));
NAND2BXL inst_cellmath__43_1_I621 (.Y(N3863), .AN(N3845), .B(N3867));
NAND2BXL inst_cellmath__43_1_I622 (.Y(N3829), .AN(N3786), .B(N3810));
NAND2BXL inst_cellmath__43_1_I623 (.Y(N3792), .AN(N3833), .B(N3854));
NAND2BXL inst_cellmath__43_1_I624 (.Y(N3858), .AN(N3879), .B(N3798));
XOR2XL inst_cellmath__43_1_I627 (.Y(N511), .A(N3800), .B(N3832));
OAI21X1 inst_cellmath__43_1_I8554 (.Y(N3880), .A0(N3793), .A1(N3888), .B0(N3874));
XOR2XL inst_cellmath__43_1_I628 (.Y(N513), .A(N3880), .B(N3863));
XNOR2X1 inst_cellmath__43_1_I629 (.Y(N515), .A(N3796), .B(N3792));
OAI21X1 inst_cellmath__43_1_I8555 (.Y(N14394), .A0(N3868), .A1(N3859), .B0(N3846));
NOR2X1 inst_cellmath__43_1_I8556 (.Y(N14397), .A(N3868), .B(N3884));
AO21X1 inst_cellmath__43_1_I8557 (.Y(N517), .A0(N14397), .A1(N3880), .B0(N14394));
INVX2 inst_cellmath__43_1_I8558 (.Y(N4022), .A(N517));
NAND2X1 inst_cellmath__43_1_I8559 (.Y(N14401), .A(N14397), .B(N3880));
INVX1 inst_cellmath__43_1_I8560 (.Y(N14406), .A(N14394));
NAND2X2 inst_cellmath__43_1_I8561 (.Y(N8754), .A(N14406), .B(N14401));
XNOR2X1 inst_cellmath__43_1_I632 (.Y(N3841), .A(N3883), .B(N3797));
XNOR2X1 inst_cellmath__43_1_I633 (.Y(N3820), .A(N3857), .B(N3797));
MX2XL inst_cellmath__43_1_I634 (.Y(N512), .A(N3820), .B(N3841), .S0(N3800));
XNOR2X1 inst_cellmath__43_1_I635 (.Y(N3808), .A(N3867), .B(N3829));
XNOR2X1 inst_cellmath__43_1_I636 (.Y(N3783), .A(N3845), .B(N3829));
MX2XL inst_cellmath__43_1_I637 (.Y(N514), .A(N3783), .B(N3808), .S0(N3880));
XNOR2X1 inst_cellmath__43_1_I638 (.Y(N3877), .A(N3854), .B(N3858));
XNOR2X1 inst_cellmath__43_1_I639 (.Y(N3852), .A(N3833), .B(N3858));
MX2XL inst_cellmath__43_1_I640 (.Y(N516), .A(N3877), .B(N3852), .S0(N3796));
NOR2X4 inst_cellmath__43_1_I3242 (.Y(N8709), .A(b_exp[0]), .B(N500));
AOI21X4 inst_cellmath__43_1_I642 (.Y(N3816), .A0(N3815), .A1(N3883), .B0(N3857));
NAND2X4 inst_cellmath__43_1_I643 (.Y(N3837), .A(N3835), .B(N3883));
AOI21X4 inst_cellmath__43_1_I644 (.Y(N3802), .A0(N3801), .A1(N3867), .B0(N3845));
NAND2X2 inst_cellmath__43_1_I645 (.Y(N3824), .A(N3823), .B(N3867));
AOI21X4 inst_cellmath__43_1_I646 (.Y(N3787), .A0(N3786), .A1(N3854), .B0(N3833));
NAND2X6 inst_cellmath__43_1_I647 (.Y(N3811), .A(N3810), .B(N3854));
INVX1 inst_cellmath__43_1_I8452 (.Y(N3806), .A(N8709));
OAI21X4 inst_cellmath__43_1_I649 (.Y(N3807), .A0(N3806), .A1(N3837), .B0(N3816));
INVXL buf1_A_I8754 (.Y(N14619), .A(N3807));
INVXL buf1_A_I8755 (.Y(N3791), .A(N14619));
OAI21XL inst_cellmath__43_1_I651 (.Y(N3851), .A0(N3824), .A1(N3816), .B0(N3802));
NOR2XL inst_cellmath__43_1_I652 (.Y(N3876), .A(N3824), .B(N3837));
OAI21X2 inst_cellmath__43_1_I653 (.Y(N3794), .A0(N3811), .A1(N3802), .B0(N3787));
NOR2X2 inst_cellmath__43_1_I654 (.Y(N3817), .A(N3811), .B(N3824));
INVXL inst_cellmath__43_1_I8453 (.Y(N3873), .A(N3806));
AOI21XL inst_cellmath__43_1_I656 (.Y(N3826), .A0(N3876), .A1(N3873), .B0(N3851));
XOR2XL inst_cellmath__43_1_I660 (.Y(inst_cellmath__44[3]), .A(N3791), .B(N3797));
XNOR2X1 inst_cellmath__43_1_I661 (.Y(inst_cellmath__44[5]), .A(N3826), .B(N3829));
AOI21X4 inst_cellmath__43_1_I8454 (.Y(N3870), .A0(N3817), .A1(N3807), .B0(N3794));
XNOR2X1 inst_cellmath__43_1_I662 (.Y(inst_cellmath__44[7]), .A(N3870), .B(N3858));
XNOR2X1 inst_cellmath__43_1_I663 (.Y(N3885), .A(N3835), .B(N3832));
XNOR2XL inst_cellmath__43_1_I664 (.Y(N3860), .A(N3815), .B(N3832));
MX2XL inst_cellmath__43_1_I665 (.Y(inst_cellmath__44[2]), .A(N3860), .B(N3885), .S0(N3873));
XNOR2X1 inst_cellmath__43_1_I666 (.Y(N3847), .A(N3823), .B(N3863));
XNOR2X1 inst_cellmath__43_1_I667 (.Y(N3825), .A(N3801), .B(N3863));
MX2XL inst_cellmath__43_1_I668 (.Y(inst_cellmath__44[4]), .A(N3825), .B(N3847), .S0(N3791));
XNOR2X1 inst_cellmath__43_1_I669 (.Y(N3812), .A(N3810), .B(N3792));
XNOR2X1 inst_cellmath__43_1_I670 (.Y(N3788), .A(N3786), .B(N3792));
MX2XL inst_cellmath__43_1_I671 (.Y(inst_cellmath__44[6]), .A(N3812), .B(N3788), .S0(N3826));
INVXL inst_cellmath__43_1_I8449 (.Y(N14232), .A(N3835));
NOR2XL inst_cellmath__43_1_I8450 (.Y(N14222), .A(N14232), .B(N3815));
NAND2XL node_cs_const1_cs_ii_A_I8756 (.Y(N14623), .A(N500), .B(b_exp[0]));
XOR2XL node_cs_const1_cs_ii_A_I8757 (.Y(N14225), .A(N14222), .B(N14623));
XOR2XL inst_cellmath__43_1_I8455 (.Y(N14214), .A(N3806), .B(N14222));
MXI2X1 inst_cellmath__43_1_I8456 (.Y(N14209), .A(N3798), .B(N3879), .S0(N3870));
INVX1 inst_cellmath__43_1_I8457 (.Y(N4474), .A(N14209));
MXI2X1 inst_cellmath__43_1_I8458 (.Y(N8716), .A(N14225), .B(N14214), .S0(N14209));
INVX2 inst_cellmath__48__10__I3309 (.Y(N8758), .A(N8754));
INVX1 inst_cellmath__48__10__I3307 (.Y(N8756), .A(N8754));
INVX1 inst_cellmath__48__10__I3306 (.Y(N8755), .A(N8754));
MX2XL inst_cellmath__48__10__I677 (.Y(inst_cellmath__48[1]), .A(b_man[0]), .B(a_man[0]), .S0(N8758));
MX2XL inst_cellmath__48__10__I678 (.Y(inst_cellmath__48[2]), .A(b_man[1]), .B(a_man[1]), .S0(N8758));
MX2XL inst_cellmath__48__10__I679 (.Y(inst_cellmath__48[3]), .A(b_man[2]), .B(a_man[2]), .S0(N8758));
MX2XL inst_cellmath__48__10__I681 (.Y(inst_cellmath__48[4]), .A(b_man[3]), .B(a_man[3]), .S0(N8755));
MX2XL inst_cellmath__48__10__I682 (.Y(inst_cellmath__48[5]), .A(b_man[4]), .B(a_man[4]), .S0(N8755));
MX2XL inst_cellmath__48__10__I683 (.Y(inst_cellmath__48[6]), .A(b_man[5]), .B(a_man[5]), .S0(N8755));
MX2XL inst_cellmath__48__10__I684 (.Y(inst_cellmath__48[7]), .A(b_man[6]), .B(a_man[6]), .S0(N8755));
MX2XL inst_cellmath__48__10__I686 (.Y(inst_cellmath__48[8]), .A(b_man[7]), .B(a_man[7]), .S0(N8758));
MX2XL inst_cellmath__48__10__I687 (.Y(inst_cellmath__48[9]), .A(b_man[8]), .B(a_man[8]), .S0(N8758));
MX2XL inst_cellmath__48__10__I688 (.Y(inst_cellmath__48[10]), .A(b_man[9]), .B(a_man[9]), .S0(N8758));
MX2XL inst_cellmath__48__10__I689 (.Y(inst_cellmath__48[11]), .A(b_man[10]), .B(a_man[10]), .S0(N8758));
MX2XL inst_cellmath__48__10__I691 (.Y(inst_cellmath__48[12]), .A(b_man[11]), .B(a_man[11]), .S0(N8756));
MX2XL inst_cellmath__48__10__I692 (.Y(inst_cellmath__48[13]), .A(b_man[12]), .B(a_man[12]), .S0(N8756));
MX2XL inst_cellmath__48__10__I693 (.Y(inst_cellmath__48[14]), .A(b_man[13]), .B(a_man[13]), .S0(N8758));
MX2XL inst_cellmath__48__10__I694 (.Y(inst_cellmath__48[15]), .A(b_man[14]), .B(a_man[14]), .S0(N8758));
MX2XL inst_cellmath__48__10__I696 (.Y(inst_cellmath__48[16]), .A(b_man[15]), .B(a_man[15]), .S0(N4022));
MX2XL inst_cellmath__48__10__I697 (.Y(inst_cellmath__48[17]), .A(b_man[16]), .B(a_man[16]), .S0(N8755));
MX2XL inst_cellmath__48__10__I698 (.Y(inst_cellmath__48[18]), .A(b_man[17]), .B(a_man[17]), .S0(N4022));
MX2XL inst_cellmath__48__10__I699 (.Y(inst_cellmath__48[19]), .A(b_man[18]), .B(a_man[18]), .S0(N8756));
MX2XL inst_cellmath__48__10__I701 (.Y(inst_cellmath__48[20]), .A(b_man[19]), .B(a_man[19]), .S0(N4022));
MX2XL inst_cellmath__48__10__I702 (.Y(inst_cellmath__48[21]), .A(b_man[20]), .B(a_man[20]), .S0(N8756));
MX2XL inst_cellmath__48__10__I703 (.Y(inst_cellmath__48[22]), .A(b_man[21]), .B(a_man[21]), .S0(N4022));
MX2XL inst_cellmath__48__10__I704 (.Y(inst_cellmath__48[23]), .A(b_man[22]), .B(a_man[22]), .S0(N8756));
INVXL cynw_cm_float_add2_I585 (.Y(N3782), .A(N500));
NOR2XL inst_cellmath__28__5__I705 (.Y(N4090), .A(N3782), .B(a_exp[1]));
NOR2XL inst_cellmath__28__5__I706 (.Y(N4094), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL inst_cellmath__28__5__I707 (.Y(N4097), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL inst_cellmath__28__5__I708 (.Y(N4085), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL inst_cellmath__28__5__I3373 (.Y(inst_cellmath__28), .A(N4094), .B(N4097), .C(N4085), .D(N4090));
NOR2XL inst_cellmath__31__7__I712 (.Y(N4112), .A(b_exp[0]), .B(b_exp[1]));
NOR2XL inst_cellmath__31__7__I713 (.Y(N4116), .A(b_exp[7]), .B(b_exp[6]));
NOR2XL inst_cellmath__31__7__I714 (.Y(N4119), .A(b_exp[5]), .B(b_exp[4]));
NOR2XL inst_cellmath__31__7__I715 (.Y(N4107), .A(b_exp[3]), .B(b_exp[2]));
NAND4XL inst_cellmath__31__7__I3374 (.Y(inst_cellmath__31), .A(N4112), .B(N4116), .C(N4119), .D(N4107));
INVX1 inst_cellmath__38__13__I3320 (.Y(N4170), .A(N517));
MXI2XL inst_cellmath__38__13__I725 (.Y(N575), .A(a_man[0]), .B(b_man[0]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I726 (.Y(N576), .A(a_man[1]), .B(b_man[1]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I727 (.Y(N577), .A(a_man[2]), .B(b_man[2]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I728 (.Y(N578), .A(a_man[3]), .B(b_man[3]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I729 (.Y(N579), .A(a_man[4]), .B(b_man[4]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I730 (.Y(N580), .A(a_man[5]), .B(b_man[5]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I731 (.Y(N581), .A(a_man[6]), .B(b_man[6]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I732 (.Y(N582), .A(a_man[7]), .B(b_man[7]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I733 (.Y(N583), .A(a_man[8]), .B(b_man[8]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I734 (.Y(N584), .A(a_man[9]), .B(b_man[9]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I735 (.Y(N585), .A(a_man[10]), .B(b_man[10]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I736 (.Y(N586), .A(a_man[11]), .B(b_man[11]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I737 (.Y(N587), .A(a_man[12]), .B(b_man[12]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I738 (.Y(N588), .A(a_man[13]), .B(b_man[13]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I739 (.Y(N589), .A(a_man[14]), .B(b_man[14]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I740 (.Y(N590), .A(a_man[15]), .B(b_man[15]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I741 (.Y(N591), .A(a_man[16]), .B(b_man[16]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I742 (.Y(N592), .A(a_man[17]), .B(b_man[17]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I743 (.Y(N593), .A(a_man[18]), .B(b_man[18]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I744 (.Y(N594), .A(a_man[19]), .B(b_man[19]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I745 (.Y(N595), .A(a_man[20]), .B(b_man[20]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I746 (.Y(N596), .A(a_man[21]), .B(b_man[21]), .S0(N4170));
MXI2XL inst_cellmath__38__13__I747 (.Y(N597), .A(a_man[22]), .B(b_man[22]), .S0(N4170));
AND4XL inst_cellmath__30_0_I8647 (.Y(N4237), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[7]), .D(b_exp[6]));
AND4XL inst_cellmath__30_0_I8648 (.Y(N4241), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND2XL inst_cellmath__30_0_I754 (.Y(inst_cellmath__30), .A(N4237), .B(N4241));
NOR2XL inst_cellmath__32__8__I760 (.Y(N4291), .A(b_man[14]), .B(b_man[13]));
NOR2XL inst_cellmath__32__8__I761 (.Y(N4301), .A(b_man[12]), .B(b_man[11]));
OR4X1 inst_cellmath__32__8__I8649 (.Y(N4279), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__32__8__I8650 (.Y(N4289), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__32__8__I8651 (.Y(N4262), .A(b_man[10]), .B(b_man[8]), .C(b_man[9]), .D(b_man[7]));
OR4X1 inst_cellmath__32__8__I8652 (.Y(N4272), .A(b_man[6]), .B(b_man[4]), .C(b_man[5]), .D(b_man[3]));
NOR4X1 inst_cellmath__32__8__I3322 (.Y(N4283), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N4279));
NAND3XL inst_cellmath__32__8__I3456 (.Y(N8764), .A(N4291), .B(N4301), .C(N4283));
OR4X1 inst_cellmath__32__8__I8653 (.Y(inst_cellmath__32), .A(N4272), .B(N4262), .C(N4289), .D(N8764));
NOR2XL cynw_cm_float_add2_I778 (.Y(inst_cellmath__24), .A(inst_cellmath__30), .B(inst_cellmath__32));
XOR2X4 cynw_cm_float_add2_I779 (.Y(inst_cellmath__55[0]), .A(a_sign), .B(b_sign));
NAND2XL inst_cellmath__27_0_I780 (.Y(N4338), .A(N3782), .B(a_exp[1]));
AND4XL inst_cellmath__27_0_I8655 (.Y(N4340), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND4BXL inst_cellmath__27_0_I8657 (.Y(inst_cellmath__27), .AN(N4338), .B(a_exp[7]), .C(N4340), .D(a_exp[6]));
NOR2XL inst_cellmath__29__6__I792 (.Y(N4390), .A(a_man[14]), .B(a_man[13]));
NOR2XL inst_cellmath__29__6__I793 (.Y(N4400), .A(a_man[12]), .B(a_man[11]));
OR4X1 inst_cellmath__29__6__I8658 (.Y(N4378), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__29__6__I8659 (.Y(N4388), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__29__6__I8660 (.Y(N4361), .A(a_man[10]), .B(a_man[8]), .C(a_man[9]), .D(a_man[7]));
OR4X1 inst_cellmath__29__6__I8661 (.Y(N4371), .A(a_man[6]), .B(a_man[4]), .C(a_man[5]), .D(a_man[3]));
NOR4X1 inst_cellmath__29__6__I3325 (.Y(N4382), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N4378));
NAND3XL inst_cellmath__29__6__I3458 (.Y(N8772), .A(N4390), .B(N4400), .C(N4382));
OR4X1 inst_cellmath__29__6__I8662 (.Y(inst_cellmath__29), .A(N4371), .B(N4361), .C(N4388), .D(N8772));
NOR2XL cynw_cm_float_add2_I810 (.Y(inst_cellmath__21), .A(inst_cellmath__27), .B(inst_cellmath__29));
NAND2BXL cynw_cm_float_add2_I3328 (.Y(inst_cellmath__20), .AN(inst_cellmath__27), .B(inst_cellmath__29));
NAND2BXL cynw_cm_float_add2_I3329 (.Y(inst_cellmath__23), .AN(inst_cellmath__30), .B(inst_cellmath__32));
NAND2XL cynw_cm_float_add2_I817 (.Y(N4450), .A(inst_cellmath__23), .B(inst_cellmath__20));
MXI2X6 cynw_cm_float_add2_I3260 (.Y(inst_cellmath__47[2]), .A(inst_cellmath__44[2]), .B(N511), .S0(N4474));
MX2XL cynw_cm_float_add2_I833 (.Y(inst_cellmath__47[3]), .A(inst_cellmath__44[3]), .B(N512), .S0(N4474));
MX2XL cynw_cm_float_add2_I3262 (.Y(inst_cellmath__47[5]), .A(inst_cellmath__44[5]), .B(N514), .S0(N4474));
MXI2XL cynw_cm_float_add2_I3263 (.Y(inst_cellmath__47[6]), .A(inst_cellmath__44[6]), .B(N515), .S0(N4474));
MX2XL cynw_cm_float_add2_I3264 (.Y(inst_cellmath__47[7]), .A(inst_cellmath__44[7]), .B(N516), .S0(N4474));
CLKBUFX6 inst_cellmath__49_0_I3265 (.Y(N4633), .A(N8716));
NOR2BXL inst_cellmath__49_0_I839 (.Y(N4651), .AN(inst_cellmath__48[2]), .B(N4633));
MX2XL inst_cellmath__49_0_I840 (.Y(N4559), .A(inst_cellmath__48[3]), .B(inst_cellmath__48[1]), .S0(N4633));
MX2XL inst_cellmath__49_0_I841 (.Y(N4594), .A(inst_cellmath__48[4]), .B(inst_cellmath__48[2]), .S0(N4633));
MX2XL inst_cellmath__49_0_I842 (.Y(N4628), .A(inst_cellmath__48[5]), .B(inst_cellmath__48[3]), .S0(N4633));
MX2XL inst_cellmath__49_0_I843 (.Y(N4666), .A(inst_cellmath__48[6]), .B(inst_cellmath__48[4]), .S0(N4633));
MXI2XL mx2a_A_I8758 (.Y(N14630), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[5]), .S0(N4633));
INVXL mx2a_A_I8759 (.Y(N4540), .A(N14630));
MX2XL inst_cellmath__49_0_I845 (.Y(N4575), .A(inst_cellmath__48[8]), .B(inst_cellmath__48[6]), .S0(N4633));
MX2XL inst_cellmath__49_0_I846 (.Y(N4607), .A(inst_cellmath__48[9]), .B(inst_cellmath__48[7]), .S0(N4633));
MX2XL inst_cellmath__49_0_I847 (.Y(N4645), .A(inst_cellmath__48[10]), .B(inst_cellmath__48[8]), .S0(N4633));
MX2XL inst_cellmath__49_0_I848 (.Y(N4520), .A(inst_cellmath__48[11]), .B(inst_cellmath__48[9]), .S0(N4633));
MX2XL inst_cellmath__49_0_I849 (.Y(N4554), .A(inst_cellmath__48[12]), .B(inst_cellmath__48[10]), .S0(N4633));
MX2XL inst_cellmath__49_0_I850 (.Y(N4589), .A(inst_cellmath__48[13]), .B(inst_cellmath__48[11]), .S0(N4633));
MX2XL inst_cellmath__49_0_I3429 (.Y(N4622), .A(inst_cellmath__48[14]), .B(inst_cellmath__48[12]), .S0(N4633));
MX2XL inst_cellmath__49_0_I852 (.Y(N4660), .A(inst_cellmath__48[15]), .B(inst_cellmath__48[13]), .S0(N4633));
MX2XL inst_cellmath__49_0_I853 (.Y(N4534), .A(inst_cellmath__48[16]), .B(inst_cellmath__48[14]), .S0(N4633));
MX2XL inst_cellmath__49_0_I854 (.Y(N4568), .A(inst_cellmath__48[17]), .B(inst_cellmath__48[15]), .S0(N4633));
MX2XL inst_cellmath__49_0_I855 (.Y(N4602), .A(inst_cellmath__48[18]), .B(inst_cellmath__48[16]), .S0(N4633));
MX2XL inst_cellmath__49_0_I856 (.Y(N4638), .A(inst_cellmath__48[19]), .B(inst_cellmath__48[17]), .S0(N4633));
MX2XL inst_cellmath__49_0_I857 (.Y(N4514), .A(inst_cellmath__48[20]), .B(inst_cellmath__48[18]), .S0(N4633));
MX2XL inst_cellmath__49_0_I858 (.Y(N4548), .A(inst_cellmath__48[21]), .B(inst_cellmath__48[19]), .S0(N4633));
MX2XL inst_cellmath__49_0_I859 (.Y(N4584), .A(inst_cellmath__48[22]), .B(inst_cellmath__48[20]), .S0(N4633));
MX2XL inst_cellmath__49_0_I860 (.Y(N4615), .A(inst_cellmath__48[23]), .B(inst_cellmath__48[21]), .S0(N4633));
NAND2BXL inst_cellmath__49_0_I861 (.Y(N4655), .AN(inst_cellmath__48[22]), .B(N4633));
AND2XL inst_cellmath__49_0_I862 (.Y(N4563), .A(N4633), .B(inst_cellmath__48[23]));
INVX6 inst_cellmath__49_0_I863 (.Y(N4578), .A(inst_cellmath__47[2]));
AOI22XL inst_cellmath__49_0_I864 (.Y(N4626), .A0(N4666), .A1(inst_cellmath__47[2]), .B0(N4651), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I865 (.Y(N4665), .A0(inst_cellmath__47[2]), .A1(N4540), .B0(N4559), .B1(N4578));
AOI22XL inst_cellmath__49_0_I866 (.Y(N4538), .A0(inst_cellmath__47[2]), .A1(N4575), .B0(N4594), .B1(N4578));
AOI22XL inst_cellmath__49_0_I867 (.Y(N4574), .A0(inst_cellmath__47[2]), .A1(N4607), .B0(N4628), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I868 (.Y(N4605), .A0(inst_cellmath__47[2]), .A1(N4645), .B0(N4666), .B1(N4578));
AOI22XL inst_cellmath__49_0_I869 (.Y(N4644), .A0(inst_cellmath__47[2]), .A1(N4520), .B0(N4540), .B1(N4578));
AOI22XL inst_cellmath__49_0_I870 (.Y(N4519), .A0(inst_cellmath__47[2]), .A1(N4554), .B0(N4575), .B1(N4578));
AOI22XL inst_cellmath__49_0_I871 (.Y(N4553), .A0(inst_cellmath__47[2]), .A1(N4589), .B0(N4607), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I872 (.Y(N4588), .A0(inst_cellmath__47[2]), .A1(N4622), .B0(N4578), .B1(N4645));
AOI22XL inst_cellmath__49_0_I873 (.Y(N4621), .A0(inst_cellmath__47[2]), .A1(N4660), .B0(N4520), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I874 (.Y(N4659), .A0(N4534), .A1(inst_cellmath__47[2]), .B0(N4578), .B1(N4554));
AOI22XL inst_cellmath__49_0_I875 (.Y(N4533), .A0(inst_cellmath__47[2]), .A1(N4568), .B0(N4589), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I876 (.Y(N4567), .A0(inst_cellmath__47[2]), .A1(N4602), .B0(N4578), .B1(N4622));
AOI22X1 inst_cellmath__49_0_I877 (.Y(N4601), .A0(inst_cellmath__47[2]), .A1(N4638), .B0(N4578), .B1(N4660));
AOI22X1 inst_cellmath__49_0_I878 (.Y(N4637), .A0(inst_cellmath__47[2]), .A1(N4514), .B0(N4578), .B1(N4534));
AOI22X1 inst_cellmath__49_0_I879 (.Y(N4513), .A0(N4548), .A1(inst_cellmath__47[2]), .B0(N4568), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I880 (.Y(N4547), .A0(inst_cellmath__47[2]), .A1(N4584), .B0(N4602), .B1(N4578));
AOI22X1 inst_cellmath__49_0_I881 (.Y(N4583), .A0(N4615), .A1(inst_cellmath__47[2]), .B0(N4578), .B1(N4638));
AOI22X1 inst_cellmath__49_0_I882 (.Y(N4614), .A0(N4655), .A1(inst_cellmath__47[2]), .B0(N4514), .B1(N4578));
AOI22XL inst_cellmath__49_0_I883 (.Y(N4654), .A0(inst_cellmath__47[2]), .A1(N4563), .B0(N4548), .B1(N4578));
AOI22XL inst_cellmath__49_0_I884 (.Y(N4527), .A0(inst_cellmath__47[2]), .A1(N4633), .B0(N4584), .B1(N4578));
NAND2XL inst_cellmath__49_0_I885 (.Y(N4561), .A(N4578), .B(N4615));
NAND2XL inst_cellmath__49_0_I886 (.Y(N4631), .A(N4655), .B(N4578));
NAND2X1 inst_cellmath__49_0_I887 (.Y(N4542), .A(N4563), .B(N4578));
NAND2XL inst_cellmath__49_0_I888 (.Y(N4609), .A(N4633), .B(N4578));
INVX2 inst_cellmath__49_0_I889 (.Y(N4610), .A(inst_cellmath__47[3]));
INVX3 inst_cellmath__49_0_I890 (.Y(N4648), .A(N4610));
AOI22XL inst_cellmath__49_0_I891 (.Y(N4572), .A0(N4610), .A1(N4626), .B0(N4648), .B1(N4588));
AOI22X1 inst_cellmath__49_0_I892 (.Y(N4603), .A0(N4610), .A1(N4665), .B0(N4648), .B1(N4621));
AOI22XL inst_cellmath__49_0_I893 (.Y(N4643), .A0(N4610), .A1(N4538), .B0(N4648), .B1(N4659));
AOI22XL inst_cellmath__49_0_I894 (.Y(N4518), .A0(N4610), .A1(N4574), .B0(N4648), .B1(N4533));
AOI22X1 inst_cellmath__49_0_I895 (.Y(N4552), .A0(N4610), .A1(N4605), .B0(N4648), .B1(N4567));
AOI22X1 inst_cellmath__49_0_I896 (.Y(N4587), .A0(N4610), .A1(N4644), .B0(N4648), .B1(N4601));
AOI22XL inst_cellmath__49_0_I897 (.Y(N4619), .A0(N4610), .A1(N4519), .B0(N4648), .B1(N4637));
AOI22X1 inst_cellmath__49_0_I898 (.Y(N4657), .A0(N4610), .A1(N4553), .B0(N4648), .B1(N4513));
AOI22XL inst_cellmath__49_0_I899 (.Y(N4532), .A0(N4610), .A1(N4588), .B0(N4648), .B1(N4547));
AOI22XL inst_cellmath__49_0_I900 (.Y(N4566), .A0(N4610), .A1(N4621), .B0(N4648), .B1(N4583));
AOI22XL inst_cellmath__49_0_I901 (.Y(N4600), .A0(N4610), .A1(N4659), .B0(N4648), .B1(N4614));
AOI22XL inst_cellmath__49_0_I902 (.Y(N4636), .A0(N4610), .A1(N4533), .B0(N4648), .B1(N4654));
AOI22X1 inst_cellmath__49_0_I903 (.Y(N4511), .A0(N4610), .A1(N4567), .B0(N4648), .B1(N4527));
AOI22X1 inst_cellmath__49_0_I904 (.Y(N4545), .A0(N4610), .A1(N4601), .B0(N4648), .B1(N4561));
AOI22XL inst_cellmath__49_0_I905 (.Y(N4582), .A0(N4610), .A1(N4637), .B0(N4648), .B1(N4631));
AOI22X1 inst_cellmath__49_0_I906 (.Y(N4613), .A0(N4610), .A1(N4513), .B0(N4648), .B1(N4542));
AOI22X1 inst_cellmath__49_0_I907 (.Y(N4653), .A0(N4610), .A1(N4547), .B0(N4648), .B1(N4609));
NOR2X1 inst_cellmath__49_0_I908 (.Y(N4526), .A(N4648), .B(N4583));
NOR2X1 inst_cellmath__49_0_I909 (.Y(N4630), .A(N4648), .B(N4614));
NOR2X1 inst_cellmath__49_0_I910 (.Y(N4577), .A(N4648), .B(N4654));
NOR2X1 inst_cellmath__49_0_I911 (.Y(N4522), .A(N4648), .B(N4527));
NOR2X1 inst_cellmath__49_0_I912 (.Y(N4624), .A(N4648), .B(N4561));
NOR2X1 inst_cellmath__49_0_I913 (.Y(N4570), .A(N4648), .B(N4631));
NOR2X1 inst_cellmath__49_0_I914 (.Y(N4516), .A(N4648), .B(N4542));
NOR2X1 inst_cellmath__49_0_I915 (.Y(N4617), .A(N4648), .B(N4609));
MX2X1 inst_cellmath__49_0_I3266 (.Y(N4556), .A(inst_cellmath__44[4]), .B(N513), .S0(N4474));
INVX1 inst_cellmath__49_0_I917 (.Y(N4592), .A(N4556));
AOI22X1 inst_cellmath__49_0_I918 (.Y(N4528), .A0(N4592), .A1(N4653), .B0(N4556), .B1(N4572));
AOI22X1 inst_cellmath__49_0_I919 (.Y(N4562), .A0(N4592), .A1(N4526), .B0(N4556), .B1(N4603));
AOI22XL inst_cellmath__49_0_I920 (.Y(N4596), .A0(N4592), .A1(N4630), .B0(N4556), .B1(N4643));
AOI22X1 inst_cellmath__49_0_I921 (.Y(N4632), .A0(N4592), .A1(N4577), .B0(N4556), .B1(N4518));
AOI22X1 inst_cellmath__49_0_I922 (.Y(N4668), .A0(N4592), .A1(N4522), .B0(N4556), .B1(N4552));
AOI22X1 inst_cellmath__49_0_I923 (.Y(N4543), .A0(N4592), .A1(N4624), .B0(N4556), .B1(N4587));
AOI22X1 inst_cellmath__49_0_I924 (.Y(N4579), .A0(N4570), .A1(N4592), .B0(N4556), .B1(N4619));
AOI22X1 inst_cellmath__49_0_I925 (.Y(N4611), .A0(N4592), .A1(N4516), .B0(N4556), .B1(N4657));
AOI22X1 inst_cellmath__49_0_I926 (.Y(N4647), .A0(N4592), .A1(N4617), .B0(N4556), .B1(N4532));
NAND2X1 inst_cellmath__49_0_I927 (.Y(N4523), .A(N4556), .B(N4566));
NAND2X1 inst_cellmath__49_0_I928 (.Y(N4591), .A(N4556), .B(N4600));
NAND2XL inst_cellmath__49_0_I929 (.Y(N4663), .A(N4556), .B(N4636));
NAND2X1 inst_cellmath__49_0_I930 (.Y(N4571), .A(N4556), .B(N4511));
NAND2X1 inst_cellmath__49_0_I931 (.Y(N4640), .A(N4556), .B(N4545));
NAND2X1 inst_cellmath__49_0_I932 (.Y(N4550), .A(N4556), .B(N4582));
NAND2XL inst_cellmath__49_0_I933 (.Y(N4618), .A(N4556), .B(N4613));
NAND2XL inst_cellmath__49_0_I934 (.Y(N4530), .A(N4556), .B(N4653));
NAND2XL inst_cellmath__49_0_I935 (.Y(N4597), .A(N4556), .B(N4526));
NAND2XL inst_cellmath__49_0_I936 (.Y(N4509), .A(N4556), .B(N4630));
NAND2XL inst_cellmath__49_0_I937 (.Y(N4580), .A(N4556), .B(N4577));
NAND2XL inst_cellmath__49_0_I938 (.Y(N4650), .A(N4556), .B(N4522));
NAND2XL inst_cellmath__49_0_I939 (.Y(N4558), .A(N4556), .B(N4624));
NAND2XL inst_cellmath__49_0_I940 (.Y(N4627), .A(N4570), .B(N4556));
NAND2XL inst_cellmath__49_0_I941 (.Y(N4539), .A(N4556), .B(N4516));
NAND2XL inst_cellmath__49_0_I942 (.Y(N4606), .A(N4556), .B(N4617));
CLKXOR2X2 inst_cellmath__49_0_I8293 (.Y(N4662), .A(b_exp[0]), .B(N500));
INVX1 inst_cellmath__49_0_I944 (.Y(N4536), .A(N4662));
AOI22XL inst_cellmath__49_0_I945 (.Y(inst_cellmath__49[0]), .A0(N4662), .A1(N4528), .B0(N4562), .B1(N4536));
AOI22XL inst_cellmath__49_0_I946 (.Y(inst_cellmath__49[1]), .A0(N4662), .A1(N4562), .B0(N4596), .B1(N4536));
AOI22XL inst_cellmath__49_0_I947 (.Y(inst_cellmath__49[2]), .A0(N4596), .A1(N4662), .B0(N4536), .B1(N4632));
AOI22XL inst_cellmath__49_0_I948 (.Y(inst_cellmath__49[3]), .A0(N4662), .A1(N4632), .B0(N4536), .B1(N4668));
AOI22XL inst_cellmath__49_0_I949 (.Y(inst_cellmath__49[4]), .A0(N4662), .A1(N4668), .B0(N4536), .B1(N4543));
AOI22X1 inst_cellmath__49_0_I950 (.Y(inst_cellmath__49[5]), .A0(N4662), .A1(N4543), .B0(N4579), .B1(N4536));
AOI22XL inst_cellmath__49_0_I951 (.Y(inst_cellmath__49[6]), .A0(N4662), .A1(N4579), .B0(N4536), .B1(N4611));
AOI22XL inst_cellmath__49_0_I952 (.Y(inst_cellmath__49[7]), .A0(N4662), .A1(N4611), .B0(N4536), .B1(N4647));
AOI22X1 inst_cellmath__49_0_I953 (.Y(inst_cellmath__49[8]), .A0(N4662), .A1(N4647), .B0(N4536), .B1(N4523));
AOI22XL inst_cellmath__49_0_I954 (.Y(inst_cellmath__49[9]), .A0(N4662), .A1(N4523), .B0(N4591), .B1(N4536));
AOI22XL inst_cellmath__49_0_I955 (.Y(inst_cellmath__49[10]), .A0(N4662), .A1(N4591), .B0(N4663), .B1(N4536));
AOI22XL inst_cellmath__49_0_I956 (.Y(inst_cellmath__49[11]), .A0(N4662), .A1(N4663), .B0(N4536), .B1(N4571));
AOI22X1 inst_cellmath__49_0_I957 (.Y(inst_cellmath__49[12]), .A0(N4662), .A1(N4571), .B0(N4536), .B1(N4640));
AOI22X1 inst_cellmath__49_0_I958 (.Y(inst_cellmath__49[13]), .A0(N4662), .A1(N4640), .B0(N4550), .B1(N4536));
AOI22XL inst_cellmath__49_0_I959 (.Y(inst_cellmath__49[14]), .A0(N4662), .A1(N4550), .B0(N4536), .B1(N4618));
AOI22XL inst_cellmath__49_0_I960 (.Y(inst_cellmath__49[15]), .A0(N4662), .A1(N4618), .B0(N4536), .B1(N4530));
AOI22X1 inst_cellmath__49_0_I961 (.Y(inst_cellmath__49[16]), .A0(N4662), .A1(N4530), .B0(N4597), .B1(N4536));
AOI22XL inst_cellmath__49_0_I962 (.Y(inst_cellmath__49[17]), .A0(N4536), .A1(N4509), .B0(N4662), .B1(N4597));
AOI22XL inst_cellmath__49_0_I963 (.Y(inst_cellmath__49[18]), .A0(N4662), .A1(N4509), .B0(N4536), .B1(N4580));
AOI22XL inst_cellmath__49_0_I964 (.Y(inst_cellmath__49[19]), .A0(N4662), .A1(N4580), .B0(N4536), .B1(N4650));
AOI22XL inst_cellmath__49_0_I965 (.Y(inst_cellmath__49[20]), .A0(N4662), .A1(N4650), .B0(N4558), .B1(N4536));
AOI22XL inst_cellmath__49_0_I966 (.Y(inst_cellmath__49[21]), .A0(N4662), .A1(N4558), .B0(N4627), .B1(N4536));
AOI22XL inst_cellmath__49_0_I967 (.Y(inst_cellmath__49[22]), .A0(N4627), .A1(N4662), .B0(N4536), .B1(N4539));
AOI22XL inst_cellmath__49_0_I968 (.Y(inst_cellmath__49[23]), .A0(N4662), .A1(N4539), .B0(N4536), .B1(N4606));
NOR3XL cynw_cm_float_add2_I970 (.Y(N4836), .A(inst_cellmath__47[6]), .B(inst_cellmath__47[5]), .C(inst_cellmath__47[7]));
AND2XL inst_cellmath__39_2mx_I996 (.Y(N4897), .A(inst_cellmath__31), .B(inst_cellmath__28));
AND2X1 cynw_cm_float_add2_I971 (.Y(N522), .A(N4897), .B(N4836));
AND2X1 inst_cellmath__39_2mx_I997 (.Y(inst_cellmath__39[0]), .A(inst_cellmath__49[0]), .B(N522));
AND2XL inst_cellmath__39_2mx_I998 (.Y(inst_cellmath__39[1]), .A(N522), .B(inst_cellmath__49[1]));
AND2X1 inst_cellmath__39_2mx_I999 (.Y(inst_cellmath__39[2]), .A(inst_cellmath__49[2]), .B(N522));
AND2X1 inst_cellmath__39_2mx_I1000 (.Y(inst_cellmath__39[3]), .A(inst_cellmath__49[3]), .B(N522));
CLKAND2X2 inst_cellmath__39_2mx_I1001 (.Y(inst_cellmath__39[4]), .A(N522), .B(inst_cellmath__49[4]));
CLKAND2X2 inst_cellmath__39_2mx_I1002 (.Y(inst_cellmath__39[5]), .A(N522), .B(inst_cellmath__49[5]));
AND2X1 inst_cellmath__39_2mx_I1003 (.Y(inst_cellmath__39[6]), .A(inst_cellmath__49[6]), .B(N522));
AND2X1 inst_cellmath__39_2mx_I1004 (.Y(inst_cellmath__39[7]), .A(inst_cellmath__49[7]), .B(N522));
CLKAND2X3 inst_cellmath__39_2mx_I1005 (.Y(inst_cellmath__39[8]), .A(N522), .B(inst_cellmath__49[8]));
CLKAND2X2 inst_cellmath__39_2mx_I1006 (.Y(inst_cellmath__39[9]), .A(N522), .B(inst_cellmath__49[9]));
CLKAND2X2 inst_cellmath__39_2mx_I1007 (.Y(inst_cellmath__39[10]), .A(N522), .B(inst_cellmath__49[10]));
CLKAND2X2 inst_cellmath__39_2mx_I1008 (.Y(inst_cellmath__39[11]), .A(N522), .B(inst_cellmath__49[11]));
CLKAND2X2 inst_cellmath__39_2mx_I1009 (.Y(inst_cellmath__39[12]), .A(N522), .B(inst_cellmath__49[12]));
AND2X1 inst_cellmath__39_2mx_I1010 (.Y(inst_cellmath__39[13]), .A(inst_cellmath__49[13]), .B(N522));
AND2X1 inst_cellmath__39_2mx_I1011 (.Y(inst_cellmath__39[14]), .A(inst_cellmath__49[14]), .B(N522));
CLKAND2X2 inst_cellmath__39_2mx_I1012 (.Y(inst_cellmath__39[15]), .A(N522), .B(inst_cellmath__49[15]));
CLKAND2X2 inst_cellmath__39_2mx_I1013 (.Y(inst_cellmath__39[16]), .A(N522), .B(inst_cellmath__49[16]));
AND2XL inst_cellmath__39_2mx_I1014 (.Y(inst_cellmath__39[17]), .A(N522), .B(inst_cellmath__49[17]));
AND2XL inst_cellmath__39_2mx_I1015 (.Y(inst_cellmath__39[18]), .A(N522), .B(inst_cellmath__49[18]));
CLKAND2X2 inst_cellmath__39_2mx_I1016 (.Y(inst_cellmath__39[19]), .A(N522), .B(inst_cellmath__49[19]));
CLKAND2X2 inst_cellmath__39_2mx_I1017 (.Y(inst_cellmath__39[20]), .A(N522), .B(inst_cellmath__49[20]));
AND2XL inst_cellmath__39_2mx_I1018 (.Y(inst_cellmath__39[21]), .A(N522), .B(inst_cellmath__49[21]));
AND3XL inst_cellmath__39_2mx_I3335 (.Y(inst_cellmath__39[22]), .A(N4836), .B(N4897), .C(inst_cellmath__49[22]));
XNOR2X1 inst_cellmath__39_2mx_I8415 (.Y(N14173), .A(N597), .B(inst_cellmath__55[0]));
INVX2 inst_cellmath__39_2mx_I8416 (.Y(inst_cellmath__55[24]), .A(inst_cellmath__55[0]));
AND3XL inst_cellmath__39_2mx_I8417 (.Y(N14169), .A(N4836), .B(N4897), .C(inst_cellmath__49[23]));
NAND2X1 inst_cellmath__39_2mx_I8419 (.Y(N5326), .A(N14173), .B(N14169));
NOR4BBX1 inst_cellmath__39_2mx_I8420 (.Y(N14181), .AN(N4836), .BN(N4897), .C(N4536), .D(N4606));
XNOR2X1 inst_cellmath__55_2mx_I1027 (.Y(inst_cellmath__55[6]), .A(inst_cellmath__55[0]), .B(N580));
NAND2X2 inst_cellmath__57__22__I1058 (.Y(N5152), .A(inst_cellmath__55[6]), .B(inst_cellmath__39[6]));
XNOR2X1 inst_cellmath__55_2mx_I1026 (.Y(inst_cellmath__55[5]), .A(N579), .B(inst_cellmath__55[0]));
NAND2X2 inst_cellmath__57__22__I1056 (.Y(N5384), .A(inst_cellmath__55[5]), .B(inst_cellmath__39[5]));
NAND2XL inst_cellmath__57__22__I1269 (.Y(N5318), .A(N5152), .B(N5384));
XNOR2X2 inst_cellmath__55_2mx_I1025 (.Y(inst_cellmath__55[4]), .A(N578), .B(inst_cellmath__55[0]));
NAND2X2 inst_cellmath__57__22__I1054 (.Y(N5211), .A(inst_cellmath__55[4]), .B(inst_cellmath__39[4]));
XNOR2X1 inst_cellmath__55_2mx_I1024 (.Y(inst_cellmath__55[3]), .A(N577), .B(inst_cellmath__55[0]));
NAND2X2 inst_cellmath__57__22__I1052 (.Y(N5437), .A(inst_cellmath__55[3]), .B(inst_cellmath__39[3]));
NAND2XL inst_cellmath__57__22__I1266 (.Y(N5369), .A(N5437), .B(N5211));
NOR2X1 inst_cellmath__57__22__I1271 (.Y(N5217), .A(N5318), .B(N5369));
XNOR2X1 inst_cellmath__55_2mx_I1023 (.Y(inst_cellmath__55[2]), .A(inst_cellmath__55[0]), .B(N576));
NAND2X2 inst_cellmath__57__22__I1050 (.Y(N5254), .A(inst_cellmath__55[2]), .B(inst_cellmath__39[2]));
XNOR2X1 inst_cellmath__55_2mx_I1022 (.Y(inst_cellmath__55[1]), .A(N575), .B(inst_cellmath__55[0]));
NAND2X1 inst_cellmath__57__22__I1048 (.Y(N5075), .A(inst_cellmath__55[1]), .B(inst_cellmath__39[1]));
NAND2XL inst_cellmath__57__22__I1263 (.Y(N5114), .A(N5254), .B(N5075));
NAND2X2 inst_cellmath__57__22__I1046 (.Y(N5311), .A(inst_cellmath__55[0]), .B(inst_cellmath__39[0]));
NOR2XL inst_cellmath__57__22__I1258 (.Y(N5350), .A(inst_cellmath__55[0]), .B(inst_cellmath__39[0]));
AOI21X1 inst_cellmath__57__22__I1260 (.Y(N5076), .A0(inst_cellmath__55[24]), .A1(N5311), .B0(N5350));
NOR2X1 inst_cellmath__57__22__I1047 (.Y(N5400), .A(inst_cellmath__55[1]), .B(inst_cellmath__39[1]));
NOR2X2 inst_cellmath__57__22__I1049 (.Y(N5169), .A(inst_cellmath__55[2]), .B(inst_cellmath__39[2]));
AOI21XL inst_cellmath__57__22__I1262 (.Y(N5439), .A0(N5254), .A1(N5400), .B0(N5169));
OAI21X1 inst_cellmath__57__22__I1264 (.Y(N5333), .A0(N5114), .A1(N5076), .B0(N5439));
NOR2X1 inst_cellmath__57__22__I1051 (.Y(N5348), .A(inst_cellmath__55[3]), .B(inst_cellmath__39[3]));
NOR2X4 inst_cellmath__57__22__I1053 (.Y(N5115), .A(inst_cellmath__55[4]), .B(inst_cellmath__39[4]));
AOI21X1 inst_cellmath__57__22__I1265 (.Y(N5273), .A0(N5211), .A1(N5348), .B0(N5115));
NOR2X1 inst_cellmath__57__22__I1055 (.Y(N5291), .A(inst_cellmath__55[5]), .B(inst_cellmath__39[5]));
NOR2X1 inst_cellmath__57__22__I1057 (.Y(N5059), .A(inst_cellmath__55[6]), .B(inst_cellmath__39[6]));
AOI21XL inst_cellmath__57__22__I1268 (.Y(N5229), .A0(N5152), .A1(N5291), .B0(N5059));
OAI21X1 inst_cellmath__57__22__I1270 (.Y(N5119), .A0(N5318), .A1(N5273), .B0(N5229));
AOI21X2 inst_cellmath__39_2mx_I8427 (.Y(N5358), .A0(N5217), .A1(N5333), .B0(N5119));
XNOR2X1 inst_cellmath__55_2mx_I1035 (.Y(inst_cellmath__55[14]), .A(N588), .B(inst_cellmath__55[0]));
XNOR2X1 inst_cellmath__55_2mx_I1034 (.Y(inst_cellmath__55[13]), .A(inst_cellmath__55[0]), .B(N587));
XNOR2X1 inst_cellmath__55_2mx_I1033 (.Y(inst_cellmath__55[12]), .A(inst_cellmath__55[0]), .B(N586));
XNOR2X1 inst_cellmath__55_2mx_I1032 (.Y(inst_cellmath__55[11]), .A(inst_cellmath__55[0]), .B(N585));
XNOR2X1 inst_cellmath__55_2mx_I1031 (.Y(inst_cellmath__55[10]), .A(inst_cellmath__55[0]), .B(N584));
XNOR2X1 inst_cellmath__55_2mx_I1030 (.Y(inst_cellmath__55[9]), .A(inst_cellmath__55[0]), .B(N583));
XNOR2X1 inst_cellmath__55_2mx_I1029 (.Y(inst_cellmath__55[8]), .A(inst_cellmath__55[0]), .B(N582));
XNOR2X1 inst_cellmath__55_2mx_I1028 (.Y(inst_cellmath__55[7]), .A(N581), .B(inst_cellmath__55[0]));
NOR2X1 inst_cellmath__39_2mx_I8563 (.Y(N5243), .A(inst_cellmath__55[7]), .B(inst_cellmath__39[7]));
NOR2X4 inst_cellmath__39_2mx_I8564 (.Y(N5420), .A(inst_cellmath__55[8]), .B(inst_cellmath__39[8]));
NAND2X4 inst_cellmath__39_2mx_I8565 (.Y(N5095), .A(inst_cellmath__55[8]), .B(inst_cellmath__39[8]));
NOR2X2 inst_cellmath__39_2mx_I8566 (.Y(N5193), .A(inst_cellmath__55[9]), .B(inst_cellmath__39[9]));
NAND2X4 inst_cellmath__39_2mx_I8567 (.Y(N5272), .A(inst_cellmath__55[9]), .B(inst_cellmath__39[9]));
NOR2X2 inst_cellmath__39_2mx_I8568 (.Y(N5370), .A(inst_cellmath__55[10]), .B(inst_cellmath__39[10]));
NAND2X4 inst_cellmath__39_2mx_I8569 (.Y(N5046), .A(inst_cellmath__55[10]), .B(inst_cellmath__39[10]));
NOR2X1 inst_cellmath__39_2mx_I8570 (.Y(N5133), .A(inst_cellmath__55[11]), .B(inst_cellmath__39[11]));
NAND2X2 inst_cellmath__39_2mx_I8571 (.Y(N5230), .A(inst_cellmath__55[11]), .B(inst_cellmath__39[11]));
NOR2X1 inst_cellmath__39_2mx_I8572 (.Y(N5317), .A(inst_cellmath__55[12]), .B(inst_cellmath__39[12]));
NAND2X2 inst_cellmath__39_2mx_I8573 (.Y(N5406), .A(inst_cellmath__55[12]), .B(inst_cellmath__39[12]));
NOR2X1 inst_cellmath__39_2mx_I8574 (.Y(N5080), .A(inst_cellmath__55[13]), .B(inst_cellmath__39[13]));
NAND2X2 inst_cellmath__39_2mx_I8575 (.Y(N5180), .A(inst_cellmath__55[13]), .B(inst_cellmath__39[13]));
NOR2X1 inst_cellmath__39_2mx_I8576 (.Y(N5260), .A(inst_cellmath__55[14]), .B(inst_cellmath__39[14]));
NAND2X2 inst_cellmath__39_2mx_I8577 (.Y(N5355), .A(inst_cellmath__55[14]), .B(inst_cellmath__39[14]));
AOI21X2 inst_cellmath__39_2mx_I8578 (.Y(N5065), .A0(N5095), .A1(N5243), .B0(N5420));
INVX2 inst_cellmath__39_2mx_I8579 (.Y(N14435), .A(N5046));
INVX2 inst_cellmath__39_2mx_I8580 (.Y(N14446), .A(N14435));
AOI21X1 inst_cellmath__39_2mx_I8581 (.Y(N14434), .A0(N5193), .A1(N14446), .B0(N5370));
NAND2X2 inst_cellmath__39_2mx_I8582 (.Y(N5106), .A(N5272), .B(N14446));
OAI21X2 inst_cellmath__39_2mx_I8583 (.Y(N5325), .A0(N5065), .A1(N5106), .B0(N14434));
INVX1 inst_cellmath__39_2mx_I8584 (.Y(N14455), .A(N5406));
INVX1 inst_cellmath__39_2mx_I8585 (.Y(N14418), .A(N14455));
AOI21X1 inst_cellmath__39_2mx_I8586 (.Y(N5265), .A0(N5133), .A1(N14418), .B0(N5317));
NAND2X1 inst_cellmath__39_2mx_I8587 (.Y(N5362), .A(N5230), .B(N14418));
AOI21XL inst_cellmath__39_2mx_I8588 (.Y(N14440), .A0(N5355), .A1(N5080), .B0(N5260));
NAND2X1 inst_cellmath__39_2mx_I8589 (.Y(N14451), .A(N5355), .B(N5180));
OAI21X2 inst_cellmath__39_2mx_I8590 (.Y(N5112), .A0(N14451), .A1(N5265), .B0(N14440));
NOR2X1 inst_cellmath__39_2mx_I8591 (.Y(N5209), .A(N14451), .B(N5362));
AOI21X2 inst_cellmath__39_2mx_I8592 (.Y(N5307), .A0(N5209), .A1(N5325), .B0(N5112));
NAND2X2 inst_cellmath__57__22__I1060 (.Y(N5332), .A(inst_cellmath__55[7]), .B(inst_cellmath__39[7]));
NAND2XL inst_cellmath__57__22__I1273 (.Y(N5161), .A(N5332), .B(N5095));
NOR2X2 inst_cellmath__57__22__I1278 (.Y(N5412), .A(N5106), .B(N5161));
NAND2X2 inst_cellmath__39_2mx_I8429 (.Y(N5398), .A(N5209), .B(N5412));
XNOR2X1 inst_cellmath__55_2mx_I1043 (.Y(inst_cellmath__55[22]), .A(N596), .B(inst_cellmath__55[0]));
NAND2X2 inst_cellmath__57__22__I1090 (.Y(N5141), .A(inst_cellmath__55[22]), .B(inst_cellmath__39[22]));
XNOR2X1 inst_cellmath__55_2mx_I1042 (.Y(inst_cellmath__55[21]), .A(N595), .B(inst_cellmath__55[0]));
NAND2X1 inst_cellmath__57__22__I1088 (.Y(N5376), .A(inst_cellmath__55[21]), .B(inst_cellmath__39[21]));
NAND2XL inst_cellmath__57__22__I1297 (.Y(N5298), .A(N5141), .B(N5376));
XNOR2X1 inst_cellmath__55_2mx_I1041 (.Y(inst_cellmath__55[20]), .A(N594), .B(inst_cellmath__55[0]));
NAND2X4 inst_cellmath__57__22__I1086 (.Y(N5201), .A(inst_cellmath__55[20]), .B(inst_cellmath__39[20]));
XNOR2X1 inst_cellmath__55_2mx_I1040 (.Y(inst_cellmath__55[19]), .A(N593), .B(inst_cellmath__55[0]));
NAND2X1 inst_cellmath__57__22__I1084 (.Y(N5426), .A(inst_cellmath__55[19]), .B(inst_cellmath__39[19]));
NAND2XL inst_cellmath__57__22__I1294 (.Y(N5354), .A(N5201), .B(N5426));
NOR2XL inst_cellmath__57__22__I1299 (.Y(N5200), .A(N5298), .B(N5354));
XNOR2X1 inst_cellmath__55_2mx_I1039 (.Y(inst_cellmath__55[18]), .A(N592), .B(inst_cellmath__55[0]));
NAND2XL inst_cellmath__57__22__I1082 (.Y(N5247), .A(inst_cellmath__55[18]), .B(inst_cellmath__39[18]));
XNOR2X1 inst_cellmath__55_2mx_I1038 (.Y(inst_cellmath__55[17]), .A(N591), .B(inst_cellmath__55[0]));
NAND2X2 inst_cellmath__57__22__I1080 (.Y(N5066), .A(inst_cellmath__55[17]), .B(inst_cellmath__39[17]));
NAND2XL inst_cellmath__57__22__I1290 (.Y(N5094), .A(N5247), .B(N5066));
XNOR2X1 inst_cellmath__55_2mx_I1037 (.Y(inst_cellmath__55[16]), .A(N590), .B(inst_cellmath__55[0]));
NAND2X2 inst_cellmath__57__22__I1078 (.Y(N5299), .A(inst_cellmath__55[16]), .B(inst_cellmath__39[16]));
XNOR2X1 inst_cellmath__55_2mx_I1036 (.Y(inst_cellmath__55[15]), .A(inst_cellmath__55[0]), .B(N589));
NOR2X1 inst_cellmath__57__22__I1075 (.Y(N5035), .A(inst_cellmath__55[15]), .B(inst_cellmath__39[15]));
NOR2X1 inst_cellmath__57__22__I1077 (.Y(N5218), .A(inst_cellmath__55[16]), .B(inst_cellmath__39[16]));
AOI21X1 inst_cellmath__57__22__I1286 (.Y(N5058), .A0(N5035), .A1(N5299), .B0(N5218));
NOR2XL inst_cellmath__57__22__I1079 (.Y(N5392), .A(inst_cellmath__55[17]), .B(inst_cellmath__39[17]));
NOR2XL inst_cellmath__57__22__I1081 (.Y(N5160), .A(inst_cellmath__55[18]), .B(inst_cellmath__39[18]));
AOI21XL inst_cellmath__57__22__I1289 (.Y(N5418), .A0(N5247), .A1(N5392), .B0(N5160));
OAI21X1 inst_cellmath__57__22__I1291 (.Y(N5316), .A0(N5094), .A1(N5058), .B0(N5418));
NOR2XL inst_cellmath__57__22__I1083 (.Y(N5340), .A(inst_cellmath__55[19]), .B(inst_cellmath__39[19]));
NOR2X1 inst_cellmath__57__22__I1085 (.Y(N5105), .A(inst_cellmath__55[20]), .B(inst_cellmath__39[20]));
AOI21XL inst_cellmath__57__22__I1293 (.Y(N5258), .A0(N5201), .A1(N5340), .B0(N5105));
NOR2XL inst_cellmath__57__22__I1087 (.Y(N5282), .A(inst_cellmath__55[21]), .B(inst_cellmath__39[21]));
NOR2XL inst_cellmath__57__22__I1089 (.Y(N5053), .A(inst_cellmath__55[22]), .B(inst_cellmath__39[22]));
AOI21XL inst_cellmath__57__22__I1296 (.Y(N5215), .A0(N5141), .A1(N5282), .B0(N5053));
OAI21XL inst_cellmath__57__22__I1298 (.Y(N5102), .A0(N5298), .A1(N5258), .B0(N5215));
AOI21X1 inst_cellmath__39_2mx_I8430 (.Y(N14148), .A0(N5200), .A1(N5316), .B0(N5102));
NAND2X2 inst_cellmath__57__22__I1076 (.Y(N5118), .A(inst_cellmath__55[15]), .B(inst_cellmath__39[15]));
NAND2X1 inst_cellmath__57__22__I1287 (.Y(N5150), .A(N5299), .B(N5118));
NOR2XL inst_cellmath__57__22__I1292 (.Y(N5405), .A(N5094), .B(N5150));
NAND2X1 inst_cellmath__39_2mx_I8431 (.Y(N14157), .A(N5200), .B(N5405));
NOR2XL inst_cellmath__39_2mx_I8594 (.Y(N5236), .A(N14173), .B(N14169));
NOR2XL inst_cellmath__39_2mx_I8595 (.Y(N5411), .A(inst_cellmath__55[24]), .B(N14181));
NAND2XL inst_cellmath__39_2mx_I8596 (.Y(N5087), .A(inst_cellmath__55[24]), .B(N14181));
NAND2XL inst_cellmath__39_2mx_I8598 (.Y(N14511), .A(N5087), .B(N5236));
NAND2XL inst_cellmath__39_2mx_I8599 (.Y(N14496), .A(N5087), .B(N5326));
INVX2 inst_cellmath__39_2mx_I8600 (.Y(N5346), .A(N5358));
OAI21X2 inst_cellmath__39_2mx_I8601 (.Y(N14508), .A0(N14157), .A1(N5307), .B0(N14148));
NOR2X2 inst_cellmath__39_2mx_I8602 (.Y(N14514), .A(N14157), .B(N5398));
AOI21X4 inst_cellmath__39_2mx_I8603 (.Y(N5352), .A0(N14514), .A1(N5346), .B0(N14508));
NOR2X4 inst_cellmath__39_2mx_I8604 (.Y(N14499), .A(N14496), .B(N5352));
NAND2BXL inst_cellmath__39_2mx_I8667 (.Y(N14504), .AN(N5411), .B(N14511));
NOR2X6 inst_cellmath__39_2mx_I8606 (.Y(N444), .A(N14504), .B(N14499));
AOI21X2 inst_cellmath__57__22__I1095 (.Y(N5361), .A0(N5075), .A1(N5311), .B0(N5400));
AOI21X1 inst_cellmath__57__22__I1096 (.Y(N5310), .A0(N5437), .A1(N5169), .B0(N5348));
NAND2XL inst_cellmath__57__22__I1097 (.Y(N5399), .A(N5437), .B(N5254));
OAI21X1 inst_cellmath__57__22__I1098 (.Y(N5208), .A0(N5399), .A1(N5361), .B0(N5310));
AOI21X2 inst_cellmath__57__22__I1099 (.Y(N5149), .A0(N5384), .A1(N5115), .B0(N5291));
NAND2X2 inst_cellmath__57__22__I1100 (.Y(N5241), .A(N5384), .B(N5211));
INVXL inst_cellmath__57__22__I1101 (.Y(N5070), .A(N5152));
AOI21X1 inst_cellmath__57__22__I1102 (.Y(N5093), .A0(N5059), .A1(N5332), .B0(N5243));
NAND2X1 inst_cellmath__57__22__I1103 (.Y(N5191), .A(N5332), .B(N5152));
OAI21X1 inst_cellmath__57__22__I1104 (.Y(N5404), .A0(N5191), .A1(N5149), .B0(N5093));
NOR2XL inst_cellmath__57__22__I1105 (.Y(N5079), .A(N5241), .B(N5191));
AOI21X2 inst_cellmath__57__22__I1106 (.Y(N5353), .A0(N5272), .A1(N5420), .B0(N5193));
NAND2X1 inst_cellmath__57__22__I1107 (.Y(N5034), .A(N5272), .B(N5095));
INVXL inst_cellmath__57__22__I1108 (.Y(N5380), .A(N5046));
AOI21X1 inst_cellmath__57__22__I1109 (.Y(N5297), .A0(N5370), .A1(N5230), .B0(N5133));
NAND2X1 inst_cellmath__57__22__I1110 (.Y(N5391), .A(N5230), .B(N5046));
OAI21X2 inst_cellmath__57__22__I1111 (.Y(N5199), .A0(N5391), .A1(N5353), .B0(N5297));
NOR2X1 inst_cellmath__57__22__I1112 (.Y(N5281), .A(N5391), .B(N5034));
AOI21X2 inst_cellmath__57__22__I8671 (.Y(N5139), .A0(N5317), .A1(N5180), .B0(N5080));
NAND2XL inst_cellmath__57__22__I1114 (.Y(N5235), .A(N5180), .B(N5406));
INVXL inst_cellmath__57__22__I1115 (.Y(N5267), .A(N5355));
AOI21X1 inst_cellmath__57__22__I1116 (.Y(N5085), .A0(N5118), .A1(N5260), .B0(N5035));
NAND2X1 inst_cellmath__57__22__I1117 (.Y(N5184), .A(N5355), .B(N5118));
OAI21X1 inst_cellmath__57__22__I1118 (.Y(N5397), .A0(N5184), .A1(N5139), .B0(N5085));
NOR2X1 inst_cellmath__57__22__I1119 (.Y(N5072), .A(N5184), .B(N5235));
AOI21X1 inst_cellmath__57__22__I1120 (.Y(N5344), .A0(N5066), .A1(N5218), .B0(N5392));
NAND2X1 inst_cellmath__57__22__I1121 (.Y(N5432), .A(N5066), .B(N5299));
INVXL inst_cellmath__57__22__I1122 (.Y(N5171), .A(N5247));
AOI21XL inst_cellmath__57__22__I1123 (.Y(N5287), .A0(N5426), .A1(N5160), .B0(N5340));
NAND2XL inst_cellmath__57__22__I1124 (.Y(N5383), .A(N5426), .B(N5247));
OAI21X1 inst_cellmath__57__22__I1125 (.Y(N5187), .A0(N5383), .A1(N5344), .B0(N5287));
NOR2XL inst_cellmath__57__22__I1126 (.Y(N5270), .A(N5383), .B(N5432));
AOI21X1 inst_cellmath__57__22__I1127 (.Y(N5129), .A0(N5376), .A1(N5105), .B0(N5282));
NAND2XL inst_cellmath__57__22__I1128 (.Y(N5228), .A(N5376), .B(N5201));
INVXL inst_cellmath__57__22__I1129 (.Y(N5060), .A(N5141));
AOI21XL inst_cellmath__57__22__I1130 (.Y(N5078), .A0(N5326), .A1(N5053), .B0(N5236));
NAND2XL inst_cellmath__57__22__I1131 (.Y(N5177), .A(N5326), .B(N5141));
OAI21XL inst_cellmath__57__22__I1132 (.Y(N5387), .A0(N5177), .A1(N5129), .B0(N5078));
NOR2XL inst_cellmath__57__22__I1133 (.Y(N5062), .A(N5177), .B(N5228));
INVXL inst_cellmath__57__22__I1134 (.Y(N5097), .A(N5208));
AOI21XL inst_cellmath__57__22__I1135 (.Y(N5336), .A0(N5079), .A1(N5208), .B0(N5404));
AOI21X1 inst_cellmath__57__22__I1136 (.Y(N5099), .A0(N5281), .A1(N5404), .B0(N5199));
NAND2X1 inst_cellmath__57__22__I1137 (.Y(N5196), .A(N5281), .B(N5079));
AOI21XL inst_cellmath__57__22__I1138 (.Y(N5276), .A0(N5072), .A1(N5199), .B0(N5397));
NAND2XL inst_cellmath__57__22__I1139 (.Y(N5373), .A(N5072), .B(N5281));
AOI21X1 inst_cellmath__57__22__I1140 (.Y(N5049), .A0(N5270), .A1(N5397), .B0(N5187));
NAND2X1 inst_cellmath__57__22__I1141 (.Y(N5136), .A(N5270), .B(N5072));
AOI21XL inst_cellmath__57__22__I1142 (.Y(N5233), .A0(N5062), .A1(N5187), .B0(N5387));
NAND2XL inst_cellmath__57__22__I1143 (.Y(N5321), .A(N5062), .B(N5270));
INVX1 inst_cellmath__57__22__I1144 (.Y(N5194), .A(N5097));
INVXL inst_cellmath__57__22__I1145 (.Y(N5274), .A(N5336));
OAI21X1 inst_cellmath__57__22__I1146 (.Y(N5303), .A0(N5136), .A1(N5099), .B0(N5049));
NOR2X1 inst_cellmath__57__22__I1147 (.Y(N5394), .A(N5136), .B(N5196));
OAI21XL inst_cellmath__57__22__I1148 (.Y(N5069), .A0(N5321), .A1(N5276), .B0(N5233));
NOR2XL inst_cellmath__57__22__I1149 (.Y(N5163), .A(N5321), .B(N5373));
INVX1 inst_cellmath__57__22__I1150 (.Y(N5371), .A(N5194));
INVX1 inst_cellmath__57__22__I1151 (.Y(N5047), .A(N5274));
OA21X1 inst_cellmath__57__22__I1152 (.Y(N5134), .A0(N5196), .A1(N5097), .B0(N5099));
OA21X1 inst_cellmath__57__22__I1153 (.Y(N5231), .A0(N5373), .A1(N5336), .B0(N5276));
AOI21X2 inst_cellmath__57__22__I1154 (.Y(N5144), .A0(N5194), .A1(N5394), .B0(N5303));
AOI21XL inst_cellmath__57__22__I1155 (.Y(N5328), .A0(N5163), .A1(N5274), .B0(N5069));
NOR2BXL inst_cellmath__57__22__I1156 (.Y(N5084), .AN(N5254), .B(N5361));
NOR2XL inst_cellmath__57__22__I1157 (.Y(N5081), .A(N5084), .B(N5169));
NOR2XL inst_cellmath__57__22__I1158 (.Y(N5306), .A(N5070), .B(N5149));
NOR2XL inst_cellmath__57__22__I1159 (.Y(N5120), .A(N5306), .B(N5059));
NOR2XL inst_cellmath__57__22__I1160 (.Y(N5110), .A(N5380), .B(N5353));
NOR2X1 inst_cellmath__57__22__I1161 (.Y(N5248), .A(N5370), .B(N5110));
AOI2BB1XL inst_cellmath__57__22__I3284 (.Y(N5377), .A0N(N5267), .A1N(N5139), .B0(N5260));
NOR2XL inst_cellmath__57__22__I1164 (.Y(N5176), .A(N5171), .B(N5344));
NOR2X1 inst_cellmath__57__22__I1165 (.Y(N5088), .A(N5176), .B(N5160));
NOR2XL inst_cellmath__57__22__I1166 (.Y(N5388), .A(N5060), .B(N5129));
NOR2X1 inst_cellmath__57__22__I1167 (.Y(N5225), .A(N5388), .B(N5053));
NAND2BXL inst_cellmath__57__22__I1168 (.Y(N5436), .AN(N5400), .B(N5075));
NAND2BXL inst_cellmath__57__22__I1169 (.Y(N5290), .AN(N5169), .B(N5254));
NAND2BXL inst_cellmath__57__22__I1170 (.Y(N5151), .AN(N5348), .B(N5437));
NAND2BXL inst_cellmath__57__22__I1171 (.Y(N5419), .AN(N5115), .B(N5211));
NAND2BXL inst_cellmath__57__22__I1172 (.Y(N5313), .AN(N5291), .B(N5384));
NAND2BXL inst_cellmath__57__22__I1173 (.Y(N5379), .AN(N5243), .B(N5332));
NAND2BXL inst_cellmath__57__22__I1174 (.Y(N5259), .AN(N5420), .B(N5095));
NAND2BXL inst_cellmath__57__22__I1175 (.Y(N5039), .AN(N5193), .B(N5272));
NAND2BXL inst_cellmath__57__22__I1176 (.Y(N5096), .AN(N5133), .B(N5230));
NAND2BXL inst_cellmath__57__22__I1177 (.Y(N5103), .AN(N5317), .B(N5406));
NAND2BXL inst_cellmath__57__22__I1178 (.Y(N5174), .AN(N5080), .B(N5180));
NAND2BXL inst_cellmath__57__22__I1179 (.Y(N5237), .AN(N5035), .B(N5118));
NAND2BXL inst_cellmath__57__22__I1180 (.Y(N5359), .AN(N5218), .B(N5299));
NAND2BXL inst_cellmath__57__22__I1181 (.Y(N5301), .AN(N5392), .B(N5066));
NAND2BXL inst_cellmath__57__22__I1182 (.Y(N5368), .AN(N5340), .B(N5426));
NAND2BXL inst_cellmath__57__22__I1183 (.Y(N5205), .AN(N5105), .B(N5201));
NAND2BXL inst_cellmath__57__22__I1184 (.Y(N5438), .AN(N5282), .B(N5376));
NAND2BXL inst_cellmath__57__22__I1185 (.Y(N5086), .AN(N5236), .B(N5326));
NAND2BXL inst_cellmath__57__22__I1186 (.Y(N5044), .AN(N5411), .B(N5087));
XNOR2X1 inst_cellmath__57__22__I1187 (.Y(N445), .A(inst_cellmath__39[0]), .B(inst_cellmath__55[0]));
XNOR2X1 inst_cellmath__57__22__I1188 (.Y(N446), .A(N5311), .B(N5436));
XNOR2X1 inst_cellmath__57__22__I1189 (.Y(N447), .A(N5361), .B(N5290));
XNOR2X1 inst_cellmath__57__22__I1190 (.Y(N448), .A(N5081), .B(N5151));
XNOR2X1 inst_cellmath__57__22__I1191 (.Y(N449), .A(N5371), .B(N5419));
XNOR2X1 inst_cellmath__57__22__I1192 (.Y(N453), .A(N5259), .B(N5047));
INVXL xnor2_A_I8760 (.Y(N14636), .A(N5103));
MXI2XL xnor2_A_I8761 (.Y(N457), .A(N5103), .B(N14636), .S0(N5134));
INVX1 xnor2_A_I3460 (.Y(N8777), .A(N5231));
MXI2X1 xnor2_A_I3461 (.Y(N461), .A(N5231), .B(N8777), .S0(N5359));
XNOR2X1 inst_cellmath__57__22__I1195 (.Y(N465), .A(N5205), .B(N5144));
XNOR2XL inst_cellmath__57__22__I1196 (.Y(N469), .A(N5044), .B(N5328));
XNOR2X1 inst_cellmath__57__22__I1197 (.Y(N5294), .A(N5211), .B(N5313));
XNOR2X1 inst_cellmath__57__22__I1198 (.Y(N5214), .A(N5115), .B(N5313));
MXI2XL inst_cellmath__57__22__I1199 (.Y(N450), .A(N5294), .B(N5214), .S0(N5371));
NOR2BXL inst_cellmath__57__22__I1200 (.Y(N5220), .AN(N5152), .B(N5059));
XNOR2X1 inst_cellmath__57__22__I1201 (.Y(N5064), .A(N5149), .B(N5220));
NAND2XL inst_cellmath__57__22__I1202 (.Y(N5037), .A(N5241), .B(N5149));
XOR2XL inst_cellmath__57__22__I1203 (.Y(N5155), .A(N5220), .B(N5037));
MXI2XL inst_cellmath__57__22__I1204 (.Y(N451), .A(N5155), .B(N5064), .S0(N5371));
XOR2XL inst_cellmath__57__22__I1205 (.Y(N5338), .A(N5379), .B(N5120));
OAI21XL inst_cellmath__57__22__I1206 (.Y(N5203), .A0(N5070), .A1(N5241), .B0(N5120));
INVXL xnor2_A_I3462 (.Y(N8783), .A(N5379));
MXI2XL xnor2_A_I3463 (.Y(N5423), .A(N5379), .B(N8783), .S0(N5203));
MXI2XL inst_cellmath__57__22__I1208 (.Y(N452), .A(N5423), .B(N5338), .S0(N5371));
XNOR2X1 inst_cellmath__57__22__I1209 (.Y(N5277), .A(N5095), .B(N5039));
XNOR2X1 inst_cellmath__57__22__I1210 (.Y(N5198), .A(N5420), .B(N5039));
MXI2XL inst_cellmath__57__22__I1211 (.Y(N454), .A(N5277), .B(N5198), .S0(N5047));
NOR2BX1 inst_cellmath__57__22__I1212 (.Y(N5349), .AN(N5046), .B(N5370));
XNOR2X1 inst_cellmath__57__22__I1213 (.Y(N5051), .A(N5353), .B(N5349));
NAND2XL inst_cellmath__57__22__I1214 (.Y(N5172), .A(N5034), .B(N5353));
XOR2XL inst_cellmath__57__22__I1215 (.Y(N5137), .A(N5349), .B(N5172));
MXI2XL inst_cellmath__57__22__I1216 (.Y(N455), .A(N5137), .B(N5051), .S0(N5047));
XOR2XL inst_cellmath__57__22__I1217 (.Y(N5323), .A(N5248), .B(N5096));
OAI21XL inst_cellmath__57__22__I1218 (.Y(N5334), .A0(N5380), .A1(N5034), .B0(N5248));
INVXL xnor2_A_I3464 (.Y(N8789), .A(N5096));
MXI2XL xnor2_A_I3465 (.Y(N5408), .A(N5096), .B(N8789), .S0(N5334));
MXI2XL inst_cellmath__57__22__I1220 (.Y(N456), .A(N5408), .B(N5323), .S0(N5047));
XNOR2X1 inst_cellmath__57__22__I1221 (.Y(N5263), .A(N5174), .B(N5406));
XNOR2X1 inst_cellmath__57__22__I1222 (.Y(N5183), .A(N5317), .B(N5174));
MXI2X1 inst_cellmath__57__22__I1223 (.Y(N458), .A(N5263), .B(N5183), .S0(N5134));
NOR2BX1 inst_cellmath__57__22__I1224 (.Y(N5067), .AN(N5355), .B(N5260));
XNOR2X1 inst_cellmath__57__22__I1225 (.Y(N5040), .A(N5139), .B(N5067));
NAND2XL inst_cellmath__57__22__I3339 (.Y(N5300), .A(N5139), .B(N5235));
XOR2XL inst_cellmath__57__22__I1227 (.Y(N5124), .A(N5067), .B(N5300));
MXI2XL inst_cellmath__57__22__I1228 (.Y(N459), .A(N5124), .B(N5040), .S0(N5134));
XOR2XL inst_cellmath__57__22__I1229 (.Y(N5305), .A(N5237), .B(N5377));
OAI21XL inst_cellmath__57__22__I1230 (.Y(N5054), .A0(N5267), .A1(N5235), .B0(N5377));
INVXL xnor2_A_I8762 (.Y(N14642), .A(N5237));
MXI2XL xnor2_A_I8763 (.Y(N5395), .A(N5237), .B(N14642), .S0(N5054));
MXI2X1 inst_cellmath__57__22__I1232 (.Y(N460), .A(N5395), .B(N5305), .S0(N5134));
XNOR2X1 inst_cellmath__57__22__I1233 (.Y(N5250), .A(N5301), .B(N5299));
XNOR2X1 inst_cellmath__57__22__I1234 (.Y(N5165), .A(N5301), .B(N5218));
MXI2XL inst_cellmath__57__22__I1235 (.Y(N462), .A(N5250), .B(N5165), .S0(N5231));
NOR2BX1 inst_cellmath__57__22__I1236 (.Y(N5210), .AN(N5247), .B(N5160));
XNOR2X1 inst_cellmath__57__22__I1237 (.Y(N5431), .A(N5210), .B(N5344));
NAND2XL inst_cellmath__57__22__I1238 (.Y(N5435), .A(N5432), .B(N5344));
XOR2XL inst_cellmath__57__22__I1239 (.Y(N5108), .A(N5210), .B(N5435));
MXI2XL inst_cellmath__57__22__I1240 (.Y(N463), .A(N5108), .B(N5431), .S0(N5231));
XOR2XL inst_cellmath__57__22__I1241 (.Y(N5286), .A(N5368), .B(N5088));
OAI21XL inst_cellmath__57__22__I1242 (.Y(N5192), .A0(N5171), .A1(N5432), .B0(N5088));
INVXL xnor2_A_I8764 (.Y(N14648), .A(N5368));
MXI2XL xnor2_A_I8765 (.Y(N5381), .A(N5368), .B(N14648), .S0(N5192));
MXI2XL inst_cellmath__57__22__I1244 (.Y(N464), .A(N5381), .B(N5286), .S0(N5231));
XNOR2X1 inst_cellmath__57__22__I1245 (.Y(N5239), .A(N5438), .B(N5201));
XNOR2X1 inst_cellmath__57__22__I1246 (.Y(N5146), .A(N5438), .B(N5105));
MXI2XL inst_cellmath__57__22__I1247 (.Y(N466), .A(N5239), .B(N5146), .S0(N5144));
NOR2BX1 inst_cellmath__57__22__I1248 (.Y(N5339), .AN(N5141), .B(N5053));
XNOR2X1 inst_cellmath__57__22__I1249 (.Y(N5415), .A(N5339), .B(N5129));
NAND2XL inst_cellmath__57__22__I1250 (.Y(N5159), .A(N5228), .B(N5129));
XOR2XL inst_cellmath__57__22__I1251 (.Y(N5090), .A(N5339), .B(N5159));
MXI2X1 inst_cellmath__57__22__I1252 (.Y(N467), .A(N5090), .B(N5415), .S0(N5144));
XOR2XL inst_cellmath__57__22__I1253 (.Y(N5269), .A(N5086), .B(N5225));
OAI21XL inst_cellmath__57__22__I1254 (.Y(N5324), .A0(N5060), .A1(N5228), .B0(N5225));
INVXL xnor2_A_I8766 (.Y(N14654), .A(N5086));
MXI2XL xnor2_A_I8767 (.Y(N5365), .A(N5086), .B(N14654), .S0(N5324));
MXI2X1 inst_cellmath__57__22__I1256 (.Y(N468), .A(N5365), .B(N5269), .S0(N5144));
INVXL inst_cellmath__57__22__I1267 (.Y(N5242), .A(N5384));
INVXL inst_cellmath__57__22__I1274 (.Y(N5132), .A(N5272));
INVXL inst_cellmath__57__22__I1281 (.Y(N5216), .A(N5180));
INVXL inst_cellmath__57__22__I1288 (.Y(N5104), .A(N5066));
INVXL inst_cellmath__57__22__I1295 (.Y(N5410), .A(N5376));
INVXL inst_cellmath__57__22__I1302 (.Y(N5167), .A(N5333));
AOI21X1 inst_cellmath__57__22__I1304 (.Y(N5126), .A0(N5412), .A1(N5119), .B0(N5325));
NAND2XL inst_cellmath__57__22__I1305 (.Y(N5222), .A(N5217), .B(N5412));
AOI21XL inst_cellmath__57__22__I1308 (.Y(N5073), .A0(N5405), .A1(N5112), .B0(N5316));
NAND2X1 inst_cellmath__57__22__I1309 (.Y(N5166), .A(N5405), .B(N5209));
INVX1 inst_cellmath__57__22__I1312 (.Y(N5253), .A(N5167));
OAI21X1 inst_cellmath__57__22__I1314 (.Y(N5330), .A0(N5166), .A1(N5126), .B0(N5073));
NOR2X1 inst_cellmath__57__22__I1315 (.Y(N5416), .A(N5166), .B(N5222));
INVX1 inst_cellmath__57__22__I1318 (.Y(N5433), .A(N5253));
INVXL inst_cellmath__57__22__I1319 (.Y(N5111), .A(N5346));
OA21X1 inst_cellmath__57__22__I1320 (.Y(N5206), .A0(N5167), .A1(N5222), .B0(N5126));
OA21X1 inst_cellmath__57__22__I1321 (.Y(N5288), .A0(N5398), .A1(N5358), .B0(N5307));
AOI21X2 inst_cellmath__57__22__I1322 (.Y(N5178), .A0(N5416), .A1(N5253), .B0(N5330));
NOR2BX1 inst_cellmath__57__22__I8676 (.Y(N5123), .AN(N5075), .B(N5076));
NOR2XL inst_cellmath__57__22__I1325 (.Y(N5147), .A(N5123), .B(N5400));
NOR2XL inst_cellmath__57__22__I1326 (.Y(N5342), .A(N5242), .B(N5273));
NOR2XL inst_cellmath__57__22__I1327 (.Y(N5189), .A(N5342), .B(N5291));
NOR2XL inst_cellmath__57__22__I1328 (.Y(N5143), .A(N5132), .B(N5065));
NOR2XL inst_cellmath__57__22__I1329 (.Y(N5314), .A(N5143), .B(N5193));
NOR2XL inst_cellmath__57__22__I1330 (.Y(N5364), .A(N5216), .B(N5265));
NOR2XL inst_cellmath__57__22__I1331 (.Y(N5032), .A(N5364), .B(N5080));
NOR2XL inst_cellmath__57__22__I1332 (.Y(N5170), .A(N5104), .B(N5058));
NOR2XL inst_cellmath__57__22__I1333 (.Y(N5157), .A(N5170), .B(N5392));
NOR2XL inst_cellmath__57__22__I1334 (.Y(N5385), .A(N5410), .B(N5258));
NOR2XL inst_cellmath__57__22__I1335 (.Y(N5279), .A(N5385), .B(N5282));
NAND2BXL inst_cellmath__57__22__I1336 (.Y(N5319), .AN(N5350), .B(N5311));
XOR2XL inst_cellmath__57__22__I1337 (.Y(N419), .A(inst_cellmath__55[24]), .B(N5319));
XNOR2X1 inst_cellmath__57__22__I1338 (.Y(N420), .A(N5076), .B(N5436));
XNOR2X1 inst_cellmath__57__22__I1341 (.Y(N426), .A(N5111), .B(N5379));
XNOR2X1 inst_cellmath__57__22__I1342 (.Y(N430), .A(N5096), .B(N5206));
XNOR2X1 inst_cellmath__57__22__I1343 (.Y(N434), .A(N5237), .B(N5288));
XNOR2XL inst_cellmath__57__22__I1344 (.Y(N438), .A(N5368), .B(N5178));
XNOR2X1 inst_cellmath__57__22__I1345 (.Y(N442), .A(N5352), .B(N5086));
XNOR2X1 inst_cellmath__57__22__I1346 (.Y(N5041), .A(N5437), .B(N5419));
XNOR2X1 inst_cellmath__57__22__I1347 (.Y(N5360), .A(N5348), .B(N5419));
MXI2XL inst_cellmath__57__22__I1348 (.Y(N423), .A(N5041), .B(N5360), .S0(N5433));
XOR2XL inst_cellmath__57__22__I1349 (.Y(N5223), .A(N5273), .B(N5313));
NAND2XL inst_cellmath__57__22__I1350 (.Y(N5130), .A(N5369), .B(N5273));
XNOR2X1 inst_cellmath__57__22__I1351 (.Y(N5308), .A(N5313), .B(N5130));
MXI2XL inst_cellmath__57__22__I1352 (.Y(N424), .A(N5308), .B(N5223), .S0(N5433));
XNOR2X1 inst_cellmath__57__22__I1353 (.Y(N5074), .A(N5220), .B(N5189));
OAI21XL inst_cellmath__57__22__I1354 (.Y(N5293), .A0(N5242), .A1(N5369), .B0(N5189));
XOR2XL inst_cellmath__57__22__I1355 (.Y(N5168), .A(N5220), .B(N5293));
MXI2XL inst_cellmath__57__22__I1356 (.Y(N425), .A(N5168), .B(N5074), .S0(N5433));
XNOR2X1 inst_cellmath__57__22__I1357 (.Y(N5434), .A(N5332), .B(N5259));
XNOR2X1 inst_cellmath__57__22__I1358 (.Y(N5347), .A(N5243), .B(N5259));
MXI2XL inst_cellmath__57__22__I1359 (.Y(N427), .A(N5434), .B(N5347), .S0(N5111));
XOR2XL inst_cellmath__57__22__I1360 (.Y(N5207), .A(N5065), .B(N5039));
NAND2XL inst_cellmath__57__22__I1361 (.Y(N5262), .A(N5065), .B(N5161));
XNOR2X1 inst_cellmath__57__22__I1362 (.Y(N5289), .A(N5039), .B(N5262));
MXI2XL inst_cellmath__57__22__I1363 (.Y(N428), .A(N5289), .B(N5207), .S0(N5111));
XNOR2X1 inst_cellmath__57__22__I1364 (.Y(N5057), .A(N5349), .B(N5314));
OAI21XL inst_cellmath__57__22__I1365 (.Y(N5430), .A0(N5132), .A1(N5161), .B0(N5314));
XOR2XL inst_cellmath__57__22__I1366 (.Y(N5148), .A(N5349), .B(N5430));
MXI2XL inst_cellmath__57__22__I1367 (.Y(N429), .A(N5148), .B(N5057), .S0(N5111));
XNOR2X1 inst_cellmath__57__22__I1368 (.Y(N5417), .A(N5103), .B(N5230));
XNOR2X1 inst_cellmath__57__22__I1369 (.Y(N5331), .A(N5133), .B(N5103));
MXI2XL inst_cellmath__57__22__I1370 (.Y(N431), .A(N5417), .B(N5331), .S0(N5206));
XOR2XL inst_cellmath__57__22__I1371 (.Y(N5190), .A(N5265), .B(N5174));
NAND2XL inst_cellmath__57__22__I1372 (.Y(N5402), .A(N5362), .B(N5265));
XNOR2X1 inst_cellmath__57__22__I1373 (.Y(N5271), .A(N5174), .B(N5402));
MXI2XL inst_cellmath__57__22__I1374 (.Y(N432), .A(N5271), .B(N5190), .S0(N5206));
XNOR2X1 inst_cellmath__57__22__I1375 (.Y(N5045), .A(N5067), .B(N5032));
OAI21XL inst_cellmath__57__22__I1376 (.Y(N5154), .A0(N5216), .A1(N5362), .B0(N5032));
XOR2XL inst_cellmath__57__22__I1377 (.Y(N5131), .A(N5067), .B(N5154));
MXI2XL inst_cellmath__57__22__I1378 (.Y(N433), .A(N5131), .B(N5045), .S0(N5206));
XNOR2X1 inst_cellmath__57__22__I1379 (.Y(N5403), .A(N5359), .B(N5118));
XNOR2X1 inst_cellmath__57__22__I1380 (.Y(N5315), .A(N5035), .B(N5359));
MXI2XL inst_cellmath__57__22__I1381 (.Y(N435), .A(N5403), .B(N5315), .S0(N5288));
XOR2XL inst_cellmath__57__22__I1382 (.Y(N5179), .A(N5301), .B(N5058));
NAND2XL inst_cellmath__57__22__I1383 (.Y(N5122), .A(N5150), .B(N5058));
XNOR2X1 inst_cellmath__57__22__I1384 (.Y(N5257), .A(N5301), .B(N5122));
MXI2XL inst_cellmath__57__22__I1385 (.Y(N436), .A(N5257), .B(N5179), .S0(N5288));
XNOR2X1 inst_cellmath__57__22__I1386 (.Y(N5033), .A(N5210), .B(N5157));
OAI21XL inst_cellmath__57__22__I1387 (.Y(N5283), .A0(N5104), .A1(N5150), .B0(N5157));
XOR2XL inst_cellmath__57__22__I1388 (.Y(N5117), .A(N5210), .B(N5283));
MXI2XL inst_cellmath__57__22__I1389 (.Y(N437), .A(N5117), .B(N5033), .S0(N5288));
XNOR2X1 inst_cellmath__57__22__I1390 (.Y(N5390), .A(N5205), .B(N5426));
XNOR2X1 inst_cellmath__57__22__I1391 (.Y(N5296), .A(N5205), .B(N5340));
MXI2XL inst_cellmath__57__22__I1392 (.Y(N439), .A(N5390), .B(N5296), .S0(N5178));
XOR2XL inst_cellmath__57__22__I1393 (.Y(N5158), .A(N5438), .B(N5258));
NAND2XL inst_cellmath__57__22__I1394 (.Y(N5255), .A(N5354), .B(N5258));
XNOR2X1 inst_cellmath__57__22__I1395 (.Y(N5246), .A(N5438), .B(N5255));
MXI2XL inst_cellmath__57__22__I1396 (.Y(N440), .A(N5246), .B(N5158), .S0(N5178));
XNOR2X1 inst_cellmath__57__22__I1397 (.Y(N5425), .A(N5339), .B(N5279));
OAI21XL inst_cellmath__57__22__I1398 (.Y(N5421), .A0(N5410), .A1(N5354), .B0(N5279));
XOR2XL inst_cellmath__57__22__I1399 (.Y(N5101), .A(N5339), .B(N5421));
MXI2XL inst_cellmath__57__22__I1400 (.Y(N441), .A(N5101), .B(N5425), .S0(N5178));
XNOR2X1 inst_cellmath__57__22__I1401 (.Y(N5375), .A(N5044), .B(N5326));
XNOR2X1 inst_cellmath__57__22__I1402 (.Y(N5280), .A(N5044), .B(N5236));
MXI2XL inst_cellmath__57__22__I1403 (.Y(N443), .A(N5375), .B(N5280), .S0(N5352));
NAND2XL cynw_cm_float_add2_I1406 (.Y(N418), .A(a_sign), .B(inst_cellmath__28));
NAND2XL cynw_cm_float_add2_I1408 (.Y(N417), .A(b_sign), .B(inst_cellmath__31));
MX2XL inst_cellmath__52_0_I1409 (.Y(N5814), .A(N417), .B(N418), .S0(N517));
MXI2XL inst_cellmath__52_0_I1410 (.Y(N5817), .A(a_sign), .B(b_sign), .S0(N517));
CLKINVX12 inst_delta_0_I8538 (.Y(inst_cellmath__56[25]), .A(N444));
MX2XL inst_cellmath__52_0_I1411 (.Y(inst_cellmath__52), .A(N5817), .B(N5814), .S0(inst_cellmath__56[25]));
NOR2XL cynw_cm_float_add2_I1412 (.Y(inst_cellmath__51[25]), .A(inst_cellmath__55[0]), .B(inst_cellmath__56[25]));
MXI2XL cynw_cm_float_add2_I1414 (.Y(N5914), .A(inst_cellmath__55[0]), .B(inst_cellmath__55[24]), .S0(N445));
MXI2XL cynw_cm_float_add2_I1415 (.Y(N5829), .A(inst_cellmath__55[0]), .B(inst_cellmath__55[24]), .S0(N446));
MXI2XL cynw_cm_float_add2_I1418 (.Y(N5901), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N449));
MXI2XL cynw_cm_float_add2_I1419 (.Y(N5927), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N450));
MXI2XL cynw_cm_float_add2_I1420 (.Y(N5840), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N451));
MXI2XL cynw_cm_float_add2_I1421 (.Y(N5863), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N452));
MXI2XL cynw_cm_float_add2_I1422 (.Y(N5887), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N453));
MXI2XL cynw_cm_float_add2_I1423 (.Y(N5911), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N454));
MXI2XL cynw_cm_float_add2_I1424 (.Y(N5936), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N455));
MXI2XL cynw_cm_float_add2_I1425 (.Y(N5849), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N456));
MXI2XL cynw_cm_float_add2_I1426 (.Y(N5873), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N457));
MXI2XL cynw_cm_float_add2_I1427 (.Y(N5895), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N458));
MXI2XL cynw_cm_float_add2_I1428 (.Y(N5922), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N459));
MXI2XL cynw_cm_float_add2_I1429 (.Y(N5836), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N460));
MXI2X1 cynw_cm_float_add2_I1430 (.Y(N5858), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N461));
MXI2XL cynw_cm_float_add2_I1431 (.Y(N5883), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N462));
MXI2XL cynw_cm_float_add2_I1432 (.Y(N5906), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N463));
MXI2XL cynw_cm_float_add2_I1433 (.Y(N5932), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N464));
MXI2X1 cynw_cm_float_add2_I8681 (.Y(N5845), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N465));
MXI2XL cynw_cm_float_add2_I1435 (.Y(N5869), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N466));
MXI2XL cynw_cm_float_add2_I1436 (.Y(N5892), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N467));
MXI2XL cynw_cm_float_add2_I1437 (.Y(N5918), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N468));
MXI2X1 cynw_cm_float_add2_I1438 (.Y(N5832), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N469));
CLKINVX12 inst_delta_0_I8540 (.Y(N5850), .A(inst_cellmath__56[25]));
AOI22XL cynw_cm_float_add2_I1447 (.Y(N474), .A0(N423), .A1(N5850), .B0(N5901), .B1(inst_cellmath__56[25]));
AOI22XL cynw_cm_float_add2_I1448 (.Y(N475), .A0(N424), .A1(N5850), .B0(N5927), .B1(inst_cellmath__56[25]));
AOI22X1 cynw_cm_float_add2_I1450 (.Y(N476), .A0(N425), .A1(N5850), .B0(N5840), .B1(inst_cellmath__56[25]));
AOI22X1 cynw_cm_float_add2_I1451 (.Y(N477), .A0(N5850), .A1(N426), .B0(inst_cellmath__56[25]), .B1(N5863));
AOI22X1 cynw_cm_float_add2_I1452 (.Y(N478), .A0(N427), .A1(N5850), .B0(N5887), .B1(inst_cellmath__56[25]));
AOI22X1 cynw_cm_float_add2_I1453 (.Y(N479), .A0(N428), .A1(N5850), .B0(N5911), .B1(inst_cellmath__56[25]));
AOI22X1 cynw_cm_float_add2_I1456 (.Y(N482), .A0(N431), .A1(N5850), .B0(N5873), .B1(inst_cellmath__56[25]));
AOI22X1 cynw_cm_float_add2_I1457 (.Y(N483), .A0(N432), .A1(N5850), .B0(N5895), .B1(inst_cellmath__56[25]));
AOI22XL cynw_cm_float_add2_I1458 (.Y(N484), .A0(N433), .A1(N5850), .B0(N5922), .B1(inst_cellmath__56[25]));
AOI22X1 cynw_cm_float_add2_I1462 (.Y(N487), .A0(N436), .A1(N5850), .B0(N5883), .B1(inst_cellmath__56[25]));
AOI22XL cynw_cm_float_add2_I1464 (.Y(N489), .A0(N438), .A1(N5850), .B0(inst_cellmath__56[25]), .B1(N5932));
AOI22X1 cynw_cm_float_add2_I1465 (.Y(N490), .A0(N439), .A1(N5850), .B0(inst_cellmath__56[25]), .B1(N5845));
AOI22XL cynw_cm_float_add2_I1466 (.Y(N491), .A0(N440), .A1(N5850), .B0(inst_cellmath__56[25]), .B1(N5869));
AOI22XL cynw_cm_float_add2_I1469 (.Y(N494), .A0(N443), .A1(N5850), .B0(inst_cellmath__56[25]), .B1(N5832));
INVX1 cynw_cm_float_add2_I42 (.Y(inst_cellmath__51[4]), .A(N474));
INVX1 cynw_cm_float_add2_I43 (.Y(inst_cellmath__51[5]), .A(N475));
INVX2 cynw_cm_float_add2_I44 (.Y(inst_cellmath__51[6]), .A(N476));
INVX2 cynw_cm_float_add2_I45 (.Y(inst_cellmath__51[7]), .A(N477));
INVX1 cynw_cm_float_add2_I46 (.Y(inst_cellmath__51[8]), .A(N478));
INVX1 cynw_cm_float_add2_I47 (.Y(inst_cellmath__51[9]), .A(N479));
AO22X1 cynw_cm_float_add2_I3347 (.Y(inst_cellmath__51[10]), .A0(inst_cellmath__56[25]), .A1(N5936), .B0(N5850), .B1(N429));
AO22X1 cynw_cm_float_add2_I3348 (.Y(inst_cellmath__51[11]), .A0(inst_cellmath__56[25]), .A1(N5849), .B0(N5850), .B1(N430));
INVX1 cynw_cm_float_add2_I50 (.Y(inst_cellmath__51[12]), .A(N482));
INVX1 cynw_cm_float_add2_I51 (.Y(inst_cellmath__51[13]), .A(N483));
INVX1 cynw_cm_float_add2_I52 (.Y(inst_cellmath__51[14]), .A(N484));
AO22X1 cynw_cm_float_add2_I3279 (.Y(inst_cellmath__51[15]), .A0(N5836), .A1(inst_cellmath__56[25]), .B0(N5850), .B1(N434));
AO22X1 cynw_cm_float_add2_I3350 (.Y(inst_cellmath__51[16]), .A0(inst_cellmath__56[25]), .A1(N5858), .B0(N435), .B1(N5850));
INVX1 cynw_cm_float_add2_I55 (.Y(inst_cellmath__51[17]), .A(N487));
AO22X1 cynw_cm_float_add2_I3352 (.Y(inst_cellmath__51[18]), .A0(inst_cellmath__56[25]), .A1(N5906), .B0(N437), .B1(N5850));
INVX1 cynw_cm_float_add2_I57 (.Y(inst_cellmath__51[19]), .A(N489));
INVX1 cynw_cm_float_add2_I58 (.Y(inst_cellmath__51[20]), .A(N490));
INVX1 cynw_cm_float_add2_I59 (.Y(inst_cellmath__51[21]), .A(N491));
AO22X1 cynw_cm_float_add2_I3355 (.Y(inst_cellmath__51[22]), .A0(N5892), .A1(inst_cellmath__56[25]), .B0(N441), .B1(N5850));
AO22X1 cynw_cm_float_add2_I3356 (.Y(inst_cellmath__51[23]), .A0(inst_cellmath__56[25]), .A1(N5918), .B0(N442), .B1(N5850));
INVX1 cynw_cm_float_add2_I62 (.Y(inst_cellmath__51[24]), .A(N494));
AOI22XL inst_delta_0_I8460 (.Y(N14264), .A0(N419), .A1(N5850), .B0(N5914), .B1(inst_cellmath__56[25]));
INVXL inst_delta_0_I8461 (.Y(inst_cellmath__51[0]), .A(N14264));
AOI22XL inst_delta_0_I8462 (.Y(N14271), .A0(N420), .A1(N5850), .B0(N5829), .B1(inst_cellmath__56[25]));
INVXL inst_delta_0_I8463 (.Y(inst_cellmath__51[1]), .A(N14271));
NOR2BX1 inst_delta_0_I1470 (.Y(N6086), .AN(inst_cellmath__51[0]), .B(inst_cellmath__51[1]));
XNOR2X1 inst_delta_0_I8539 (.Y(N14358), .A(N5147), .B(N5290));
MXI2XL inst_delta_0_I8541 (.Y(N14368), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N447));
INVXL inst_delta_0_I8542 (.Y(N14377), .A(N5850));
AOI22XL inst_delta_0_I8543 (.Y(N14360), .A0(N14358), .A1(N5850), .B0(N14368), .B1(N14377));
INVXL inst_delta_0_I8544 (.Y(inst_cellmath__51[2]), .A(N14360));
XNOR2X1 inst_delta_0_I8545 (.Y(N14362), .A(N5433), .B(N5151));
MXI2XL inst_delta_0_I8546 (.Y(N14373), .A(inst_cellmath__55[24]), .B(inst_cellmath__55[0]), .S0(N448));
AOI22XL inst_delta_0_I8547 (.Y(N14365), .A0(N14362), .A1(N5850), .B0(N14373), .B1(N14377));
INVX1 inst_delta_0_I8548 (.Y(inst_cellmath__51[3]), .A(N14365));
NOR2BX1 inst_delta_0_I1472 (.Y(N6011), .AN(inst_cellmath__51[2]), .B(inst_cellmath__51[3]));
INVXL inst_delta_0_I1473 (.Y(N6030), .A(inst_cellmath__51[5]));
OAI21XL inst_delta_0_I1474 (.Y(N6052), .A0(inst_cellmath__51[4]), .A1(N6011), .B0(N6030));
NOR2BX1 inst_delta_0_I1477 (.Y(N6040), .AN(inst_cellmath__51[6]), .B(inst_cellmath__51[7]));
INVXL inst_delta_0_I1478 (.Y(N6060), .A(inst_cellmath__51[9]));
OAI21XL inst_delta_0_I1479 (.Y(N6083), .A0(inst_cellmath__51[8]), .A1(N6040), .B0(N6060));
NOR2BXL inst_delta_0_I1482 (.Y(N6070), .AN(inst_cellmath__51[10]), .B(inst_cellmath__51[11]));
INVXL inst_delta_0_I1483 (.Y(N6090), .A(inst_cellmath__51[13]));
OAI21XL inst_delta_0_I1484 (.Y(N6017), .A0(inst_cellmath__51[12]), .A1(N6070), .B0(N6090));
NOR2X2 inst_delta_0_I1485 (.Y(N6037), .A(inst_cellmath__51[11]), .B(inst_cellmath__51[10]));
NOR2X2 inst_delta_0_I1486 (.Y(N6057), .A(inst_cellmath__51[13]), .B(inst_cellmath__51[12]));
NOR2BXL inst_delta_0_I1487 (.Y(N6003), .AN(inst_cellmath__51[14]), .B(inst_cellmath__51[15]));
INVXL inst_delta_0_I1488 (.Y(N6024), .A(inst_cellmath__51[17]));
OAI21XL inst_delta_0_I1489 (.Y(N6045), .A0(inst_cellmath__51[16]), .A1(N6003), .B0(N6024));
NOR2X2 inst_delta_0_I1490 (.Y(N6067), .A(inst_cellmath__51[15]), .B(inst_cellmath__51[14]));
NOR2X4 inst_delta_0_I1491 (.Y(N6088), .A(inst_cellmath__51[17]), .B(inst_cellmath__51[16]));
NOR2BX1 inst_delta_0_I1492 (.Y(N6032), .AN(inst_cellmath__51[18]), .B(inst_cellmath__51[19]));
INVXL inst_delta_0_I1493 (.Y(N6054), .A(inst_cellmath__51[21]));
OAI21XL inst_delta_0_I1494 (.Y(N6076), .A0(inst_cellmath__51[20]), .A1(N6032), .B0(N6054));
NOR2X2 inst_delta_0_I1495 (.Y(N6000), .A(inst_cellmath__51[19]), .B(inst_cellmath__51[18]));
NOR2X2 inst_delta_0_I1496 (.Y(N6021), .A(inst_cellmath__51[21]), .B(inst_cellmath__51[20]));
NOR2BXL inst_delta_0_I1497 (.Y(N6062), .AN(inst_cellmath__51[22]), .B(inst_cellmath__51[23]));
INVXL inst_delta_0_I1498 (.Y(N6085), .A(inst_cellmath__51[25]));
OAI21XL inst_delta_0_I1499 (.Y(N6009), .A0(inst_cellmath__51[24]), .A1(N6062), .B0(N6085));
NOR2X4 inst_delta_0_I1500 (.Y(N6028), .A(inst_cellmath__51[23]), .B(inst_cellmath__51[22]));
NOR2X2 inst_delta_0_I1501 (.Y(N6050), .A(inst_cellmath__51[25]), .B(inst_cellmath__51[24]));
MXI2XL inst_delta_0_I8549 (.Y(N14357), .A(N14362), .B(N14373), .S0(inst_cellmath__56[25]));
MXI2XL inst_delta_0_I8550 (.Y(N14367), .A(N14358), .B(N14368), .S0(inst_cellmath__56[25]));
AND2X1 inst_delta_0_I8686 (.Y(N6074), .A(N14357), .B(N14367));
NOR2X4 inst_delta_0_I8466 (.Y(N5998), .A(inst_cellmath__51[5]), .B(inst_cellmath__51[4]));
NAND2BXL inst_delta_0_I1502 (.Y(N6046), .AN(N6074), .B(N5998));
NAND2BXL inst_delta_0_I1505 (.Y(N6077), .AN(N6037), .B(N6057));
INVXL inst_delta_0_I1506 (.Y(N6001), .A(N6088));
AOI21XL inst_delta_0_I1507 (.Y(N6022), .A0(N6067), .A1(N6077), .B0(N6001));
NAND2X2 inst_delta_0_I1508 (.Y(N6042), .A(N6057), .B(N6037));
NAND2X4 inst_delta_0_I1509 (.Y(N6063), .A(N6067), .B(N6088));
NAND2BXL inst_delta_0_I1510 (.Y(N6010), .AN(N6000), .B(N6021));
INVXL inst_delta_0_I1511 (.Y(N6029), .A(N6050));
AOI21X1 inst_delta_0_I1512 (.Y(N6051), .A0(N6028), .A1(N6010), .B0(N6029));
NAND2X2 inst_delta_0_I1513 (.Y(N6073), .A(N6021), .B(N6000));
NAND2X4 inst_delta_0_I1514 (.Y(N5997), .A(N6050), .B(N6028));
NOR2X4 inst_delta_0_I8467 (.Y(N14270), .A(inst_cellmath__51[6]), .B(inst_cellmath__51[7]));
NOR2X4 inst_delta_0_I8468 (.Y(N6026), .A(inst_cellmath__51[9]), .B(inst_cellmath__51[8]));
NAND2X6 inst_delta_0_I8470 (.Y(N6033), .A(N14270), .B(N6026));
NAND2X6 inst_delta_0_I8469 (.Y(N6014), .A(N6074), .B(N5998));
NAND2BXL inst_delta_0_I1515 (.Y(N6082), .AN(N6033), .B(N6014));
NOR2BXL inst_delta_0_I1517 (.Y(N6016), .AN(N6042), .B(N6063));
INVXL inst_delta_0_I1518 (.Y(N6036), .A(N5997));
OAI21XL inst_delta_0_I1519 (.Y(N6055), .A0(N6073), .A1(N6016), .B0(N6036));
NOR2X4 inst_delta_0_I1520 (.Y(N6080), .A(N6042), .B(N6063));
NOR2X4 inst_delta_0_I1521 (.Y(N6034), .A(N5997), .B(N6073));
NOR2XL inst_delta_0_I8464 (.Y(N6064), .A(inst_cellmath__51[1]), .B(inst_cellmath__51[0]));
NOR2X6 inst_delta_0_I8471 (.Y(N6069), .A(N6033), .B(N6014));
NAND2X1 inst_delta_0_I8472 (.Y(N14283), .A(N14271), .B(N14264));
NAND2X4 inst_delta_0_I8473 (.Y(N6044), .A(N14283), .B(N6069));
INVXL buf1_A_I8768 (.Y(N14662), .A(N14270));
INVXL buf1_A_I8769 (.Y(N6007), .A(N14662));
INVX2 inst_delta_0_I1523 (.Y(N6066), .A(N6034));
AOI21X4 inst_delta_0_I1524 (.Y(inst_delta[3]), .A0(N6080), .A1(N6044), .B0(N6066));
NAND2XL inst_delta_0_I1525 (.Y(N6013), .A(N6069), .B(N6064));
NAND2X2 inst_cellmath__63_0_I8608 (.Y(N6079), .A(N6080), .B(N6034));
NOR2BX2 inst_delta_0_I1527 (.Y(inst_delta[4]), .AN(N6013), .B(N6079));
NOR2XL inst_delta_0_I1528 (.Y(inst_delta[5]), .A(N6013), .B(N6079));
OAI21XL inst_delta_0_I1533 (.Y(N6072), .A0(N6033), .A1(N6052), .B0(N6083));
OAI21XL inst_delta_0_I1534 (.Y(N6019), .A0(N6017), .A1(N6063), .B0(N6045));
OAI21XL inst_delta_0_I1535 (.Y(N6059), .A0(N5997), .A1(N6076), .B0(N6009));
AOI21XL inst_delta_0_I1536 (.Y(N6005), .A0(N6069), .A1(N6086), .B0(N6072));
AOI21XL inst_delta_0_I1537 (.Y(N6047), .A0(N6034), .A1(N6019), .B0(N6059));
OA21X1 cynw_cm_float_add2_I8688 (.Y(N2396), .A0(N6082), .A1(N6079), .B0(N6055));
OR2XL cynw_cm_float_add2_I1540 (.Y(N496), .A(inst_cellmath__52), .B(inst_delta[5]));
OAI2BB1X1 cynw_cm_float_add2_I3359 (.Y(N6171), .A0N(a_sign), .A1N(b_sign), .B0(N496));
AOI31X1 inst_cellmath__63_0_I8477 (.Y(N14317), .A0(inst_cellmath__21), .A1(inst_cellmath__24), .A2(inst_cellmath__55[0]), .B0(N4450));
INVXL inst_cellmath__63_0_I8478 (.Y(inst_cellmath__62), .A(N14317));
NOR2BX1 cynw_cm_float_add2_I3360 (.Y(x[31]), .AN(N6171), .B(inst_cellmath__62));
INVXL cynw_cm_float_add2_I1546 (.Y(N6223), .A(b_exp[0]));
INVXL cynw_cm_float_add2_I1547 (.Y(N6189), .A(b_exp[1]));
INVXL cynw_cm_float_add2_I1548 (.Y(N6198), .A(b_exp[2]));
INVXL cynw_cm_float_add2_I1549 (.Y(N6207), .A(b_exp[3]));
INVXL cynw_cm_float_add2_I1550 (.Y(N6217), .A(b_exp[4]));
INVXL cynw_cm_float_add2_I1551 (.Y(N6227), .A(b_exp[5]));
INVXL cynw_cm_float_add2_I1552 (.Y(N6192), .A(b_exp[6]));
INVXL cynw_cm_float_add2_I1553 (.Y(N6201), .A(b_exp[7]));
INVXL cynw_cm_float_add2_I1554 (.Y(N6211), .A(N3782));
INVXL cynw_cm_float_add2_I1564 (.Y(N6186), .A(N4170));
AOI22XL cynw_cm_float_add2_I1566 (.Y(inst_cellmath__40[0]), .A0(N6186), .A1(N6211), .B0(N6223), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1567 (.Y(inst_cellmath__40[1]), .A0(N501), .A1(N6186), .B0(N6189), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1568 (.Y(inst_cellmath__40[2]), .A0(N502), .A1(N6186), .B0(N6198), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1569 (.Y(inst_cellmath__40[3]), .A0(N503), .A1(N6186), .B0(N6207), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1570 (.Y(inst_cellmath__40[4]), .A0(N6186), .A1(N504), .B0(N6217), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1571 (.Y(inst_cellmath__40[5]), .A0(N505), .A1(N6186), .B0(N6227), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1572 (.Y(inst_cellmath__40[6]), .A0(N506), .A1(N6186), .B0(N6192), .B1(N4170));
AOI22XL cynw_cm_float_add2_I1573 (.Y(inst_cellmath__40[7]), .A0(N6186), .A1(N507), .B0(N6201), .B1(N4170));
INVXL inst_cellmath__73_0_I1574 (.Y(N6264), .A(inst_cellmath__40[1]));
INVXL inst_cellmath__73_0_I1575 (.Y(N6279), .A(inst_cellmath__40[2]));
INVXL inst_cellmath__73_0_I1576 (.Y(N6259), .A(inst_cellmath__40[3]));
INVXL inst_cellmath__73_0_I1577 (.Y(N6274), .A(inst_cellmath__40[4]));
OAI21X1 inst_cellmath__63_0_I8615 (.Y(inst_delta[0]), .A0(N6005), .A1(N6079), .B0(N6047));
NAND2BXL inst_cellmath__73_0_I1578 (.Y(N6260), .AN(inst_cellmath__40[0]), .B(inst_delta[0]));
OAI2BB1XL inst_cellmath__63_0_I8609 (.Y(N14573), .A0N(N6007), .A1N(N6046), .B0(N6026));
AOI21X1 inst_cellmath__63_0_I8610 (.Y(N14535), .A0(N6034), .A1(N6022), .B0(N6051));
OAI21X2 inst_cellmath__63_0_I8614 (.Y(inst_delta[1]), .A0(N14573), .A1(N6079), .B0(N14535));
NAND2XL inst_cellmath__73_0_I1579 (.Y(N6284), .A(N6264), .B(inst_delta[1]));
NOR2X1 inst_cellmath__73_0_I1580 (.Y(N6275), .A(N6264), .B(inst_delta[1]));
INVX1 inst_cellmath__63_0_I8476 (.Y(N2397), .A(N2396));
NAND2X1 inst_cellmath__73_0_I1581 (.Y(N6270), .A(N6279), .B(N2397));
NAND2XL inst_cellmath__73_0_I1583 (.Y(N6257), .A(N6259), .B(inst_delta[3]));
NOR2XL inst_cellmath__73_0_I1584 (.Y(N6288), .A(N6259), .B(inst_delta[3]));
NOR2XL inst_cellmath__73_0_I1586 (.Y(N6273), .A(N6274), .B(inst_delta[4]));
NOR2XL inst_cellmath__73_0_I1587 (.Y(N6277), .A(inst_cellmath__40[7]), .B(inst_cellmath__40[6]));
NAND4BX1 inst_cellmath__73_0_I8690 (.Y(N6266), .AN(inst_cellmath__40[5]), .B(N6274), .C(N6277), .D(inst_delta[4]));
NOR2XL inst_cellmath__73_0_I1589 (.Y(N6265), .A(inst_cellmath__40[5]), .B(N6273));
OAI21X1 inst_cellmath__73_0_I1590 (.Y(N6272), .A0(N6288), .A1(N6270), .B0(N6257));
AOI2BB1X1 inst_cellmath__73_0_I3270 (.Y(N6280), .A0N(N6279), .A1N(N2397), .B0(N6288));
OAI21X1 inst_cellmath__73_0_I1592 (.Y(N6290), .A0(N6275), .A1(N6260), .B0(N6284));
NAND2X1 inst_cellmath__73_0_I1594 (.Y(N6286), .A(N6277), .B(N6265));
AOI21X2 inst_cellmath__73_0_I1595 (.Y(N6256), .A0(N6280), .A1(N6290), .B0(N6272));
OAI21X2 inst_cellmath__73_0_I1596 (.Y(inst_cellmath__73), .A0(N6286), .A1(N6256), .B0(N6266));
AND4XL inst_cellmath__75__32__I1597 (.Y(N6325), .A(inst_cellmath__40[7]), .B(inst_cellmath__40[2]), .C(inst_cellmath__40[4]), .D(inst_cellmath__40[3]));
NAND2XL inst_cellmath__75__32__I1598 (.Y(N6315), .A(N6325), .B(inst_cellmath__40[6]));
NAND3XL hyperpropagate_4_1_A_I3472 (.Y(N8813), .A(inst_cellmath__40[5]), .B(inst_cellmath__40[1]), .C(inst_cellmath__51[25]));
NOR2XL hyperpropagate_4_1_A_I3473 (.Y(N499), .A(N6315), .B(N8813));
OR4X1 cynw_cm_float_add2_I3363 (.Y(inst_cellmath__77), .A(inst_cellmath__21), .B(inst_cellmath__24), .C(inst_cellmath__62), .D(N499));
NOR2XL cynw_cm_float_add2_I1604 (.Y(N498), .A(inst_cellmath__31), .B(inst_cellmath__28));
OR3X1 inst_cellmath__72_0_I3364 (.Y(N6354), .A(N498), .B(inst_cellmath__77), .C(inst_delta[5]));
NOR2X2 inst_cellmath__63_0_I8490 (.Y(N14301), .A(N6354), .B(inst_cellmath__73));
INVX2 inst_cellmath__63_0_I8491 (.Y(N6348), .A(N14301));
INVX1 inst_cellmath__72_0_I3310 (.Y(N8759), .A(N6348));
INVX2 inst_cellmath__72_0_I3311 (.Y(N8760), .A(N8759));
INVXL inst_cellmath__66_0_I1611 (.Y(N6399), .A(inst_delta[0]));
INVXL inst_cellmath__66_0_I1613 (.Y(N6423), .A(inst_delta[3]));
INVX1 inst_cellmath__66_0_I1614 (.Y(N6381), .A(inst_delta[4]));
ADDHX1 inst_cellmath__66_0_I1615 (.CO(N6417), .S(N6398), .A(inst_cellmath__40[2]), .B(inst_cellmath__40[1]));
ADDHX1 inst_cellmath__66_0_I1616 (.CO(N6375), .S(N6437), .A(inst_cellmath__40[3]), .B(N6417));
ADDHX1 inst_cellmath__66_0_I1617 (.CO(N6407), .S(N6389), .A(inst_cellmath__40[4]), .B(N6375));
INVXL inst_cellmath__66_0_I1618 (.Y(N6422), .A(inst_cellmath__40[5]));
NAND2X1 inst_cellmath__66_0_I1619 (.Y(N6395), .A(inst_cellmath__40[0]), .B(N6399));
AND2XL inst_cellmath__66_0_I1620 (.Y(N6412), .A(inst_cellmath__40[1]), .B(inst_delta[1]));
OR2XL inst_cellmath__66_0_I1621 (.Y(N6430), .A(inst_cellmath__40[1]), .B(inst_delta[1]));
NOR2X1 inst_cellmath__66_0_I1622 (.Y(N6370), .A(N6398), .B(N2396));
NAND2X1 inst_cellmath__66_0_I1623 (.Y(N6385), .A(N6398), .B(N2396));
NOR2X1 inst_cellmath__66_0_I1624 (.Y(N6400), .A(N6437), .B(N6423));
NAND2X1 inst_cellmath__66_0_I1625 (.Y(N6418), .A(N6437), .B(N6423));
NOR2XL inst_cellmath__66_0_I1626 (.Y(N6439), .A(N6389), .B(N6381));
NAND2X1 inst_cellmath__66_0_I1627 (.Y(N6376), .A(N6389), .B(N6381));
NOR2XL inst_cellmath__66_0_I1628 (.Y(N6391), .A(N6422), .B(N6407));
NAND2XL inst_cellmath__66_0_I1629 (.Y(N6408), .A(N6422), .B(N6407));
INVXL inst_cellmath__66_0_I1630 (.Y(N6377), .A(inst_cellmath__40[6]));
NOR2XL inst_cellmath__66_0_I1631 (.Y(N6425), .A(inst_cellmath__40[5]), .B(N6377));
NAND2XL inst_cellmath__66_0_I1632 (.Y(N6367), .A(inst_cellmath__40[5]), .B(N6377));
INVX1 inst_cellmath__66_0_I1633 (.Y(N6392), .A(N6395));
AOI21XL inst_cellmath__66_0_I1634 (.Y(N6372), .A0(N6430), .A1(N6395), .B0(N6412));
AOI21X1 inst_cellmath__66_0_I1635 (.Y(N6404), .A0(N6412), .A1(N6385), .B0(N6370));
NAND2XL inst_cellmath__66_0_I1636 (.Y(N6419), .A(N6385), .B(N6430));
AOI21XL inst_cellmath__66_0_I1637 (.Y(N6363), .A0(N6418), .A1(N6370), .B0(N6400));
NAND2XL inst_cellmath__66_0_I1638 (.Y(N6380), .A(N6418), .B(N6385));
AOI21X1 inst_cellmath__66_0_I1639 (.Y(N6396), .A0(N6376), .A1(N6400), .B0(N6439));
NAND2X1 inst_cellmath__66_0_I1640 (.Y(N6414), .A(N6376), .B(N6418));
AOI21XL inst_cellmath__66_0_I1641 (.Y(N6431), .A0(N6408), .A1(N6439), .B0(N6391));
NAND2XL inst_cellmath__66_0_I1642 (.Y(N6371), .A(N6408), .B(N6376));
AOI21XL inst_cellmath__66_0_I1643 (.Y(N6387), .A0(N6367), .A1(N6391), .B0(N6425));
NAND2XL inst_cellmath__66_0_I1644 (.Y(N6402), .A(N6367), .B(N6408));
INVXL inst_cellmath__66_0_I1645 (.Y(N6409), .A(N6392));
INVXL inst_cellmath__66_0_I1646 (.Y(N6424), .A(N6372));
OAI21XL inst_cellmath__66_0_I1647 (.Y(N6369), .A0(N6419), .A1(N6392), .B0(N6404));
OAI21XL inst_cellmath__66_0_I1648 (.Y(N6436), .A0(N6414), .A1(N6404), .B0(N6396));
NOR2XL inst_cellmath__66_0_I1649 (.Y(N6374), .A(N6414), .B(N6419));
OAI21XL inst_cellmath__66_0_I1650 (.Y(N6388), .A0(N6371), .A1(N6363), .B0(N6431));
NOR2XL inst_cellmath__66_0_I1651 (.Y(N6405), .A(N6371), .B(N6380));
OAI21XL inst_cellmath__66_0_I1652 (.Y(N6421), .A0(N6402), .A1(N6396), .B0(N6387));
NOR2XL inst_cellmath__66_0_I1653 (.Y(N6365), .A(N6402), .B(N6414));
OA21X1 inst_cellmath__66_0_I1654 (.Y(N6415), .A0(N6380), .A1(N6372), .B0(N6363));
AOI21XL inst_cellmath__66_0_I1655 (.Y(N6394), .A0(N6374), .A1(N6409), .B0(N6436));
AOI21XL inst_cellmath__66_0_I1656 (.Y(N6429), .A0(N6405), .A1(N6424), .B0(N6388));
AOI21XL inst_cellmath__66_0_I1657 (.Y(N6384), .A0(N6365), .A1(N6369), .B0(N6421));
NAND2BXL inst_cellmath__66_0_I1658 (.Y(N6362), .AN(N6412), .B(N6430));
NAND2BXL inst_cellmath__66_0_I1659 (.Y(N6413), .AN(N6370), .B(N6385));
NAND2BXL inst_cellmath__66_0_I1660 (.Y(N6386), .AN(N6400), .B(N6418));
NAND2BXL inst_cellmath__66_0_I1661 (.Y(N6361), .AN(N6439), .B(N6376));
NAND2BXL inst_cellmath__66_0_I1662 (.Y(N6411), .AN(N6391), .B(N6408));
NAND2BXL inst_cellmath__66_0_I1663 (.Y(N6382), .AN(N6425), .B(N6367));
XNOR2X1 inst_cellmath__66_0_I1664 (.Y(N6434), .A(inst_cellmath__40[7]), .B(N6377));
XNOR2X1 inst_cellmath__66_0_I1665 (.Y(inst_cellmath__66[0]), .A(inst_cellmath__40[0]), .B(N6399));
XNOR2X1 inst_cellmath__66_0_I1666 (.Y(inst_cellmath__66[1]), .A(N6409), .B(N6362));
XNOR2X1 inst_cellmath__66_0_I1667 (.Y(inst_cellmath__66[2]), .A(N6424), .B(N6413));
XNOR2X1 inst_cellmath__66_0_I1668 (.Y(inst_cellmath__66[3]), .A(N6369), .B(N6386));
XOR2XL inst_cellmath__66_0_I3368 (.Y(inst_cellmath__66[4]), .A(N6415), .B(N6361));
XOR2XL inst_cellmath__66_0_I1672 (.Y(inst_cellmath__66[6]), .A(N6382), .B(N6429));
XOR2XL inst_cellmath__66_0_I1673 (.Y(inst_cellmath__66[7]), .A(N6434), .B(N6384));
INVXL inst_cellmath__60_0_I1674 (.Y(N6512), .A(inst_cellmath__77));
XOR2XL inst_cellmath__60_0_I3286 (.Y(N6511), .A(N6411), .B(N6394));
INVX2 inst_cellmath__60_0_I1683 (.Y(N6518), .A(N8760));
AOI22XL inst_cellmath__60_0_I1684 (.Y(x[23]), .A0(N6518), .A1(inst_cellmath__66[0]), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1685 (.Y(x[24]), .A0(N6518), .A1(inst_cellmath__66[1]), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1686 (.Y(x[25]), .A0(N6518), .A1(inst_cellmath__66[2]), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1687 (.Y(x[26]), .A0(N6518), .A1(inst_cellmath__66[3]), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1688 (.Y(x[27]), .A0(N6518), .A1(inst_cellmath__66[4]), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1689 (.Y(x[28]), .A0(N6518), .A1(N6511), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1690 (.Y(x[29]), .A0(N6518), .A1(inst_cellmath__66[6]), .B0(N6512), .B1(N8760));
AOI22XL inst_cellmath__60_0_I1691 (.Y(x[30]), .A0(N6518), .A1(inst_cellmath__66[7]), .B0(N6512), .B1(N8760));
INVX8 inst_cellmath__63_0_I1693 (.Y(N6715), .A(inst_delta[3]));
AND2XL inst_cellmath__63_0_I1701 (.Y(N6559), .A(N6715), .B(inst_cellmath__51[3]));
AND2XL inst_cellmath__63_0_I1702 (.Y(N6637), .A(N6715), .B(inst_cellmath__51[4]));
AND2XL inst_cellmath__63_0_I1703 (.Y(N6712), .A(N6715), .B(inst_cellmath__51[5]));
AND2XL inst_cellmath__63_0_I1704 (.Y(N6613), .A(N6715), .B(inst_cellmath__51[6]));
AND2XL inst_cellmath__63_0_I1705 (.Y(N6688), .A(N6715), .B(inst_cellmath__51[7]));
MX2XL inst_cellmath__63_0_I1706 (.Y(N6592), .A(inst_cellmath__51[0]), .B(inst_cellmath__51[8]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1707 (.Y(N6630), .A(inst_cellmath__51[1]), .B(inst_cellmath__51[9]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1708 (.Y(N6666), .A(inst_cellmath__51[2]), .B(inst_cellmath__51[10]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1709 (.Y(N6705), .A(inst_cellmath__51[3]), .B(inst_cellmath__51[11]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1710 (.Y(N6569), .A(inst_cellmath__51[4]), .B(inst_cellmath__51[12]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1711 (.Y(N6608), .A(inst_cellmath__51[5]), .B(inst_cellmath__51[13]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1712 (.Y(N6647), .A(inst_cellmath__51[6]), .B(inst_cellmath__51[14]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1717 (.Y(N6661), .A(inst_cellmath__51[11]), .B(inst_cellmath__51[19]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1718 (.Y(N6700), .A(inst_cellmath__51[12]), .B(inst_cellmath__51[20]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1719 (.Y(N6564), .A(inst_cellmath__51[13]), .B(inst_cellmath__51[21]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1720 (.Y(N6602), .A(inst_cellmath__51[14]), .B(inst_cellmath__51[22]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1721 (.Y(N6642), .A(inst_cellmath__51[15]), .B(inst_cellmath__51[23]), .S0(N6715));
MX2XL inst_cellmath__63_0_I1722 (.Y(N6677), .A(inst_cellmath__51[16]), .B(inst_cellmath__51[24]), .S0(N6715));
AND2XL inst_cellmath__63_0_I8616 (.Y(N6679), .A(N6715), .B(inst_cellmath__51[0]));
CLKINVX6 inst_cellmath__63_0_I8623 (.Y(N6634), .A(inst_delta[4]));
NAND2XL inst_cellmath__63_0_I1728 (.Y(N6672), .A(N6679), .B(N6634));
AND2XL inst_cellmath__63_0_I8617 (.Y(N6581), .A(N6715), .B(inst_cellmath__51[1]));
NAND2XL inst_cellmath__63_0_I1729 (.Y(N6575), .A(N6581), .B(N6634));
AND2XL inst_cellmath__63_0_I8618 (.Y(N6658), .A(N6715), .B(inst_cellmath__51[2]));
NAND2XL inst_cellmath__63_0_I1730 (.Y(N6652), .A(N6658), .B(N6634));
NAND2XL inst_cellmath__63_0_I1731 (.Y(N6554), .A(N6559), .B(N6634));
NAND2XL inst_cellmath__63_0_I1732 (.Y(N6629), .A(N6637), .B(N6634));
NAND2XL inst_cellmath__63_0_I1733 (.Y(N6704), .A(N6712), .B(N6634));
NAND2XL inst_cellmath__63_0_I1734 (.Y(N6606), .A(N6613), .B(N6634));
NAND2XL inst_cellmath__63_0_I1735 (.Y(N6681), .A(N6688), .B(N6634));
NAND2XL inst_cellmath__63_0_I1736 (.Y(N6583), .A(N6592), .B(N6634));
NAND2XL inst_cellmath__63_0_I1737 (.Y(N6660), .A(N6630), .B(N6634));
NAND2XL inst_cellmath__63_0_I1738 (.Y(N6563), .A(N6666), .B(N6634));
NAND2XL inst_cellmath__63_0_I1739 (.Y(N6641), .A(N6705), .B(N6634));
NAND2XL inst_cellmath__63_0_I1740 (.Y(N6716), .A(N6634), .B(N6569));
NAND2XL inst_cellmath__63_0_I1741 (.Y(N6618), .A(N6634), .B(N6608));
NAND2XL inst_cellmath__63_0_I1742 (.Y(N6693), .A(N6647), .B(N6634));
MXI2X1 inst_cellmath__63_0_I1747 (.Y(N6611), .A(N6559), .B(N6661), .S0(N6634));
MXI2X1 inst_cellmath__63_0_I1748 (.Y(N6650), .A(N6637), .B(N6700), .S0(N6634));
MXI2XL inst_cellmath__63_0_I1749 (.Y(N6686), .A(N6712), .B(N6564), .S0(N6634));
MXI2XL inst_cellmath__63_0_I1750 (.Y(N6552), .A(N6613), .B(N6602), .S0(N6634));
MXI2XL inst_cellmath__63_0_I1751 (.Y(N6589), .A(N6688), .B(N6642), .S0(N6634));
MXI2XL inst_cellmath__63_0_I1752 (.Y(N6627), .A(N6592), .B(N6677), .S0(N6634));
BUFX4 inst_cellmath__63_0_I8628 (.Y(N6588), .A(inst_delta[0]));
NOR2XL inst_cellmath__63_0_I1754 (.Y(N6621), .A(N6672), .B(N6588));
MXI2XL inst_cellmath__63_0_I1755 (.Y(N6696), .A(N6575), .B(N6672), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1756 (.Y(N6561), .A(N6652), .B(N6575), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1757 (.Y(N6600), .A(N6554), .B(N6652), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1758 (.Y(N6639), .A(N6629), .B(N6554), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1759 (.Y(N6676), .A(N6704), .B(N6629), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1760 (.Y(N6713), .A(N6606), .B(N6704), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1761 (.Y(N6577), .A(N6681), .B(N6606), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1762 (.Y(N6616), .A(N6583), .B(N6681), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1763 (.Y(N6655), .A(N6660), .B(N6583), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1764 (.Y(N6691), .A(N6563), .B(N6660), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1765 (.Y(N6557), .A(N6641), .B(N6563), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1766 (.Y(N6593), .A(N6716), .B(N6641), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1767 (.Y(N6632), .A(N6618), .B(N6716), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1768 (.Y(N6669), .A(N6693), .B(N6618), .S0(N6588));
MX2XL inst_cellmath__63_0_I8619 (.Y(N14550), .A(inst_cellmath__51[7]), .B(inst_cellmath__51[15]), .S0(N6715));
NAND2XL inst_cellmath__63_0_I8624 (.Y(N6596), .A(N6634), .B(N14550));
MXI2XL inst_cellmath__63_0_I1769 (.Y(N6708), .A(N6596), .B(N6693), .S0(N6588));
MX2XL inst_cellmath__63_0_I8621 (.Y(N14570), .A(inst_cellmath__51[9]), .B(inst_cellmath__51[17]), .S0(N6715));
MXI2X1 inst_cellmath__63_0_I8626 (.Y(N6709), .A(N6581), .B(N14570), .S0(N6634));
MX2XL inst_cellmath__63_0_I8620 (.Y(N14560), .A(inst_cellmath__51[8]), .B(inst_cellmath__51[16]), .S0(N6715));
MXI2X1 inst_cellmath__63_0_I8625 (.Y(N6670), .A(N6679), .B(N14560), .S0(N6634));
MXI2X1 inst_cellmath__63_0_I1771 (.Y(N6610), .A(N6709), .B(N6670), .S0(N6588));
MX2XL inst_cellmath__63_0_I8622 (.Y(N14533), .A(inst_cellmath__51[10]), .B(inst_cellmath__51[18]), .S0(N6715));
MXI2X1 inst_cellmath__63_0_I8627 (.Y(N6573), .A(N6658), .B(N14533), .S0(N6634));
MXI2X1 inst_cellmath__63_0_I1773 (.Y(N6684), .A(N6611), .B(N6573), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1775 (.Y(N6587), .A(N6686), .B(N6650), .S0(N6588));
MXI2XL inst_cellmath__63_0_I1777 (.Y(N6663), .A(N6589), .B(N6552), .S0(N6588));
MXI2X1 inst_cellmath__63_0_I8480 (.Y(N6722), .A(N6650), .B(N6611), .S0(N6588));
MXI2XL inst_cellmath__63_0_I8481 (.Y(N6625), .A(N6552), .B(N6686), .S0(N6588));
MXI2XL inst_cellmath__63_0_I8482 (.Y(N14303), .A(N6627), .B(N6589), .S0(N6588));
OA21X1 inst_cellmath__63_0_I8724 (.Y(N14539), .A0(N14573), .A1(N6079), .B0(N14535));
MXI2X1 inst_cellmath__63_0_I8629 (.Y(N6572), .A(N6670), .B(N6596), .S0(N6588));
MXI2X1 inst_cellmath__63_0_I8630 (.Y(N6648), .A(N6573), .B(N6709), .S0(N6588));
INVX1 inst_cellmath__63_0_I8631 (.Y(N6579), .A(inst_delta[1]));
MXI2XL inst_cellmath__63_0_I8632 (.Y(N6585), .A(N6572), .B(N6648), .S0(N14539));
MXI2XL inst_cellmath__63_0_I8484 (.Y(N6662), .A(N6648), .B(N6722), .S0(N6579));
MXI2XL inst_cellmath__63_0_I8485 (.Y(N14319), .A(N6625), .B(N14303), .S0(N6579));
BUFX2 inst_cellmath__63_0_I8486 (.Y(N6635), .A(N2397));
INVXL inst_cellmath__63_0_I8487 (.Y(N14309), .A(N6635));
MX2XL inst_cellmath__63_0_I8488 (.Y(N14334), .A(N6662), .B(N14319), .S0(N14309));
INVXL inst_cellmath__63_0_I8489 (.Y(N6906), .A(inst_cellmath__62));
CLKBUFX6 inst_cellmath__63_0_I8492 (.Y(N6921), .A(N6348));
CLKINVX8 inst_cellmath__63_0_I8493 (.Y(N6888), .A(N6921));
MXI2XL inst_cellmath__63_0_I8494 (.Y(x[22]), .A(N14317), .B(N14334), .S0(N6888));
NAND2XL inst_cellmath__63_0_I1781 (.Y(N6695), .A(N6621), .B(N6579));
NAND2XL inst_cellmath__63_0_I1782 (.Y(N6598), .A(N6696), .B(N6579));
MXI2XL inst_cellmath__63_0_I1783 (.Y(N6673), .A(N6621), .B(N6561), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1784 (.Y(N6711), .A(N6696), .B(N6600), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1785 (.Y(N6576), .A(N6561), .B(N6639), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1786 (.Y(N6614), .A(N6600), .B(N6676), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1787 (.Y(N6653), .A(N6639), .B(N6713), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1788 (.Y(N6689), .A(N6676), .B(N6577), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1789 (.Y(N6555), .A(N6713), .B(N6616), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1790 (.Y(N6591), .A(N6577), .B(N6655), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1791 (.Y(N6631), .A(N6616), .B(N6691), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1792 (.Y(N6667), .A(N6655), .B(N6557), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1793 (.Y(N6706), .A(N6691), .B(N6593), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1794 (.Y(N6570), .A(N6557), .B(N6632), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1795 (.Y(N6607), .A(N6593), .B(N6669), .S0(N6579));
MXI2X1 inst_cellmath__63_0_I1796 (.Y(N6646), .A(N6632), .B(N6708), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1797 (.Y(N6683), .A(N6669), .B(N6572), .S0(N6579));
MXI2X1 inst_cellmath__63_0_I1798 (.Y(N6720), .A(N6708), .B(N6610), .S0(N6579));
MXI2X1 inst_cellmath__63_0_I1800 (.Y(N6623), .A(N6610), .B(N6684), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1802 (.Y(N6699), .A(N6684), .B(N6587), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1803 (.Y(N6565), .A(N6722), .B(N6625), .S0(N6579));
MXI2XL inst_cellmath__63_0_I1804 (.Y(N6603), .A(N6587), .B(N6663), .S0(N6579));
OR2XL inst_cellmath__63_0_I1809 (.Y(inst_cellmath__63[2]), .A(N6673), .B(N6635));
OR2XL inst_cellmath__63_0_I1810 (.Y(inst_cellmath__63[3]), .A(N6711), .B(N6635));
MX2XL inst_cellmath__63_0_I1811 (.Y(inst_cellmath__63[4]), .A(N6576), .B(N6695), .S0(N6635));
MX2XL inst_cellmath__63_0_I1812 (.Y(inst_cellmath__63[5]), .A(N6614), .B(N6598), .S0(N6635));
MX2XL inst_cellmath__63_0_I1814 (.Y(inst_cellmath__63[7]), .A(N6689), .B(N6711), .S0(N6635));
MX2XL inst_cellmath__63_0_I1815 (.Y(inst_cellmath__63[8]), .A(N6555), .B(N6576), .S0(N6635));
MX2XL inst_cellmath__63_0_I1816 (.Y(inst_cellmath__63[9]), .A(N6591), .B(N6614), .S0(N6635));
MX2XL inst_cellmath__63_0_I1817 (.Y(inst_cellmath__63[10]), .A(N6631), .B(N6653), .S0(N6635));
MX2XL inst_cellmath__63_0_I1818 (.Y(inst_cellmath__63[11]), .A(N6667), .B(N6689), .S0(N6635));
MX2XL inst_cellmath__63_0_I1819 (.Y(inst_cellmath__63[12]), .A(N6706), .B(N6555), .S0(N6635));
MX2XL inst_cellmath__63_0_I1820 (.Y(inst_cellmath__63[13]), .A(N6570), .B(N6591), .S0(N6635));
MX2XL inst_cellmath__63_0_I1821 (.Y(inst_cellmath__63[14]), .A(N6607), .B(N6631), .S0(N6635));
MX2XL inst_cellmath__63_0_I1822 (.Y(inst_cellmath__63[15]), .A(N6646), .B(N6667), .S0(N6635));
MX2XL inst_cellmath__63_0_I1823 (.Y(inst_cellmath__63[16]), .A(N6683), .B(N6706), .S0(N6635));
MX2XL inst_cellmath__63_0_I1824 (.Y(inst_cellmath__63[17]), .A(N6720), .B(N6570), .S0(N6635));
MX2XL inst_cellmath__63_0_I1825 (.Y(inst_cellmath__63[18]), .A(N6585), .B(N6607), .S0(N6635));
MX2XL inst_cellmath__63_0_I1826 (.Y(inst_cellmath__63[19]), .A(N6623), .B(N6646), .S0(N6635));
MX2XL inst_cellmath__63_0_I1827 (.Y(inst_cellmath__63[20]), .A(N6662), .B(N6683), .S0(N6635));
MX2XL inst_cellmath__63_0_I1828 (.Y(inst_cellmath__63[21]), .A(N6699), .B(N6720), .S0(N6635));
MX2XL inst_cellmath__63_0_I1829 (.Y(inst_cellmath__63[22]), .A(N6565), .B(N6585), .S0(N6635));
MX2XL inst_cellmath__63_0_I1830 (.Y(inst_cellmath__63[23]), .A(N6603), .B(N6623), .S0(N6635));
MX2XL cynw_cm_float_add2_I3280 (.Y(N6922), .A(N6653), .B(N6673), .S0(N6635));
AOI22XL cynw_cm_float_add2_I1858 (.Y(x[0]), .A0(N6888), .A1(inst_cellmath__63[2]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1859 (.Y(x[1]), .A0(N6888), .A1(inst_cellmath__63[3]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1860 (.Y(x[2]), .A0(N6888), .A1(inst_cellmath__63[4]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1861 (.Y(x[3]), .A0(N6888), .A1(inst_cellmath__63[5]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1862 (.Y(x[4]), .A0(N6888), .A1(N6922), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1863 (.Y(x[5]), .A0(N6888), .A1(inst_cellmath__63[7]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I3274 (.Y(x[6]), .A0(N6906), .A1(N6921), .B0(inst_cellmath__63[8]), .B1(N6888));
AOI22XL cynw_cm_float_add2_I1865 (.Y(x[7]), .A0(N6888), .A1(inst_cellmath__63[9]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1866 (.Y(x[8]), .A0(N6888), .A1(inst_cellmath__63[10]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1867 (.Y(x[9]), .A0(N6888), .A1(inst_cellmath__63[11]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1868 (.Y(x[10]), .A0(N6888), .A1(inst_cellmath__63[12]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1869 (.Y(x[11]), .A0(N6888), .A1(inst_cellmath__63[13]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1870 (.Y(x[12]), .A0(N6888), .A1(inst_cellmath__63[14]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1871 (.Y(x[13]), .A0(N6888), .A1(inst_cellmath__63[15]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1872 (.Y(x[14]), .A0(N6888), .A1(inst_cellmath__63[16]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1873 (.Y(x[15]), .A0(N6888), .A1(inst_cellmath__63[17]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1874 (.Y(x[16]), .A0(N6888), .A1(inst_cellmath__63[18]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1875 (.Y(x[17]), .A0(N6888), .A1(inst_cellmath__63[19]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1876 (.Y(x[18]), .A0(N6888), .A1(inst_cellmath__63[20]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1877 (.Y(x[19]), .A0(N6888), .A1(inst_cellmath__63[21]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1878 (.Y(x[20]), .A0(N6888), .A1(inst_cellmath__63[22]), .B0(N6906), .B1(N6921));
AOI22XL cynw_cm_float_add2_I1879 (.Y(x[21]), .A0(N6888), .A1(inst_cellmath__63[23]), .B0(N6906), .B1(N6921));
assign inst_cellmath__39[23] = 1'B0;
assign inst_cellmath__39[24] = 1'B0;
assign inst_cellmath__44[0] = 1'B0;
assign inst_cellmath__44[1] = 1'B0;
assign inst_cellmath__44[8] = 1'B0;
assign inst_cellmath__47[0] = 1'B0;
assign inst_cellmath__47[1] = 1'B0;
assign inst_cellmath__47[4] = 1'B0;
assign inst_cellmath__48[0] = 1'B0;
assign inst_cellmath__48[24] = 1'B1;
assign inst_cellmath__49[24] = 1'B0;
assign inst_delta[2] = 1'B0;
assign inst_cellmath__55[23] = 1'B0;
assign inst_cellmath__56[0] = 1'B0;
assign inst_cellmath__56[1] = 1'B0;
assign inst_cellmath__56[2] = 1'B0;
assign inst_cellmath__56[3] = 1'B0;
assign inst_cellmath__56[4] = 1'B0;
assign inst_cellmath__56[5] = 1'B0;
assign inst_cellmath__56[6] = 1'B0;
assign inst_cellmath__56[7] = 1'B0;
assign inst_cellmath__56[8] = 1'B0;
assign inst_cellmath__56[9] = 1'B0;
assign inst_cellmath__56[10] = 1'B0;
assign inst_cellmath__56[11] = 1'B0;
assign inst_cellmath__56[12] = 1'B0;
assign inst_cellmath__56[13] = 1'B0;
assign inst_cellmath__56[14] = 1'B0;
assign inst_cellmath__56[15] = 1'B0;
assign inst_cellmath__56[16] = 1'B0;
assign inst_cellmath__56[17] = 1'B0;
assign inst_cellmath__56[18] = 1'B0;
assign inst_cellmath__56[19] = 1'B0;
assign inst_cellmath__56[20] = 1'B0;
assign inst_cellmath__56[21] = 1'B0;
assign inst_cellmath__56[22] = 1'B0;
assign inst_cellmath__56[23] = 1'B0;
assign inst_cellmath__56[24] = 1'B0;
assign inst_cellmath__63[0] = 1'B0;
assign inst_cellmath__63[1] = 1'B0;
assign inst_cellmath__63[6] = 1'B0;
assign inst_cellmath__63[24] = 1'B0;
assign inst_cellmath__66[5] = 1'B0;
endmodule

/* CADENCE  urL2QwjWrxk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




