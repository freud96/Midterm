/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:23:19 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__68,
	inst_cellmath__82;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire  inst_cellmath__219;
wire N487,N541,N542,N543,N544,N577,N578 
	,N579,N580,N608,N609,N610,N611,N612,N613 
	,N614,N615,N616,N617,N618,N619,N620,N621 
	,N622,N623,N624,N625,N626,N627,N628,N629 
	,N630,N631,N632,N633,N634,N635,N636,N637 
	,N639,N640,N641,N642,N643,N644,N645,N646 
	,N647,N648,N649,N650,N651,N652,N653,N654 
	,N655,N656,N657,N658,N659,N660,N661,N662 
	,N663,N664,N665,N666,N667,N668,N669,N670 
	,N679,N680,N681,N682,N683,N684,N685,N686 
	,N687,N688,N689,N690,N691,N692,N693,N694 
	,N695,N696,N697,N698,N699,N700,N701,N733 
	,N734,N735,N736,N737,N738,N739,N740,N741 
	,N742,N743,N744,N745,N746,N747,N748,N749 
	,N750,N751,N752,N753,N754,N755,N757,N759 
	,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923 
	,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934 
	,N3935,N3936,N3937,N3938,N3940,N3941,N3942,N3943 
	,N3944,N3945,N3946,N3948,N3949,N3951,N3952,N3953 
	,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961 
	,N3962,N3963,N3966,N3967,N3968,N3969,N3970,N3971 
	,N3972,N3973,N3975,N3976,N3977,N3978,N3979,N3981 
	,N3982,N3983,N3984,N3985,N3987,N3988,N3989,N3990 
	,N3991,N3992,N3994,N3995,N3996,N3997,N3998,N3999 
	,N4000,N4001,N4004,N4005,N4006,N4007,N4008,N4010 
	,N4011,N4012,N4013,N4014,N4015,N4016,N4019,N4020 
	,N4021,N4022,N4023,N4024,N4025,N4026,N4028,N4029 
	,N4030,N4031,N4032,N4034,N4035,N4036,N4037,N4038 
	,N4039,N4040,N4041,N4042,N4045,N4046,N4047,N4048 
	,N4049,N4050,N4052,N4053,N4054,N4055,N4056,N4058 
	,N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066 
	,N4068,N4069,N4071,N4072,N4073,N4074,N4075,N4076 
	,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085 
	,N4086,N4087,N4088,N4090,N4092,N4093,N4095,N4096 
	,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104 
	,N4106,N4107,N4109,N4110,N4111,N4112,N4113,N4114 
	,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122 
	,N4124,N4125,N4128,N4129,N4130,N4131,N4132,N4133 
	,N4134,N4137,N4138,N4139,N4140,N4141,N4143,N4144 
	,N4145,N4146,N4148,N4149,N4150,N4152,N4153,N4154 
	,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162 
	,N4164,N4165,N4166,N4167,N4168,N4169,N4170,N4173 
	,N4174,N4175,N4176,N4177,N4178,N4180,N4181,N4182 
	,N4183,N4184,N4185,N4187,N4188,N4189,N4190,N4191 
	,N4192,N4193,N4194,N4196,N4197,N4198,N4199,N4200 
	,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208 
	,N4209,N4210,N4212,N4213,N4214,N4215,N4217,N4218 
	,N4219,N4220,N4221,N4222,N4224,N4225,N4226,N4227 
	,N4228,N4229,N4230,N4231,N4232,N4233,N4235,N4236 
	,N4237,N4238,N4239,N4240,N4241,N4243,N4244,N4245 
	,N4246,N4247,N4249,N4251,N4253,N4254,N4255,N4256 
	,N4257,N4258,N4259,N4262,N4263,N4265,N4266,N4267 
	,N4268,N4269,N4270,N4271,N4273,N4274,N4275,N4276 
	,N4277,N4278,N4280,N4281,N4282,N4283,N4284,N4285 
	,N4287,N4288,N4289,N4291,N4292,N4293,N4294,N4295 
	,N4296,N4297,N4299,N4300,N4301,N4302,N4303,N4305 
	,N4306,N4307,N4308,N4309,N4312,N4313,N4314,N4316 
	,N4317,N4318,N4319,N4320,N4321,N4322,N4324,N4326 
	,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334 
	,N4335,N4336,N4338,N4339,N4342,N4343,N4344,N4346 
	,N4347,N4348,N4349,N4350,N4351,N4352,N4354,N4355 
	,N4356,N4359,N4360,N4361,N4362,N4363,N4364,N4365 
	,N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4374 
	,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382 
	,N4383,N4385,N4386,N4387,N4389,N4390,N4392,N4393 
	,N4394,N4396,N4397,N4398,N4400,N4401,N4402,N4403 
	,N4404,N4405,N4406,N4408,N4409,N4410,N4411,N4412 
	,N4413,N4414,N4415,N4416,N4417,N4418,N4420,N4421 
	,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429 
	,N4430,N4431,N4432,N4434,N4435,N4436,N4437,N4438 
	,N4439,N4440,N4441,N4442,N4443,N4446,N4447,N4449 
	,N4450,N4451,N4453,N4454,N4455,N4456,N4457,N4459 
	,N4461,N4462,N4463,N4464,N4465,N4467,N4468,N4469 
	,N4471,N4472,N4473,N4476,N4477,N4478,N4479,N4480 
	,N4481,N4482,N4483,N4484,N4486,N4487,N4488,N4489 
	,N4490,N4491,N4492,N4493,N4494,N4496,N4497,N4498 
	,N4499,N4501,N4502,N4503,N4504,N4505,N4507,N4508 
	,N4509,N4510,N4512,N4513,N4515,N4516,N4517,N4518 
	,N4519,N4520,N4521,N4523,N4524,N4525,N4526,N4528 
	,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4537 
	,N4538,N4539,N4540,N4542,N4543,N4545,N4546,N4548 
	,N4549,N4550,N4551,N4552,N4554,N4556,N4557,N4558 
	,N4559,N4560,N4562,N4563,N4564,N4565,N4567,N4569 
	,N4570,N4571,N4573,N4574,N4575,N4577,N4578,N4579 
	,N4580,N4582,N4583,N4584,N4585,N4586,N4587,N4588 
	,N4589,N4590,N4591,N4592,N4594,N4595,N4596,N4597 
	,N4598,N4600,N4601,N4602,N4604,N4605,N4606,N4607 
	,N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615 
	,N4617,N4618,N4619,N4621,N4622,N4623,N4624,N4626 
	,N4628,N4630,N4631,N4632,N4633,N4634,N4635,N4636 
	,N4637,N4638,N4640,N4641,N5345,N5347,N5348,N5349 
	,N5360,N5373,N5374,N5375,N5377,N5378,N5379,N5381 
	,N5382,N5383,N5385,N5386,N5388,N5389,N5390,N5392 
	,N5394,N5395,N5397,N5399,N5400,N5401,N5402,N5404 
	,N5406,N5407,N5408,N5409,N5410,N5411,N5413,N5414 
	,N5415,N5417,N5418,N5420,N5421,N5422,N5424,N5425 
	,N5427,N5428,N5429,N5430,N5432,N5433,N5434,N5436 
	,N5437,N5439,N5441,N5442,N5443,N5446,N5447,N5448 
	,N5449,N5451,N5453,N5454,N5455,N5456,N5457,N5459 
	,N5460,N5462,N5463,N5465,N5467,N5468,N5470,N5472 
	,N5473,N5474,N5476,N5477,N5478,N5480,N5481,N5483 
	,N5485,N5486,N5488,N5489,N5490,N5492,N5493,N5494 
	,N5495,N5497,N5499,N5500,N5501,N5502,N5504,N5505 
	,N5506,N5508,N5509,N5511,N5513,N5514,N5515,N5516 
	,N5519,N5520,N5521,N5522,N5524,N5525,N5527,N5528 
	,N5529,N5530,N5531,N5533,N5534,N5536,N5537,N5539 
	,N5540,N5541,N5542,N5544,N5545,N5547,N5548,N5549 
	,N5550,N5552,N5553,N5555,N5556,N5558,N5560,N5561 
	,N5562,N5565,N5566,N5567,N5568,N5570,N5571,N5573 
	,N5574,N5575,N5576,N5578,N5579,N5580,N5581,N5583 
	,N5584,N5586,N5778,N5837,N5838,N5839,N5840,N5842 
	,N5843,N5845,N5846,N5847,N5848,N5850,N5851,N5852 
	,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860 
	,N5861,N5862,N5863,N5865,N5866,N5867,N5868,N5869 
	,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5878 
	,N5879,N5881,N5882,N5883,N5884,N5885,N5886,N5887 
	,N5888,N5889,N5890,N5891,N5892,N5893,N5894,N5895 
	,N5897,N5898,N5899,N5900,N5901,N5902,N5903,N5905 
	,N5906,N5907,N5908,N5909,N5911,N5912,N5913,N5914 
	,N5916,N5917,N5918,N5919,N5920,N5921,N5922,N5923 
	,N5924,N5925,N5926,N5927,N5928,N5929,N5931,N5932 
	,N5933,N5935,N5936,N5937,N5938,N5939,N5940,N5941 
	,N5942,N5943,N5944,N5945,N5946,N5947,N5948,N5950 
	,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958 
	,N5959,N5960,N5961,N5963,N5964,N5965,N5966,N5969 
	,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977 
	,N5978,N5979,N5980,N5981,N5982,N5984,N5986,N5987 
	,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995 
	,N5997,N5998,N6000,N6001,N6002,N6003,N6004,N6005 
	,N6006,N6007,N6008,N6009,N6010,N6012,N6014,N6015 
	,N6016,N6017,N6018,N6019,N6020,N6021,N6022,N6023 
	,N6024,N6026,N6027,N6028,N6029,N6030,N6031,N6032 
	,N6033,N6034,N6036,N6037,N6038,N6039,N6040,N6041 
	,N6042,N6043,N6044,N6045,N6047,N6050,N6051,N6052 
	,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060 
	,N6061,N6062,N6063,N6064,N6066,N6067,N6069,N6070 
	,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078 
	,N6079,N6080,N6082,N6083,N6084,N6085,N6086,N6087 
	,N6088,N6089,N6090,N6092,N6093,N6094,N6095,N6096 
	,N6098,N6099,N6102,N6103,N6104,N6105,N6106,N6107 
	,N6108,N6109,N6110,N6111,N6112,N6114,N6115,N6116 
	,N6117,N6118,N6119,N6120,N6121,N6123,N6124,N6125 
	,N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133 
	,N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142 
	,N6144,N6145,N6146,N6147,N6149,N6150,N6151,N6152 
	,N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160 
	,N6161,N6162,N6164,N6165,N6166,N6167,N6168,N6169 
	,N6170,N6171,N6172,N6173,N6174,N6175,N6178,N6180 
	,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188 
	,N6189,N6191,N6192,N6193,N6195,N6196,N6197,N6198 
	,N6199,N6200,N6201,N6202,N6203,N6206,N6208,N6209 
	,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218 
	,N6219,N6220,N6221,N6222,N6223,N6225,N6226,N6227 
	,N6228,N6229,N6230,N6231,N6232,N6233,N6234,N6236 
	,N6237,N6239,N6241,N6242,N6243,N6244,N6245,N6247 
	,N6248,N6249,N6250,N6251,N6252,N6253,N6254,N6255 
	,N6257,N6258,N6260,N6261,N6262,N6263,N6264,N6265 
	,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6274 
	,N6275,N6276,N6277,N6278,N6279,N6280,N6281,N6282 
	,N6284,N6285,N6287,N6288,N6289,N6291,N6292,N6293 
	,N6294,N6295,N6296,N6297,N6298,N6299,N6300,N6301 
	,N6302,N6304,N6305,N6306,N6307,N6308,N6309,N6310 
	,N6311,N6312,N6313,N6314,N6315,N6316,N6317,N6318 
	,N6319,N6321,N6322,N6323,N6324,N6325,N6326,N6327 
	,N6328,N6329,N6331,N6332,N6334,N6335,N6336,N6338 
	,N6339,N6340,N6341,N6342,N6343,N6344,N6345,N6346 
	,N6347,N6350,N6351,N6352,N6353,N6354,N6355,N6356 
	,N6357,N6358,N6359,N6361,N6362,N6364,N6365,N6366 
	,N6367,N6368,N6370,N6371,N6372,N6373,N6374,N6375 
	,N6376,N6377,N6378,N6379,N6380,N6382,N6383,N6385 
	,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393 
	,N6395,N6396,N6397,N6399,N6400,N6401,N6402,N6403 
	,N6404,N6406,N6407,N6408,N6409,N6411,N6413,N6414 
	,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422 
	,N6423,N6424,N6425,N6426,N6428,N6429,N6430,N6432 
	,N6433,N6434,N6435,N6436,N6437,N6438,N6439,N6440 
	,N6441,N6442,N6443,N6444,N6446,N6447,N6448,N6449 
	,N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457 
	,N6458,N6460,N6461,N6464,N6465,N6466,N6467,N6468 
	,N6470,N6471,N6472,N6473,N6474,N6476,N6477,N6478 
	,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486 
	,N6487,N6488,N6490,N6491,N6492,N6493,N6494,N6496 
	,N6497,N6498,N6499,N6500,N6502,N6503,N6504,N6505 
	,N6507,N6508,N6509,N6510,N6511,N6512,N6513,N6514 
	,N6517,N6518,N6519,N6520,N6521,N6522,N6523,N6524 
	,N6525,N6526,N6527,N6530,N6532,N6533,N6534,N6535 
	,N6536,N6537,N6538,N6540,N6541,N6542,N6543,N6544 
	,N6545,N6547,N6548,N6549,N6550,N6551,N6552,N6553 
	,N6554,N6555,N6556,N6557,N6558,N6560,N6562,N6563 
	,N6565,N6566,N6567,N6568,N6569,N6570,N6571,N6572 
	,N6573,N6574,N6576,N6577,N6578,N6580,N6582,N6583 
	,N6584,N6585,N6586,N6587,N6588,N6589,N6590,N6591 
	,N6592,N6595,N6596,N6597,N6598,N6599,N6600,N6601 
	,N6603,N6604,N6605,N6606,N6608,N6609,N6610,N6611 
	,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620 
	,N6621,N6622,N6623,N6625,N6626,N6628,N6629,N6630 
	,N6631,N6633,N6634,N6635,N6636,N6638,N6639,N6640 
	,N6641,N6643,N6645,N6646,N6647,N6648,N6649,N6650 
	,N6651,N6653,N6654,N6655,N6658,N6659,N6660,N6661 
	,N6662,N6663,N6664,N6665,N6666,N6667,N6668,N6669 
	,N6670,N6671,N6672,N6673,N6674,N6676,N6677,N6678 
	,N7515,N7516,N7517,N7518,N7520,N7521,N7522,N7523 
	,N7524,N7526,N7527,N7528,N7529,N7530,N7531,N7532 
	,N7533,N7534,N7536,N7537,N7538,N7539,N7540,N7541 
	,N7542,N7543,N7544,N7545,N7546,N7548,N7549,N7550 
	,N7551,N7552,N7553,N7554,N7555,N7556,N7557,N7558 
	,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567 
	,N7568,N7569,N7570,N7571,N7572,N7573,N7574,N7575 
	,N7576,N7577,N7578,N7579,N7580,N7582,N7583,N7584 
	,N7586,N7587,N7588,N7589,N7591,N7592,N7593,N7594 
	,N7595,N7596,N7597,N7598,N7599,N7600,N7601,N7602 
	,N7604,N7605,N7606,N7608,N7609,N7610,N7611,N7612 
	,N7613,N7615,N7616,N7617,N7618,N7619,N7620,N7621 
	,N7622,N7623,N7624,N7626,N7627,N7628,N7630,N7631 
	,N7633,N7634,N7635,N7636,N7637,N7639,N7641,N7642 
	,N7643,N7644,N7645,N7646,N7648,N7649,N7650,N7651 
	,N7652,N7654,N7655,N7656,N7657,N7660,N7662,N7664 
	,N7665,N7667,N7668,N7669,N7670,N7672,N7673,N7674 
	,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7683 
	,N7684,N7685,N7686,N7687,N7689,N7690,N7691,N7692 
	,N7693,N7694,N7695,N7696,N7697,N7698,N7699,N7700 
	,N7701,N7702,N7703,N7704,N7705,N7706,N7708,N7709 
	,N7710,N7711,N7712,N7713,N7714,N7715,N7716,N7718 
	,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726 
	,N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7736 
	,N7737,N7738,N7741,N7742,N7743,N7744,N7745,N7747 
	,N7748,N7749,N7750,N7751,N7752,N7753,N7754,N7755 
	,N7756,N7757,N7759,N7760,N7761,N7762,N7764,N7765 
	,N7766,N7767,N7768,N7769,N7770,N7771,N7772,N7773 
	,N7774,N7776,N7777,N7778,N7779,N7780,N7782,N7783 
	,N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792 
	,N7793,N7794,N7795,N7796,N7797,N7798,N7799,N7800 
	,N7801,N7802,N7803,N7804,N7806,N7807,N7808,N7809 
	,N7810,N7811,N7813,N7814,N7815,N7816,N7817,N7818 
	,N7819,N7820,N7821,N7822,N7823,N7824,N7825,N7826 
	,N7828,N7829,N7830,N7832,N7833,N7834,N7836,N7838 
	,N7839,N7840,N7841,N7842,N7843,N7844,N7846,N7847 
	,N7848,N7849,N7850,N7851,N7853,N7855,N7858,N7859 
	,N7860,N7861,N7862,N7864,N7865,N7866,N7867,N7868 
	,N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876 
	,N7877,N7878,N7880,N7881,N7882,N7883,N7884,N7885 
	,N7886,N7887,N7888,N7889,N7890,N7891,N7892,N7894 
	,N7895,N7896,N7897,N7898,N7900,N7901,N7902,N7903 
	,N7905,N7906,N7907,N7909,N7910,N7911,N7912,N7913 
	,N7914,N7915,N7916,N7918,N7919,N7920,N7921,N7922 
	,N7923,N7924,N7925,N7926,N7927,N7929,N7930,N7931 
	,N7932,N7933,N7934,N7935,N7936,N7937,N7938,N7939 
	,N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947 
	,N7948,N7949,N7951,N7952,N7953,N7954,N7955,N7956 
	,N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7965 
	,N7966,N7967,N7968,N7970,N7971,N7972,N7973,N7974 
	,N7975,N7976,N7977,N7978,N7981,N7982,N7983,N7984 
	,N7986,N7987,N7989,N7990,N7991,N7992,N7993,N7994 
	,N7995,N7996,N7997,N7998,N8000,N8001,N8002,N8003 
	,N8005,N8006,N8007,N8009,N8010,N8011,N8012,N8013 
	,N8014,N8015,N8016,N8017,N8019,N8020,N8021,N8024 
	,N8025,N8026,N8027,N8029,N8030,N8031,N8033,N8034 
	,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042 
	,N8043,N8044,N8045,N8046,N8047,N8048,N8049,N8052 
	,N8053,N8054,N8056,N8057,N8058,N8059,N8060,N8061 
	,N8062,N8064,N8065,N8066,N8067,N8068,N8069,N8070 
	,N8072,N8073,N8074,N8075,N8076,N8077,N8078,N8081 
	,N8082,N8083,N8084,N8086,N8088,N8089,N8648,N8649 
	,N8650,N8651,N8652,N8654,N8655,N8656,N8657,N8658 
	,N8659,N8660,N8661,N8662,N8663,N8664,N8665,N8666 
	,N8667,N8668,N8669,N8670,N8671,N8672,N8673,N8675 
	,N8676,N8677,N8678,N8679,N8680,N8681,N8683,N8685 
	,N8686,N8687,N8688,N8689,N8690,N8691,N8692,N8693 
	,N8694,N8695,N8696,N8697,N8699,N8700,N8701,N8702 
	,N8704,N8705,N8707,N8708,N8709,N8710,N8711,N8712 
	,N8713,N8714,N8715,N8716,N8717,N8718,N8719,N8720 
	,N8721,N8723,N8725,N8726,N8727,N8728,N8729,N8730 
	,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738 
	,N8740,N8741,N8742,N8743,N8744,N8745,N8746,N8748 
	,N8749,N8750,N8751,N8752,N8755,N8756,N8757,N8758 
	,N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766 
	,N8767,N8768,N8769,N8770,N8771,N8773,N8774,N8775 
	,N8776,N8777,N8778,N8780,N8781,N8782,N8783,N8784 
	,N8785,N8786,N8787,N8789,N8791,N8792,N8793,N8794 
	,N8795,N8796,N8797,N8798,N8800,N8801,N8802,N8803 
	,N8804,N8805,N8806,N8809,N8810,N8811,N8812,N8813 
	,N8814,N8815,N8816,N8817,N8818,N8819,N8820,N8821 
	,N8822,N8823,N8824,N8826,N8827,N8828,N8830,N8832 
	,N8833,N8834,N8835,N8836,N8837,N8838,N8839,N8840 
	,N8841,N8842,N8843,N8844,N8845,N8846,N8847,N8848 
	,N8849,N8850,N8851,N8852,N8853,N8854,N8855,N8857 
	,N8858,N8859,N8860,N8861,N8862,N8863,N8865,N8866 
	,N8867,N8868,N8869,N8870,N8872,N8873,N8874,N8875 
	,N8876,N8877,N8878,N8879,N8880,N8881,N8882,N8883 
	,N8884,N8886,N8887,N8888,N8890,N8892,N8893,N8894 
	,N8895,N8896,N8897,N8898,N8899,N8901,N8902,N8903 
	,N8904,N8905,N8906,N8907,N8908,N8909,N8910,N8911 
	,N8912,N8914,N8915,N8916,N8917,N8919,N8920,N8921 
	,N8922,N8923,N8924,N8925,N8926,N8927,N8928,N8929 
	,N8930,N8932,N8933,N8934,N8935,N8936,N8937,N8938 
	,N8939,N8940,N8941,N8942,N8943,N8945,N8946,N8947 
	,N8950,N8951,N8952,N8953,N8954,N8955,N8956,N8957 
	,N8958,N8959,N8960,N8961,N8962,N8963,N8964,N8965 
	,N8966,N8967,N8968,N8969,N8970,N8971,N8972,N8974 
	,N8975,N8976,N8977,N8978,N8980,N8981,N8982,N8983 
	,N8984,N8985,N8986,N8987,N8988,N8989,N8990,N8991 
	,N8992,N8993,N8994,N8995,N8996,N8997,N8998,N8999 
	,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007 
	,N9008,N9010,N9011,N9012,N9013,N9015,N9016,N9017 
	,N9018,N9019,N9021,N9022,N9023,N9024,N9025,N9026 
	,N9027,N9028,N9029,N9030,N9031,N9032,N9033,N9035 
	,N9036,N9037,N9039,N9040,N9042,N9043,N9044,N9045 
	,N9046,N9047,N9048,N9049,N9050,N9051,N9052,N9053 
	,N9054,N9055,N9056,N9057,N9058,N9059,N9060,N9061 
	,N9062,N9064,N9065,N9066,N9067,N9068,N9069,N9070 
	,N9071,N9072,N9073,N9074,N9075,N9076,N9077,N9078 
	,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087 
	,N9088,N9089,N9090,N9091,N9092,N9093,N9094,N9095 
	,N9097,N9098,N9099,N9101,N9102,N9103,N9104,N9105 
	,N9106,N9107,N9108,N9109,N9110,N9111,N9112,N9113 
	,N9114,N9115,N9116,N9117,N9118,N9119,N9120,N9121 
	,N9122,N9123,N9125,N9126,N9127,N9128,N9129,N9130 
	,N9131,N9133,N9134,N9135,N9136,N9137,N9138,N9139 
	,N9140,N9142,N9143,N9144,N9145,N9146,N9147,N9148 
	,N9149,N9150,N9151,N9152,N9153,N9154,N9155,N9156 
	,N9157,N9158,N9160,N9161,N9162,N9163,N9164,N9165 
	,N9167,N9169,N9170,N9171,N9172,N9173,N9174,N9175 
	,N9176,N9177,N9178,N9179,N9180,N9181,N9182,N9183 
	,N9184,N9185,N9186,N9187,N9188,N9190,N9191,N9192 
	,N9193,N9194,N9195,N9196,N9198,N9200,N9201,N9202 
	,N9203,N9204,N9205,N9206,N9207,N9208,N9209,N9210 
	,N9211,N9212,N9213,N9215,N9216,N9217,N9218,N9219 
	,N9220,N9221,N9222,N9223,N9224,N9225,N9227,N9228 
	,N9229,N9230,N9231,N9234,N9235,N9236,N9237,N9238 
	,N9240,N9241,N9243,N9244,N9245,N9246,N9247,N9248 
	,N9249,N9250,N9251,N9252,N9253,N9254,N9256,N9257 
	,N9258,N9259,N9260,N9261,N9263,N9265,N9266,N9267 
	,N9268,N9269,N9270,N9271,N9272,N9273,N9274,N9275 
	,N9276,N9277,N9278,N9279,N9280,N9281,N9283,N9284 
	,N9285,N9286,N9287,N9288,N9289,N9291,N9292,N9293 
	,N9294,N9295,N9296,N9297,N9298,N9299,N9300,N9301 
	,N9302,N9304,N9305,N9306,N9307,N9308,N9309,N9310 
	,N9311,N9312,N9313,N9314,N9315,N9316,N9317,N9318 
	,N9319,N9320,N9321,N9322,N9324,N9325,N9326,N9327 
	,N9328,N9329,N9330,N9333,N9334,N9335,N9336,N9337 
	,N9338,N9339,N9340,N9341,N9342,N9343,N9344,N9345 
	,N9346,N9347,N9348,N9349,N9351,N9352,N9353,N9354 
	,N9355,N9356,N9357,N9359,N9360,N9361,N9362,N9363 
	,N9364,N9365,N9366,N9367,N9368,N9369,N9370,N9372 
	,N9373,N9374,N9375,N9376,N9377,N9378,N9379,N9380 
	,N9381,N9382,N9383,N9384,N9385,N9386,N9387,N9389 
	,N9390,N9391,N9392,N9393,N9394,N9395,N9396,N9397 
	,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407 
	,N9408,N9409,N9410,N9411,N9412,N9413,N9414,N9415 
	,N9417,N9418,N9419,N9420,N9421,N9423,N9424,N9426 
	,N9427,N9428,N9429,N9430,N9431,N9432,N9433,N9434 
	,N9435,N9436,N9437,N9438,N9439,N9440,N9441,N9442 
	,N9443,N9444,N9446,N9447,N9448,N9449,N9450,N9451 
	,N9452,N9454,N9455,N9456,N9457,N9458,N9459,N9460 
	,N9462,N9463,N9464,N9465,N9467,N9468,N9469,N9470 
	,N9471,N9472,N9473,N9474,N9475,N9476,N9477,N9478 
	,N9479,N9480,N9481,N9482,N9484,N9485,N9486,N9487 
	,N9488,N9489,N9490,N9492,N9493,N9494,N9495,N9496 
	,N9497,N9498,N9499,N9501,N9502,N9503,N9504,N9505 
	,N9506,N9507,N9508,N9509,N9510,N9511,N9512,N9513 
	,N9514,N9516,N9517,N9518,N9519,N9520,N9521,N9522 
	,N9524,N9525,N9526,N9527,N9528,N9529,N9530,N9531 
	,N9532,N9533,N9536,N9537,N9538,N9539,N9540,N9541 
	,N9542,N9543,N9544,N9545,N9546,N9547,N9548,N9549 
	,N9550,N9551,N9552,N9554,N9555,N9556,N9557,N9558 
	,N9559,N9562,N9563,N9564,N9565,N9566,N9567,N9568 
	,N9569,N9570,N9571,N9572,N9573,N9574,N9575,N9576 
	,N9577,N9579,N9580,N9581,N9582,N9583,N9585,N9586 
	,N9587,N9589,N9590,N9591,N9592,N9593,N9594,N9595 
	,N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603 
	,N9604,N9605,N9606,N9607,N9608,N9609,N9610,N9611 
	,N9612,N9613,N9614,N9615,N9617,N9618,N9619,N9620 
	,N9621,N9623,N9624,N9625,N9627,N9628,N9629,N9631 
	,N9632,N9633,N9634,N9635,N9636,N9637,N9638,N9639 
	,N9640,N9641,N9642,N9643,N9644,N9645,N9647,N9648 
	,N9649,N9650,N9651,N9653,N9654,N9655,N9657,N9658 
	,N9659,N9660,N9661,N9662,N9663,N9664,N9665,N9666 
	,N9667,N9668,N9669,N9670,N9671,N9672,N9673,N9674 
	,N9676,N9677,N9678,N9679,N9680,N9681,N9682,N9683 
	,N9684,N9685,N9686,N9687,N9688,N9689,N9690,N9691 
	,N9692,N9693,N9694,N9695,N9697,N9698,N9699,N9700 
	,N9701,N9702,N9703,N9704,N9705,N9706,N9707,N9708 
	,N9709,N9710,N9711,N9712,N9714,N9715,N9716,N9717 
	,N9718,N9719,N9720,N9722,N9724,N9725,N9726,N9727 
	,N9728,N9729,N9730,N9731,N9732,N9733,N9734,N9735 
	,N9736,N9737,N9738,N9739,N9740,N9741,N9742,N9744 
	,N9745,N9746,N9747,N9748,N9749,N9750,N9752,N9753 
	,N9754,N9755,N9756,N9757,N9758,N9759,N9760,N9761 
	,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769 
	,N9770,N9771,N9772,N9773,N9774,N9776,N9777,N9778 
	,N9779,N9780,N9781,N9782,N9784,N9786,N9787,N9788 
	,N9789,N9790,N9791,N9792,N9793,N9794,N9795,N9796 
	,N9797,N9798,N9799,N9800,N9801,N9802,N9804,N9805 
	,N9806,N9807,N9808,N9810,N9811,N9813,N9814,N9815 
	,N9816,N9817,N9818,N9819,N9820,N9821,N9823,N9824 
	,N9825,N9826,N9827,N9828,N9829,N9831,N9832,N9833 
	,N9834,N9835,N9836,N9837,N9838,N9840,N9841,N9842 
	,N9843,N9844,N9845,N9846,N9847,N9848,N9850,N9851 
	,N9852,N9853,N9854,N9856,N9857,N9858,N9859,N9860 
	,N9861,N9862,N9863,N9864,N9865,N9866,N9868,N9869 
	,N9870,N9871,N9872,N9873,N9874,N9876,N9877,N9878 
	,N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886 
	,N9887,N9888,N9889,N9890,N9891,N9893,N9894,N9895 
	,N9896,N9897,N9898,N9899,N9901,N9902,N9903,N9904 
	,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9912 
	,N9913,N9914,N9915,N9917,N9918,N9919,N9920,N9921 
	,N9922,N9923,N9924,N9925,N9926,N9927,N9928,N9930 
	,N9931,N9932,N9933,N9934,N9935,N9936,N9939,N9940 
	,N9941,N9942,N9943,N9944,N9945,N9946,N9947,N9948 
	,N9949,N9950,N9951,N9952,N9953,N9954,N9955,N9956 
	,N9958,N9959,N9960,N9961,N9962,N9964,N9965,N9966 
	,N9967,N9968,N9969,N9970,N9971,N9972,N9973,N9974 
	,N9975,N9976,N9977,N9978,N9979,N9980,N9981,N9982 
	,N9983,N9984,N9985,N9986,N9988,N9989,N9990,N9991 
	,N9992,N9993,N9994,N9995,N9996,N9998,N9999,N10000 
	,N10001,N10003,N10004,N10005,N10006,N10007,N10008,N10009 
	,N10010,N10011,N10012,N10013,N10015,N10016,N10017,N10018 
	,N10020,N10021,N10023,N10024,N10025,N10026,N10027,N10028 
	,N10029,N10030,N10031,N10032,N10033,N10034,N10035,N10036 
	,N10037,N10038,N10039,N10040,N10041,N10042,N10044,N10045 
	,N10046,N10047,N10048,N10049,N10050,N10051,N10052,N10053 
	,N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061 
	,N10062,N10064,N10065,N10066,N10067,N10068,N10069,N10070 
	,N10071,N10072,N10073,N10074,N10075,N10076,N10078,N10079 
	,N10080,N10081,N10082,N10085,N10086,N10087,N10088,N10089 
	,N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097 
	,N10098,N10099,N10100,N10101,N10102,N10103,N10104,N10105 
	,N10106,N10108,N10109,N10110,N10111,N10112,N10114,N10115 
	,N10116,N10117,N10118,N10119,N10120,N10121,N10122,N10123 
	,N10124,N10125,N10126,N10127,N10128,N10129,N10130,N10131 
	,N10132,N10133,N10134,N10135,N10137,N10138,N10139,N10142 
	,N10143,N10144,N10145,N10146,N10147,N10148,N10149,N10150 
	,N10151,N10152,N10153,N10154,N10155,N10156,N10157,N10158 
	,N10159,N10160,N10161,N10163,N10164,N10165,N10167,N10169 
	,N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177 
	,N10178,N10179,N10181,N10182,N10183,N10184,N10185,N10186 
	,N10187,N10188,N10189,N10190,N10191,N10192,N10193,N10194 
	,N10195,N10196,N10197,N10199,N10200,N10201,N10202,N10203 
	,N10205,N10206,N10207,N10208,N10209,N10211,N10212,N10213 
	,N10214,N10215,N10216,N10217,N10218,N10219,N10220,N10221 
	,N10222,N10223,N10224,N10226,N10227,N10228,N10229,N10231 
	,N10232,N10234,N10235,N10236,N10237,N10238,N10239,N10240 
	,N10241,N10242,N10243,N10244,N10245,N10246,N10247,N10248 
	,N10249,N10250,N10251,N10252,N10253,N10255,N10256,N10257 
	,N10258,N10259,N10261,N10262,N10263,N10264,N10265,N10266 
	,N10267,N10268,N10269,N10271,N10272,N10273,N10274,N10275 
	,N10276,N10277,N10278,N10279,N10280,N10281,N10282,N10284 
	,N10285,N10286,N10287,N10288,N10290,N10292,N10293,N10294 
	,N10295,N10296,N10297,N10298,N10299,N10300,N10301,N10302 
	,N10303,N10304,N10305,N10306,N10307,N10308,N10310,N11898 
	,N11899,N11901,N11902,N11906,N11907,N11909,N11910,N11911 
	,N11912,N11914,N11915,N11918,N11919,N11920,N11921,N11923 
	,N11925,N11927,N11928,N11929,N11931,N11933,N11935,N11936 
	,N11937,N11941,N11942,N11943,N11944,N11945,N11946,N11948 
	,N11950,N11951,N11953,N11956,N11958,N11959,N11961,N11965 
	,N11966,N11968,N11969,N11970,N11972,N11973,N11975,N11976 
	,N11977,N11981,N11983,N11984,N11985,N11988,N11989,N11990 
	,N11991,N11992,N11993,N11995,N11996,N11998,N11999,N12000 
	,N12002,N12005,N12007,N12008,N12009,N12011,N12013,N12014 
	,N12015,N12017,N12020,N12021,N12022,N12023,N12024,N12027 
	,N12028,N12030,N12031,N12033,N12035,N12036,N12037,N12040 
	,N12042,N12043,N12044,N12045,N12047,N12048,N12051,N12052 
	,N12054,N12055,N12057,N12059,N12060,N12061,N12062,N12063 
	,N12065,N12066,N12068,N12069,N12072,N12073,N12075,N12076 
	,N12077,N12080,N12082,N12083,N12084,N12086,N12087,N12090 
	,N12094,N12095,N12097,N12099,N12100,N12101,N12102,N12103 
	,N12104,N12107,N12108,N12110,N12112,N12113,N12115,N12116 
	,N12117,N12120,N12121,N12123,N12124,N12125,N12126,N12127 
	,N12128,N12131,N12132,N12133,N12135,N12137,N12138,N12140 
	,N12143,N12146,N12148,N12149,N12150,N12151,N12154,N12155 
	,N12156,N12157,N12158,N12160,N12161,N12163,N12164,N12168 
	,N12169,N12171,N12172,N12174,N12177,N12178,N12179,N12180 
	,N12181,N12182,N12184,N12185,N12187,N12188,N12189,N12192 
	,N12194,N12196,N12197,N12198,N12201,N12202,N12203,N12204 
	,N12206,N12207,N12209,N12210,N12211,N12212,N12213,N12214 
	,N12217,N12218,N12220,N12222,N12225,N12226,N12227,N12229 
	,N12230,N12232,N12234,N12235,N12236,N12239,N12240,N12242 
	,N12243,N12245,N12246,N12249,N12250,N12251,N12252,N12254 
	,N12255,N12257,N12258,N12259,N12260,N12261,N12263,N12264 
	,N12265,N12266,N12269,N12270,N12272,N12273,N12276,N12278 
	,N12279,N12281,N12282,N12283,N12284,N12285,N12286,N12288 
	,N12290,N12291,N12294,N12295,N12297,N12298,N12299,N12300 
	,N12302,N12305,N12307,N12308,N12310,N12311,N12313,N12317 
	,N12318,N12320,N12321,N12322,N12323,N12324,N12328,N12329 
	,N12330,N12331,N12333,N12335,N12336,N12337,N12341,N12344 
	,N12345,N12346,N12347,N12348,N12349,N12350,N12353,N12354 
	,N12355,N12356,N12357,N12360,N12362,N12364,N12365,N12367 
	,N12371,N12373,N12374,N12375,N12376,N12380,N12381,N12382 
	,N12383,N12384,N12385,N12387,N12390,N12391,N12392,N12394 
	,N12397,N12399,N12400,N12401,N12404,N12405,N12406,N12407 
	,N12408,N12410,N12411,N12414,N12415,N12416,N12418,N12421 
	,N12423,N12424,N12426,N12427,N12429,N12431,N12432,N12434 
	,N12435,N12436,N12437,N12440,N12441,N12443,N12444,N12446 
	,N12448,N12449,N12450,N12451,N12453,N12456,N12457,N12458 
	,N12459,N12460,N12463,N12464,N12466,N12467,N12469,N12470 
	,N12472,N12473,N12475,N12476,N12478,N12479,N12481,N12484 
	,N12485,N12487,N12491,N12492,N12494,N12495,N12497,N12498 
	,N12501,N12503,N12504,N12506,N12508,N12509,N12512,N12513 
	,N12515,N12516,N12517,N12518,N12519,N12522,N12524,N13041 
	,N13185,N13187,N13208,N13216,N13219,N13221,N13225,N13227 
	,N13230,N13236,N13240,N13288,N13292,N13316,N13332,N13334 
	,N13337,N13339,N13340,N13341,N13343,N13346,N13347,N13348 
	,N13349,N13351,N13352,N13354,N13355,N13356,N13358,N13359 
	,N13360,N13362,N13365,N13367,N13368,N13370,N13371,N13373 
	,N13374,N13375,N13376,N13377,N13379,N13380,N13383,N13384 
	,N13386,N13387,N13388,N13391,N13392,N13393,N13394,N13395 
	,N13397,N13398,N13399,N13402,N13404,N13405,N13406,N13407 
	,N13409,N13411,N13470,N13472,N13475,N13490,N13491,N13492 
	,N13495,N13496,N13497,N13498,N13501,N13502,N13503,N13506 
	,N13507,N13509,N13510,N13511,N13512,N13513,N13516,N13517 
	,N13518,N13521,N13522,N13525,N13526,N13527,N13528,N13531 
	,N13532,N13533,N13534,N13535,N13539,N13540,N13541,N13542 
	,N13545,N13546,N13547,N13548,N13549,N13551,N13553,N13554 
	,N13555,N13556,N13558,N13560,N13562,N13563,N13564,N13565 
	,N13566,N13569,N13570,N13571,N13574,N13575,N13576,N13577 
	,N13578,N13581,N13582,N13583,N13584,N13587,N13588,N13589 
	,N13591,N13594,N13595,N13596,N13597,N13598,N13601,N13602 
	,N13603,N13604,N13605,N13608,N13609,N13610,N13611,N13612 
	,N13615,N13616,N13617,N13618,N13621,N13622,N13623,N13627 
	,N13628,N13629,N13630,N13633,N13634,N13635,N13638,N13639 
	,N13640,N13786,N13800,N13809,N13818,N13822,N13832,N13845 
	,N13863,N13877,N13925,N13934,N13937,N13939,N13940,N13943 
	,N13947,N13955,N13957,N13969,N13970,N14019,N14026,N19007 
	,N19009,N19011,N19018,N19025,N19032,N19047,N19054,N37704 
	,N37712,N37720;
INVXL inst_blk01_cellmath__39_I170 (.Y(N3949), .A(a_man[0]));
INVXL inst_blk01_cellmath__39_I171 (.Y(N4417), .A(a_man[1]));
INVXL inst_blk01_cellmath__39_I172 (.Y(N4381), .A(a_man[2]));
INVXL inst_blk01_cellmath__39_I173 (.Y(N4428), .A(a_man[3]));
INVXL inst_blk01_cellmath__39_I174 (.Y(N4287), .A(a_man[4]));
INVXL inst_blk01_cellmath__39_I175 (.Y(N4614), .A(a_man[5]));
INVXL inst_blk01_cellmath__39_I176 (.Y(N4080), .A(a_man[6]));
INVXL inst_blk01_cellmath__39_I177 (.Y(N4508), .A(a_man[7]));
INVXL inst_blk01_cellmath__39_I178 (.Y(N4104), .A(a_man[8]));
INVXL inst_blk01_cellmath__39_I179 (.Y(N4415), .A(a_man[9]));
INVXL inst_blk01_cellmath__39_I180 (.Y(N4015), .A(a_man[10]));
INVXL inst_blk01_cellmath__39_I181 (.Y(N4322), .A(a_man[11]));
INVXL inst_blk01_cellmath__39_I182 (.Y(N3922), .A(a_man[12]));
INVXL inst_blk01_cellmath__39_I183 (.Y(N4236), .A(a_man[13]));
INVXL inst_blk01_cellmath__39_I184 (.Y(N4548), .A(a_man[14]));
INVXL inst_blk01_cellmath__39_I185 (.Y(N4145), .A(a_man[15]));
INVXL inst_blk01_cellmath__39_I186 (.Y(N4454), .A(a_man[16]));
INVXL inst_blk01_cellmath__39_I187 (.Y(N4052), .A(a_man[17]));
INVXL inst_blk01_cellmath__39_I188 (.Y(N4368), .A(a_man[18]));
INVXL inst_blk01_cellmath__39_I189 (.Y(N3958), .A(a_man[19]));
INVXL inst_blk01_cellmath__39_I190 (.Y(N4274), .A(a_man[20]));
INVXL inst_blk01_cellmath__39_I191 (.Y(N4595), .A(a_man[21]));
INVXL inst_blk01_cellmath__39_I192 (.Y(N4181), .A(a_man[22]));
INVXL inst_blk01_cellmath__39_I193 (.Y(N4273), .A(N4428));
ADDHX1 inst_blk01_cellmath__39_I194 (.CO(N4335), .S(N4182), .A(N4287), .B(N4428));
ADDHX1 inst_blk01_cellmath__39_I195 (.CO(N3933), .S(N4496), .A(N4614), .B(N4381));
ADDFX1 inst_blk01_cellmath__39_I196 (.CO(N4157), .S(N4004), .A(N3949), .B(N4428), .CI(a_man[6]));
ADDHX1 inst_blk01_cellmath__39_I197 (.CO(N4467), .S(N4308), .A(N4508), .B(N4080));
ADDFX1 inst_blk01_cellmath__39_I198 (.CO(N4063), .S(N4635), .A(N4417), .B(N4287), .CI(N4308));
ADDHX1 inst_blk01_cellmath__39_I199 (.CO(N4379), .S(N4217), .A(N4104), .B(N4614));
ADDFX1 inst_blk01_cellmath__39_I200 (.CO(N3968), .S(N4531), .A(N4467), .B(N4381), .CI(N4217));
ADDFX1 inst_blk01_cellmath__39_I201 (.CO(N4439), .S(N4350), .A(N4080), .B(a_man[0]), .CI(N4415));
ADDFX1 inst_blk01_cellmath__39_I202 (.CO(N4284), .S(N4131), .A(N4428), .B(N4379), .CI(N4350));
ADDFX1 inst_blk01_cellmath__39_I203 (.CO(N4191), .S(N4233), .A(N4015), .B(a_man[1]), .CI(N4508));
ADDFX1 inst_blk01_cellmath__39_I204 (.CO(N4038), .S(N4611), .A(N4287), .B(N4439), .CI(N4233));
ADDFX1 inst_blk01_cellmath__39_I205 (.CO(N3945), .S(N4119), .A(N4104), .B(a_man[2]), .CI(N4322));
ADDFX1 inst_blk01_cellmath__39_I206 (.CO(N4505), .S(N4349), .A(N4614), .B(N4191), .CI(N4119));
ADDFX1 inst_blk01_cellmath__39_I207 (.CO(N4412), .S(N3998), .A(N3922), .B(a_man[3]), .CI(N4415));
ADDFX1 inst_blk01_cellmath__39_I208 (.CO(N4257), .S(N4100), .A(N3945), .B(N4080), .CI(N3998));
ADDFX1 inst_blk01_cellmath__39_I209 (.CO(N4167), .S(N4609), .A(N4236), .B(a_man[4]), .CI(N4015));
ADDFX1 inst_blk01_cellmath__39_I210 (.CO(N4013), .S(N4573), .A(N4508), .B(N4412), .CI(N4609));
XNOR2X1 inst_blk01_cellmath__39_I211 (.Y(N4320), .A(a_man[5]), .B(N3949));
OR2XL inst_blk01_cellmath__39_I212 (.Y(N4481), .A(a_man[5]), .B(N3949));
ADDFX1 inst_blk01_cellmath__39_I213 (.CO(N4543), .S(N3978), .A(N4322), .B(N4548), .CI(N4104));
ADDFX1 inst_blk01_cellmath__39_I214 (.CO(N4389), .S(N4231), .A(N4167), .B(N4320), .CI(N3978));
ADDFX1 inst_blk01_cellmath__39_I215 (.CO(N4143), .S(N3982), .A(N4417), .B(a_man[6]), .CI(N4145));
ADDFX1 inst_blk01_cellmath__39_I216 (.CO(N4622), .S(N4587), .A(N4415), .B(N3922), .CI(N4481));
ADDFX1 inst_blk01_cellmath__39_I217 (.CO(N4450), .S(N4296), .A(N4543), .B(N3982), .CI(N4587));
ADDHX1 inst_blk01_cellmath__39_I218 (.CO(N4202), .S(N4049), .A(a_man[7]), .B(N4381));
ADDFX1 inst_blk01_cellmath__39_I219 (.CO(N4519), .S(N4365), .A(N4454), .B(a_man[0]), .CI(N4236));
ADDFX1 inst_blk01_cellmath__39_I220 (.CO(N4270), .S(N4461), .A(N4049), .B(N4015), .CI(N4143));
ADDFX1 inst_blk01_cellmath__39_I221 (.CO(N4117), .S(N3955), .A(N4365), .B(N4622), .CI(N4461));
ADDFX1 inst_blk01_cellmath__39_I222 (.CO(N4024), .S(N4343), .A(N4428), .B(a_man[8]), .CI(N4052));
ADDFX1 inst_blk01_cellmath__39_I223 (.CO(N4591), .S(N4425), .A(N4202), .B(N4519), .CI(N4343));
ADDFX1 inst_blk01_cellmath__39_I224 (.CO(N4490), .S(N4225), .A(N4322), .B(a_man[1]), .CI(N4548));
ADDFX1 inst_blk01_cellmath__39_I225 (.CO(N4333), .S(N4177), .A(N4425), .B(N4270), .CI(N4225));
XNOR2X1 inst_blk01_cellmath__39_I226 (.Y(N3931), .A(a_man[9]), .B(N4287));
OR2XL inst_blk01_cellmath__39_I227 (.Y(N4087), .A(a_man[9]), .B(N4287));
ADDFX1 inst_blk01_cellmath__39_I228 (.CO(N4155), .S(N4326), .A(N4368), .B(a_man[2]), .CI(N4145));
ADDFX1 inst_blk01_cellmath__39_I229 (.CO(N3997), .S(N4556), .A(N4490), .B(N4024), .CI(N4326));
ADDFX1 inst_blk01_cellmath__39_I230 (.CO(N4632), .S(N4208), .A(N3949), .B(N3922), .CI(N3931));
ADDFX1 inst_blk01_cellmath__39_I231 (.CO(N4463), .S(N4305), .A(N4556), .B(N4591), .CI(N4208));
ADDFX1 inst_blk01_cellmath__39_I232 (.CO(N4213), .S(N4059), .A(N4614), .B(a_man[10]), .CI(N3958));
ADDFX1 inst_blk01_cellmath__39_I233 (.CO(N3967), .S(N4092), .A(N4454), .B(a_man[3]), .CI(N4236));
ADDFX1 inst_blk01_cellmath__39_I234 (.CO(N4529), .S(N4376), .A(N4155), .B(N4059), .CI(N4092));
ADDFX1 inst_blk01_cellmath__39_I235 (.CO(N4436), .S(N3971), .A(N4087), .B(N4417), .CI(N4632));
ADDFX1 inst_blk01_cellmath__39_I236 (.CO(N4281), .S(N4128), .A(N3997), .B(N4376), .CI(N3971));
ADDFX1 inst_blk01_cellmath__39_I237 (.CO(N4035), .S(N4607), .A(N4080), .B(a_man[11]), .CI(N4274));
ADDFX1 inst_blk01_cellmath__39_I238 (.CO(N4502), .S(N4575), .A(N4052), .B(a_man[4]), .CI(N4548));
ADDFX1 inst_blk01_cellmath__39_I239 (.CO(N4347), .S(N4189), .A(N3967), .B(N4607), .CI(N4575));
ADDFX1 inst_blk01_cellmath__39_I240 (.CO(N4254), .S(N4455), .A(N4213), .B(N4381), .CI(N4529));
ADDFX1 inst_blk01_cellmath__39_I241 (.CO(N4097), .S(N3941), .A(N4436), .B(N4189), .CI(N4455));
ADDFX1 inst_blk01_cellmath__39_I242 (.CO(N4569), .S(N4410), .A(N4508), .B(a_man[12]), .CI(N4595));
ADDFX1 inst_blk01_cellmath__39_I243 (.CO(N4318), .S(N4336), .A(N4145), .B(a_man[5]), .CI(N4368));
ADDFX1 inst_blk01_cellmath__39_I244 (.CO(N4165), .S(N4010), .A(N4502), .B(N4410), .CI(N4336));
ADDFX1 inst_blk01_cellmath__39_I245 (.CO(N4073), .S(N4218), .A(N4035), .B(N4428), .CI(N4347));
ADDFX1 inst_blk01_cellmath__39_I246 (.CO(N4641), .S(N4477), .A(N4010), .B(N4254), .CI(N4218));
ADDFX1 inst_blk01_cellmath__39_I247 (.CO(N4386), .S(N4227), .A(N4104), .B(a_man[13]), .CI(N4181));
ADDFX1 inst_blk01_cellmath__39_I248 (.CO(N4139), .S(N4099), .A(N3958), .B(a_man[6]), .CI(N4454));
ADDFX1 inst_blk01_cellmath__39_I249 (.CO(N3976), .S(N4539), .A(N4318), .B(N4099), .CI(N4227));
ADDFX1 inst_blk01_cellmath__39_I250 (.CO(N4619), .S(N3983), .A(N4569), .B(N4287), .CI(N4165));
ADDFX1 inst_blk01_cellmath__39_I251 (.CO(N4446), .S(N4292), .A(N4539), .B(N4073), .CI(N3983));
ADDFX1 inst_blk01_cellmath__39_I252 (.CO(N4197), .S(N4047), .A(N4274), .B(N4548), .CI(N4415));
ADDFX1 inst_blk01_cellmath__39_I253 (.CO(N4267), .S(N4557), .A(N4052), .B(a_man[7]), .CI(N4614));
ADDFX1 inst_blk01_cellmath__39_I254 (.CO(N4112), .S(N3952), .A(N4386), .B(N4139), .CI(N4557));
ADDFX1 inst_blk01_cellmath__39_I255 (.CO(N4020), .S(N4437), .A(N4047), .B(N3949), .CI(N3976));
ADDFX1 inst_blk01_cellmath__39_I256 (.CO(N4586), .S(N4421), .A(N4619), .B(N3952), .CI(N4437));
XNOR2X1 inst_blk01_cellmath__39_I257 (.Y(N4316), .A(a_man[15]), .B(N4015));
OR2XL inst_blk01_cellmath__39_I258 (.Y(N4488), .A(a_man[15]), .B(N4015));
ADDFX1 inst_blk01_cellmath__39_I259 (.CO(N4329), .S(N4174), .A(N4267), .B(N4197), .CI(N4316));
ADDFX1 inst_blk01_cellmath__39_I260 (.CO(N4241), .S(N4198), .A(N4595), .B(a_man[8]), .CI(N4368));
ADDFX1 inst_blk01_cellmath__39_I261 (.CO(N4083), .S(N3927), .A(N4417), .B(N4080), .CI(N4198));
ADDFX1 inst_blk01_cellmath__39_I262 (.CO(N3992), .S(N4084), .A(N4112), .B(a_man[14]), .CI(N4174));
ADDFX1 inst_blk01_cellmath__39_I263 (.CO(N4552), .S(N4397), .A(N3927), .B(N4020), .CI(N4084));
ADDFX1 inst_blk01_cellmath__39_I264 (.CO(N4303), .S(N4149), .A(N4181), .B(N4322), .CI(N4454));
ADDFX1 inst_blk01_cellmath__39_I265 (.CO(N4210), .S(N4056), .A(N3958), .B(a_man[9]), .CI(N4508));
ADDFX1 inst_blk01_cellmath__39_I266 (.CO(N3963), .S(N3936), .A(N4381), .B(a_man[0]), .CI(N4488));
ADDFX1 inst_blk01_cellmath__39_I267 (.CO(N4526), .S(N4371), .A(N4056), .B(N4149), .CI(N3936));
ADDFX1 inst_blk01_cellmath__39_I268 (.CO(N4432), .S(N4533), .A(N4329), .B(N4241), .CI(N4083));
ADDFX1 inst_blk01_cellmath__39_I269 (.CO(N4278), .S(N4124), .A(N4371), .B(N3992), .CI(N4533));
ADDFX1 inst_blk01_cellmath__39_I270 (.CO(N4032), .S(N4601), .A(N4274), .B(N3922), .CI(N4052));
ADDFX1 inst_blk01_cellmath__39_I271 (.CO(N3938), .S(N4499), .A(N4104), .B(a_man[10]), .CI(N4428));
ADDFX1 inst_blk01_cellmath__39_I272 (.CO(N4406), .S(N4393), .A(a_man[16]), .B(a_man[1]), .CI(N4210));
ADDFX1 inst_blk01_cellmath__39_I273 (.CO(N4251), .S(N4093), .A(N4601), .B(N3963), .CI(N4393));
ADDFX1 inst_blk01_cellmath__39_I274 (.CO(N4162), .S(N4276), .A(N4499), .B(N4303), .CI(N4526));
ADDFX1 inst_blk01_cellmath__39_I275 (.CO(N4007), .S(N4567), .A(N4432), .B(N4093), .CI(N4276));
ADDFX1 inst_blk01_cellmath__39_I276 (.CO(N4638), .S(N4158), .A(N4236), .B(a_man[18]), .CI(N4595));
ADDFX1 inst_blk01_cellmath__39_I277 (.CO(N4472), .S(N4314), .A(N3938), .B(N4032), .CI(N4158));
ADDFX1 inst_blk01_cellmath__39_I278 (.CO(N4383), .S(N4039), .A(N4287), .B(a_man[11]), .CI(N4415));
ADDFX1 inst_blk01_cellmath__39_I279 (.CO(N4221), .S(N4069), .A(a_man[17]), .B(a_man[2]), .CI(N4039));
ADDFX1 inst_blk01_cellmath__39_I280 (.CO(N4134), .S(N3920), .A(N4314), .B(N4406), .CI(N4069));
ADDFX1 inst_blk01_cellmath__39_I281 (.CO(N3972), .S(N4535), .A(N4251), .B(N4162), .CI(N3920));
ADDFX1 inst_blk01_cellmath__39_I282 (.CO(N4441), .S(N4289), .A(N4181), .B(N4548), .CI(N3958));
ADDFX1 inst_blk01_cellmath__39_I283 (.CO(N4355), .S(N4194), .A(N4015), .B(a_man[12]), .CI(N4614));
ADDFX1 inst_blk01_cellmath__39_I284 (.CO(N4107), .S(N4494), .A(a_man[0]), .B(a_man[3]), .CI(N4638));
ADDFX1 inst_blk01_cellmath__39_I285 (.CO(N3948), .S(N4510), .A(N4194), .B(N4289), .CI(N4494));
ADDFX1 inst_blk01_cellmath__39_I286 (.CO(N4580), .S(N4377), .A(N4472), .B(N4383), .CI(N4221));
ADDFX1 inst_blk01_cellmath__39_I287 (.CO(N4416), .S(N4263), .A(N4134), .B(N4510), .CI(N4377));
ADDFX1 inst_blk01_cellmath__39_I288 (.CO(N4170), .S(N4016), .A(N4322), .B(N4145), .CI(N4274));
ADDFX1 inst_blk01_cellmath__39_I289 (.CO(N4079), .S(N3923), .A(a_man[4]), .B(a_man[13]), .CI(N4080));
ADDFX1 inst_blk01_cellmath__39_I290 (.CO(N4549), .S(N4230), .A(a_man[19]), .B(a_man[1]), .CI(N4355));
ADDFX1 inst_blk01_cellmath__39_I291 (.CO(N4392), .S(N4238), .A(N4016), .B(N4107), .CI(N4230));
ADDFX1 inst_blk01_cellmath__39_I292 (.CO(N4300), .S(N4115), .A(N3923), .B(N4441), .CI(N3948));
ADDFX1 inst_blk01_cellmath__39_I293 (.CO(N4146), .S(N3988), .A(N4580), .B(N4238), .CI(N4115));
ADDHX1 inst_blk01_cellmath__39_I294 (.CO(N4624), .S(N4456), .A(a_man[21]), .B(N4454));
ADDFX1 inst_blk01_cellmath__39_I295 (.CO(N4369), .S(N3995), .A(N3922), .B(a_man[14]), .CI(N4508));
ADDFX1 inst_blk01_cellmath__39_I296 (.CO(N4207), .S(N4053), .A(N4079), .B(N4170), .CI(N3995));
ADDFX1 inst_blk01_cellmath__39_I297 (.CO(N4121), .S(N4604), .A(a_man[2]), .B(a_man[5]), .CI(a_man[0]));
ADDFX1 inst_blk01_cellmath__39_I298 (.CO(N3960), .S(N4524), .A(a_man[20]), .B(N4456), .CI(N4604));
ADDFX1 inst_blk01_cellmath__39_I299 (.CO(N4597), .S(N4476), .A(N4524), .B(N4549), .CI(N4053));
ADDFX1 inst_blk01_cellmath__39_I300 (.CO(N4430), .S(N4275), .A(N4392), .B(N4300), .CI(N4476));
XNOR2X1 inst_blk01_cellmath__39_I301 (.Y(N4029), .A(N4052), .B(N4236));
OR2XL inst_blk01_cellmath__39_I302 (.Y(N4183), .A(N4052), .B(N4236));
ADDFX1 inst_blk01_cellmath__39_I303 (.CO(N4249), .S(N4584), .A(a_man[15]), .B(a_man[22]), .CI(N4104));
ADDFX1 inst_blk01_cellmath__39_I304 (.CO(N4090), .S(N3935), .A(N4369), .B(N4029), .CI(N4584));
ADDFX1 inst_blk01_cellmath__39_I305 (.CO(N4006), .S(N4457), .A(a_man[3]), .B(a_man[6]), .CI(a_man[1]));
ADDFX1 inst_blk01_cellmath__39_I306 (.CO(N4564), .S(N4404), .A(N4624), .B(N4121), .CI(N4457));
ADDFX1 inst_blk01_cellmath__39_I307 (.CO(N4469), .S(N4338), .A(N4207), .B(N3960), .CI(N4404));
ADDFX1 inst_blk01_cellmath__39_I308 (.CO(N4309), .S(N4160), .A(N3935), .B(N4597), .CI(N4338));
ADDFX1 inst_blk01_cellmath__39_I309 (.CO(N4219), .S(N4220), .A(N4368), .B(a_man[16]), .CI(N4548));
ADDFX1 inst_blk01_cellmath__39_I310 (.CO(N4065), .S(N4636), .A(N4006), .B(N4249), .CI(N4220));
ADDFX1 inst_blk01_cellmath__39_I311 (.CO(N3970), .S(N4106), .A(N4415), .B(a_man[7]), .CI(a_man[4]));
ADDFX1 inst_blk01_cellmath__39_I312 (.CO(N4532), .S(N4380), .A(a_man[2]), .B(N4183), .CI(N4106));
ADDFX1 inst_blk01_cellmath__39_I313 (.CO(N4440), .S(N3987), .A(N4090), .B(N4564), .CI(N4636));
ADDFX1 inst_blk01_cellmath__39_I314 (.CO(N4285), .S(N4132), .A(N4380), .B(N4469), .CI(N3987));
ADDHX1 inst_blk01_cellmath__39_I315 (.CO(N4041), .S(N4613), .A(a_man[17]), .B(N3958));
ADDFX1 inst_blk01_cellmath__39_I316 (.CO(N4352), .S(N4193), .A(N4145), .B(a_man[8]), .CI(N4015));
ADDFX1 inst_blk01_cellmath__39_I317 (.CO(N4103), .S(N4596), .A(a_man[3]), .B(a_man[5]), .CI(N4613));
ADDFX1 inst_blk01_cellmath__39_I318 (.CO(N3946), .S(N4507), .A(N4219), .B(N4193), .CI(N4596));
ADDFX1 inst_blk01_cellmath__39_I319 (.CO(N4574), .S(N4468), .A(N4065), .B(N3970), .CI(N4532));
ADDFX1 inst_blk01_cellmath__39_I320 (.CO(N4413), .S(N4259), .A(N4440), .B(N4507), .CI(N4468));
ADDHX1 inst_blk01_cellmath__39_I321 (.CO(N4169), .S(N4014), .A(a_man[18]), .B(N4274));
ADDFX1 inst_blk01_cellmath__39_I322 (.CO(N4483), .S(N4321), .A(N4454), .B(a_man[9]), .CI(N4322));
ADDFX1 inst_blk01_cellmath__39_I323 (.CO(N4235), .S(N4351), .A(a_man[4]), .B(a_man[6]), .CI(N4041));
ADDFX1 inst_blk01_cellmath__39_I324 (.CO(N4076), .S(N3919), .A(N4321), .B(N4103), .CI(N4351));
ADDFX1 inst_blk01_cellmath__39_I325 (.CO(N3985), .S(N4232), .A(N4352), .B(N4014), .CI(N3946));
ADDFX1 inst_blk01_cellmath__39_I326 (.CO(N4545), .S(N4390), .A(N3919), .B(N4574), .CI(N4232));
ADDHX1 inst_blk01_cellmath__39_I327 (.CO(N4297), .S(N4144), .A(a_man[19]), .B(N4595));
ADDFX1 inst_blk01_cellmath__39_I328 (.CO(N4623), .S(N4453), .A(N4052), .B(a_man[10]), .CI(N3922));
ADDFX1 inst_blk01_cellmath__39_I329 (.CO(N4366), .S(N4118), .A(a_man[5]), .B(a_man[7]), .CI(N4169));
ADDFX1 inst_blk01_cellmath__39_I330 (.CO(N4204), .S(N4050), .A(N4453), .B(N4235), .CI(N4118));
ADDFX1 inst_blk01_cellmath__39_I331 (.CO(N4120), .S(N3999), .A(N4483), .B(N4144), .CI(N4076));
ADDFX1 inst_blk01_cellmath__39_I332 (.CO(N3957), .S(N4521), .A(N4050), .B(N3985), .CI(N3999));
ADDHX1 inst_blk01_cellmath__39_I333 (.CO(N4427), .S(N4271), .A(a_man[20]), .B(N4181));
ADDFX1 inst_blk01_cellmath__39_I334 (.CO(N4026), .S(N4592), .A(N4368), .B(a_man[11]), .CI(N4236));
ADDFX1 inst_blk01_cellmath__39_I335 (.CO(N4493), .S(N4608), .A(a_man[6]), .B(a_man[8]), .CI(N4297));
ADDFX1 inst_blk01_cellmath__39_I336 (.CO(N4334), .S(N4180), .A(N4592), .B(N4366), .CI(N4608));
ADDFX1 inst_blk01_cellmath__39_I337 (.CO(N4247), .S(N4478), .A(N4623), .B(N4271), .CI(N4204));
ADDFX1 inst_blk01_cellmath__39_I338 (.CO(N4088), .S(N3932), .A(N4180), .B(N4120), .CI(N4478));
ADDFX1 inst_blk01_cellmath__39_I339 (.CO(N4560), .S(N4403), .A(N3958), .B(a_man[21]), .CI(N4548));
ADDFX1 inst_blk01_cellmath__39_I340 (.CO(N4307), .S(N4360), .A(a_man[9]), .B(a_man[12]), .CI(a_man[7]));
ADDFX1 inst_blk01_cellmath__39_I341 (.CO(N4156), .S(N4001), .A(N4403), .B(N4493), .CI(N4360));
ADDFX1 inst_blk01_cellmath__39_I342 (.CO(N4061), .S(N4243), .A(N4026), .B(N4427), .CI(N4334));
ADDFX1 inst_blk01_cellmath__39_I343 (.CO(N4634), .S(N4465), .A(N4001), .B(N4247), .CI(N4243));
XNOR2X1 inst_blk01_cellmath__39_I344 (.Y(N4215), .A(N4274), .B(N4145));
OR2XL inst_blk01_cellmath__39_I345 (.Y(N4378), .A(N4274), .B(N4145));
ADDFX1 inst_blk01_cellmath__39_I346 (.CO(N4438), .S(N4342), .A(a_man[13]), .B(a_man[22]), .CI(a_man[10]));
ADDFX1 inst_blk01_cellmath__39_I347 (.CO(N4283), .S(N4130), .A(N4560), .B(N4215), .CI(N4342));
ADDFX1 inst_blk01_cellmath__39_I348 (.CO(N4190), .S(N4224), .A(N4307), .B(a_man[8]), .CI(N4156));
ADDFX1 inst_blk01_cellmath__39_I349 (.CO(N4036), .S(N4610), .A(N4130), .B(N4061), .CI(N4224));
ADDFX1 inst_blk01_cellmath__39_I350 (.CO(N3943), .S(N4109), .A(N4595), .B(a_man[14]), .CI(N4454));
ADDFX1 inst_blk01_cellmath__39_I351 (.CO(N4504), .S(N4348), .A(N4378), .B(N4438), .CI(N4109));
ADDFX1 inst_blk01_cellmath__39_I352 (.CO(N4411), .S(N3989), .A(a_man[9]), .B(a_man[11]), .CI(N4283));
ADDFX1 inst_blk01_cellmath__39_I353 (.CO(N4256), .S(N4098), .A(N4348), .B(N4190), .CI(N3989));
ADDHX1 inst_blk01_cellmath__39_I354 (.CO(N4012), .S(N4571), .A(a_man[15]), .B(N4181));
ADDFX1 inst_blk01_cellmath__39_I355 (.CO(N4319), .S(N4166), .A(a_man[10]), .B(a_man[12]), .CI(N4052));
ADDFX1 inst_blk01_cellmath__39_I356 (.CO(N4075), .S(N4600), .A(N3943), .B(N4571), .CI(N4166));
ADDFX1 inst_blk01_cellmath__39_I357 (.CO(N3917), .S(N4479), .A(N4411), .B(N4504), .CI(N4600));
ADDFX1 inst_blk01_cellmath__39_I358 (.CO(N4387), .S(N4229), .A(N4368), .B(a_man[16]), .CI(a_man[13]));
ADDFX1 inst_blk01_cellmath__39_I359 (.CO(N4141), .S(N4471), .A(N4319), .B(a_man[11]), .CI(N4012));
ADDFX1 inst_blk01_cellmath__39_I360 (.CO(N3979), .S(N4540), .A(N4229), .B(N4075), .CI(N4471));
XNOR2X1 inst_blk01_cellmath__39_I361 (.Y(N4294), .A(N3958), .B(a_man[17]));
OR2XL inst_blk01_cellmath__39_I362 (.Y(N4449), .A(N3958), .B(a_man[17]));
ADDFX1 inst_blk01_cellmath__39_I363 (.CO(N4516), .S(N4577), .A(a_man[12]), .B(a_man[14]), .CI(N4387));
ADDFX1 inst_blk01_cellmath__39_I364 (.CO(N4361), .S(N4201), .A(N4294), .B(N4141), .CI(N4577));
XNOR2X1 inst_blk01_cellmath__39_I365 (.Y(N3953), .A(N4274), .B(a_man[18]));
OR2XL inst_blk01_cellmath__39_I366 (.Y(N4113), .A(N4274), .B(a_man[18]));
ADDFX1 inst_blk01_cellmath__39_I367 (.CO(N4176), .S(N3959), .A(a_man[13]), .B(a_man[15]), .CI(N4449));
ADDFX1 inst_blk01_cellmath__39_I368 (.CO(N4022), .S(N4588), .A(N3953), .B(N4516), .CI(N3959));
XNOR2X1 inst_blk01_cellmath__39_I369 (.Y(N4331), .A(N4595), .B(a_man[19]));
OR2XL inst_blk01_cellmath__39_I370 (.Y(N4489), .A(N4595), .B(a_man[19]));
ADDFX1 inst_blk01_cellmath__39_I371 (.CO(N4554), .S(N4064), .A(a_man[14]), .B(a_man[16]), .CI(N4113));
ADDFX1 inst_blk01_cellmath__39_I372 (.CO(N4400), .S(N4245), .A(N4331), .B(N4176), .CI(N4064));
XNOR2X1 inst_blk01_cellmath__39_I373 (.Y(N3994), .A(N4181), .B(a_man[20]));
OR2XL inst_blk01_cellmath__39_I374 (.Y(N4153), .A(N4181), .B(a_man[20]));
ADDFX1 inst_blk01_cellmath__39_I375 (.CO(N4212), .S(N4168), .A(a_man[15]), .B(a_man[17]), .CI(N4489));
ADDFX1 inst_blk01_cellmath__39_I376 (.CO(N4058), .S(N4630), .A(N3994), .B(N4554), .CI(N4168));
ADDFX1 inst_blk01_cellmath__39_I377 (.CO(N4528), .S(N4374), .A(a_man[16]), .B(a_man[18]), .CI(N4595));
ADDFX1 inst_blk01_cellmath__39_I378 (.CO(N4434), .S(N4280), .A(N4212), .B(N4153), .CI(N4374));
ADDFX1 inst_blk01_cellmath__39_I379 (.CO(N4187), .S(N4025), .A(a_man[19]), .B(a_man[22]), .CI(a_man[17]));
ADDFX1 inst_blk01_cellmath__39_I380 (.CO(N4034), .S(N4605), .A(a_man[21]), .B(N4528), .CI(N4025));
ADDFX1 inst_blk01_cellmath__39_I381 (.CO(N4501), .S(N4344), .A(a_man[18]), .B(a_man[20]), .CI(N4187));
ADDHX1 inst_blk01_cellmath__39_I382 (.CO(N4095), .S(N3940), .A(a_man[21]), .B(a_man[19]));
ADDHX1 inst_blk01_cellmath__39_I383 (.CO(N4408), .S(N4253), .A(a_man[22]), .B(a_man[20]));
INVXL inst_blk01_cellmath__39_I384 (.Y(N4071), .A(N4381));
NOR2XL inst_blk01_cellmath__39_I385 (.Y(N4226), .A(N3949), .B(N4273));
NAND2XL inst_blk01_cellmath__39_I386 (.Y(N4385), .A(N3949), .B(N4273));
NOR2XL inst_blk01_cellmath__39_I387 (.Y(N4537), .A(N4417), .B(N4182));
NAND2XL inst_blk01_cellmath__39_I388 (.Y(N3975), .A(N4417), .B(N4182));
NOR2XL inst_blk01_cellmath__39_I389 (.Y(N4137), .A(N4496), .B(N4335));
NAND2XL inst_blk01_cellmath__39_I390 (.Y(N4291), .A(N4335), .B(N4496));
AND2XL inst_blk01_cellmath__39_I392 (.Y(N4617), .A(N3933), .B(N4004));
NOR2XL inst_blk01_cellmath__39_I393 (.Y(N4045), .A(N4157), .B(N4635));
NAND2XL inst_blk01_cellmath__39_I394 (.Y(N4196), .A(N4157), .B(N4635));
AND2XL inst_blk01_cellmath__39_I396 (.Y(N4513), .A(N4063), .B(N4531));
NOR2XL inst_blk01_cellmath__39_I397 (.Y(N3951), .A(N3968), .B(N4131));
NAND2XL inst_blk01_cellmath__39_I398 (.Y(N4110), .A(N3968), .B(N4131));
NOR2XL inst_blk01_cellmath__39_I399 (.Y(N4265), .A(N4284), .B(N4611));
NAND2XL inst_blk01_cellmath__39_I400 (.Y(N4420), .A(N4284), .B(N4611));
NOR2XL inst_blk01_cellmath__39_I401 (.Y(N4582), .A(N4038), .B(N4349));
NOR2XL inst_blk01_cellmath__39_I403 (.Y(N4173), .A(N4505), .B(N4100));
NAND2XL inst_blk01_cellmath__39_I404 (.Y(N4327), .A(N4505), .B(N4100));
NOR2XL inst_blk01_cellmath__39_I405 (.Y(N4486), .A(N4257), .B(N4573));
NOR2XL inst_blk01_cellmath__39_I407 (.Y(N4081), .A(N4013), .B(N4231));
NAND2XL inst_blk01_cellmath__39_I408 (.Y(N4239), .A(N4013), .B(N4231));
NOR2XL inst_blk01_cellmath__39_I409 (.Y(N4396), .A(N4389), .B(N4296));
NAND2XL inst_blk01_cellmath__39_I410 (.Y(N4550), .A(N4389), .B(N4296));
NOR2XL inst_blk01_cellmath__39_I411 (.Y(N3990), .A(N4450), .B(N3955));
NAND2XL inst_blk01_cellmath__39_I412 (.Y(N4148), .A(N4450), .B(N3955));
NOR2XL inst_blk01_cellmath__39_I413 (.Y(N4301), .A(N4117), .B(N4177));
NOR2XL inst_blk01_cellmath__39_I415 (.Y(N4626), .A(N4333), .B(N4305));
NAND2XL inst_blk01_cellmath__39_I416 (.Y(N4054), .A(N4333), .B(N4305));
NOR2XL inst_blk01_cellmath__39_I417 (.Y(N3961), .A(a_man[1]), .B(a_man[0]));
AOI21XL inst_blk01_cellmath__39_I418 (.Y(N4030), .A0(N4385), .A1(N4071), .B0(N4226));
INVXL inst_blk01_cellmath__39_I419 (.Y(N4184), .A(N4385));
OAI21XL inst_blk01_cellmath__39_I420 (.Y(N4312), .A0(N4184), .A1(N3961), .B0(N4030));
AO21XL inst_blk01_cellmath__39_I421 (.Y(N4497), .A0(N4291), .A1(N4537), .B0(N4137));
AOI31X1 inst_blk01_cellmath__39_I423 (.Y(N4578), .A0(N4291), .A1(N3975), .A2(N4312), .B0(N4497));
OAI22XL inst_blk01_cellmath__39_I8415 (.Y(N4205), .A0(N4617), .A1(N4578), .B0(N3933), .B1(N4004));
AOI21XL inst_blk01_cellmath__39_I427 (.Y(N4563), .A0(N4196), .A1(N4205), .B0(N4045));
OAI22XL inst_blk01_cellmath__39_I8416 (.Y(N4101), .A0(N4513), .A1(N4563), .B0(N4063), .B1(N4531));
AO21XL inst_blk01_cellmath__39_I431 (.Y(N4546), .A0(N4420), .A1(N3951), .B0(N4265));
AOI31X1 inst_blk01_cellmath__39_I433 (.Y(N4491), .A0(N4420), .A1(N4110), .A2(N4101), .B0(N4546));
AOI21XL inst_blk01_cellmath__39_I434 (.Y(N4401), .A0(N4327), .A1(N4582), .B0(N4173));
OAI2BB1X1 inst_blk01_cellmath__39_I8417 (.Y(N4559), .A0N(N4038), .A1N(N4349), .B0(N4327));
AOI21XL inst_blk01_cellmath__39_I437 (.Y(N4306), .A0(N4239), .A1(N4486), .B0(N4081));
OAI2BB1X1 inst_blk01_cellmath__39_I8418 (.Y(N4464), .A0N(N4257), .A1N(N4573), .B0(N4239));
OAI21XL inst_blk01_cellmath__39_I442 (.Y(N4583), .A0(N4464), .A1(N4401), .B0(N4306));
NOR3XL inst_blk01_cellmath__39_I443 (.Y(N4266), .A(N4464), .B(N4559), .C(N4491));
OR2XL inst_blk01_cellmath__39_I444 (.Y(N4330), .A(N4266), .B(N4583));
AO21XL inst_blk01_cellmath__39_I445 (.Y(N3944), .A0(N4148), .A1(N4396), .B0(N3990));
AOI31X1 inst_blk01_cellmath__39_I452 (.Y(N4443), .A0(N4148), .A1(N4550), .A2(N4330), .B0(N3944));
AOI21XL inst_blk01_cellmath__39_I455 (.Y(N4356), .A0(N4054), .A1(N4301), .B0(N4626));
OAI2BB1X1 inst_blk01_cellmath__39_I8419 (.Y(N4512), .A0N(N4117), .A1N(N4177), .B0(N4054));
OAI21XL inst_blk01_cellmath__39_I458 (.Y(N3918), .A0(N4512), .A1(N4443), .B0(N4356));
NOR2XL inst_blk01_cellmath__39_I494 (.Y(N4542), .A(N4281), .B(N3941));
XOR2XL inst_blk01_cellmath__39_I495 (.Y(N3984), .A(N4281), .B(N3941));
XOR2XL inst_blk01_cellmath__39_I496 (.Y(N4295), .A(N4097), .B(N4477));
NOR2XL inst_blk01_cellmath__39_I497 (.Y(N4451), .A(N4641), .B(N4292));
XOR2XL inst_blk01_cellmath__39_I498 (.Y(N4621), .A(N4641), .B(N4292));
XOR2XL inst_blk01_cellmath__39_I499 (.Y(N4203), .A(N4446), .B(N4421));
NOR2XL inst_blk01_cellmath__39_I500 (.Y(N4364), .A(N4586), .B(N4397));
XOR2XL inst_blk01_cellmath__39_I501 (.Y(N4518), .A(N4586), .B(N4397));
XOR2XL inst_blk01_cellmath__39_I502 (.Y(N4116), .A(N4552), .B(N4124));
NOR2XL inst_blk01_cellmath__39_I503 (.Y(N4269), .A(N4278), .B(N4567));
XOR2XL inst_blk01_cellmath__39_I504 (.Y(N4426), .A(N4278), .B(N4567));
XOR2XL inst_blk01_cellmath__39_I505 (.Y(N4023), .A(N4007), .B(N4535));
NOR2XL inst_blk01_cellmath__39_I506 (.Y(N4178), .A(N3972), .B(N4263));
XOR2XL inst_blk01_cellmath__39_I507 (.Y(N4332), .A(N3972), .B(N4263));
XOR2XL inst_blk01_cellmath__39_I508 (.Y(N3930), .A(N4416), .B(N3988));
NOR2XL inst_blk01_cellmath__39_I509 (.Y(N4086), .A(N4146), .B(N4275));
XOR2XL inst_blk01_cellmath__39_I510 (.Y(N4246), .A(N4146), .B(N4275));
XOR2XL inst_blk01_cellmath__39_I511 (.Y(N4558), .A(N4430), .B(N4160));
NOR2XL inst_blk01_cellmath__39_I512 (.Y(N3996), .A(N4309), .B(N4132));
XOR2XL inst_blk01_cellmath__39_I513 (.Y(N4154), .A(N4309), .B(N4132));
XOR2XL inst_blk01_cellmath__39_I514 (.Y(N4462), .A(N4285), .B(N4259));
NOR2XL inst_blk01_cellmath__39_I515 (.Y(N4631), .A(N4413), .B(N4390));
XOR2XL inst_blk01_cellmath__39_I516 (.Y(N4060), .A(N4413), .B(N4390));
XOR2XL inst_blk01_cellmath__39_I517 (.Y(N4375), .A(N4545), .B(N4521));
NOR2XL inst_blk01_cellmath__39_I518 (.Y(N4530), .A(N3957), .B(N3932));
XOR2XL inst_blk01_cellmath__39_I519 (.Y(N3966), .A(N3957), .B(N3932));
XOR2XL inst_blk01_cellmath__39_I520 (.Y(N4282), .A(N4088), .B(N4465));
NOR2XL inst_blk01_cellmath__39_I521 (.Y(N4435), .A(N4634), .B(N4610));
XOR2XL inst_blk01_cellmath__39_I522 (.Y(N4606), .A(N4634), .B(N4610));
XOR2XL inst_blk01_cellmath__39_I523 (.Y(N4188), .A(N4036), .B(N4098));
NOR2XL inst_blk01_cellmath__39_I524 (.Y(N4346), .A(N4256), .B(N4479));
XOR2XL inst_blk01_cellmath__39_I525 (.Y(N4503), .A(N4256), .B(N4479));
XOR2XL inst_blk01_cellmath__39_I526 (.Y(N4096), .A(N4540), .B(N3917));
NOR2XL inst_blk01_cellmath__39_I527 (.Y(N4255), .A(N3979), .B(N4201));
XOR2XL inst_blk01_cellmath__39_I528 (.Y(N4409), .A(N3979), .B(N4201));
XOR2XL inst_blk01_cellmath__39_I529 (.Y(N4011), .A(N4361), .B(N4588));
NOR2XL inst_blk01_cellmath__39_I530 (.Y(N4164), .A(N4022), .B(N4245));
XOR2XL inst_blk01_cellmath__39_I531 (.Y(N4317), .A(N4022), .B(N4245));
XOR2XL inst_blk01_cellmath__39_I532 (.Y(N4640), .A(N4400), .B(N4630));
NOR2XL inst_blk01_cellmath__39_I533 (.Y(N4072), .A(N4280), .B(N4058));
XOR2XL inst_blk01_cellmath__39_I534 (.Y(N4228), .A(N4280), .B(N4058));
XOR2XL inst_blk01_cellmath__39_I535 (.Y(N4538), .A(N4434), .B(N4605));
NOR2XL inst_blk01_cellmath__39_I536 (.Y(N3977), .A(N4344), .B(N4034));
XOR2XL inst_blk01_cellmath__39_I537 (.Y(N4138), .A(N4344), .B(N4034));
XOR2XL inst_blk01_cellmath__39_I538 (.Y(N4447), .A(N3940), .B(N4501));
NOR2XL inst_blk01_cellmath__39_I539 (.Y(N4618), .A(N4095), .B(N4253));
XOR2XL inst_blk01_cellmath__39_I540 (.Y(N4046), .A(N4095), .B(N4253));
XOR2XL inst_blk01_cellmath__39_I541 (.Y(N4359), .A(N4595), .B(N4408));
XNOR2X1 inst_blk01_cellmath__39_I542 (.Y(N4152), .A(a_man[22]), .B(a_man[21]));
INVXL cmpii_A_I8511 (.Y(N19009), .A(N4463));
INVXL cmpii_A_I8512 (.Y(N19011), .A(N4128));
AND2XL cmpii_A_I8513 (.Y(N19007), .A(N19009), .B(N19011));
OAI22XL cmpii_A_I8514 (.Y(N4111), .A0(N19007), .A1(N3918), .B0(N19009), .B1(N19011));
AOI2BB2X1 inst_blk01_cellmath__39_I544 (.Y(N4422), .A0N(N4097), .A1N(N4477), .B0(N4542), .B1(N4295));
NAND2XL inst_blk01_cellmath__39_I545 (.Y(N4585), .A(N4295), .B(N3984));
AOI2BB2X1 inst_blk01_cellmath__39_I546 (.Y(N4019), .A0N(N4446), .A1N(N4421), .B0(N4451), .B1(N4203));
NAND2XL inst_blk01_cellmath__39_I547 (.Y(N4175), .A(N4203), .B(N4621));
AOI2BB2X1 inst_blk01_cellmath__39_I548 (.Y(N4328), .A0N(N4552), .A1N(N4124), .B0(N4364), .B1(N4116));
NAND2XL inst_blk01_cellmath__39_I549 (.Y(N4487), .A(N4116), .B(N4518));
AOI2BB2X1 inst_blk01_cellmath__39_I550 (.Y(N3928), .A0N(N4007), .A1N(N4535), .B0(N4269), .B1(N4023));
NAND2XL inst_blk01_cellmath__39_I551 (.Y(N4082), .A(N4023), .B(N4426));
AOI2BB2X1 inst_blk01_cellmath__39_I552 (.Y(N4240), .A0N(N4416), .A1N(N3988), .B0(N4178), .B1(N3930));
NAND2XL inst_blk01_cellmath__39_I553 (.Y(N4398), .A(N3930), .B(N4332));
AOI2BB2X1 inst_blk01_cellmath__39_I554 (.Y(N4551), .A0N(N4430), .A1N(N4160), .B0(N4086), .B1(N4558));
NAND2XL inst_blk01_cellmath__39_I555 (.Y(N3991), .A(N4558), .B(N4246));
AOI2BB2X1 inst_blk01_cellmath__39_I556 (.Y(N4150), .A0N(N4285), .A1N(N4259), .B0(N3996), .B1(N4462));
NAND2XL inst_blk01_cellmath__39_I557 (.Y(N4302), .A(N4462), .B(N4154));
AOI2BB2X1 inst_blk01_cellmath__39_I558 (.Y(N4459), .A0N(N4545), .A1N(N4521), .B0(N4631), .B1(N4375));
NAND2XL inst_blk01_cellmath__39_I559 (.Y(N4628), .A(N4375), .B(N4060));
AOI2BB2X1 inst_blk01_cellmath__39_I560 (.Y(N4055), .A0N(N4088), .A1N(N4465), .B0(N4530), .B1(N4282));
NAND2XL inst_blk01_cellmath__39_I561 (.Y(N4209), .A(N4282), .B(N3966));
AOI2BB2X1 inst_blk01_cellmath__39_I562 (.Y(N4372), .A0N(N4036), .A1N(N4098), .B0(N4435), .B1(N4188));
NAND2XL inst_blk01_cellmath__39_I563 (.Y(N4525), .A(N4188), .B(N4606));
AOI2BB2X1 inst_blk01_cellmath__39_I564 (.Y(N3962), .A0N(N4540), .A1N(N3917), .B0(N4346), .B1(N4096));
NAND2XL inst_blk01_cellmath__39_I565 (.Y(N4125), .A(N4096), .B(N4503));
AOI2BB2X1 inst_blk01_cellmath__39_I566 (.Y(N4277), .A0N(N4361), .A1N(N4588), .B0(N4255), .B1(N4011));
NAND2XL inst_blk01_cellmath__39_I567 (.Y(N4431), .A(N4011), .B(N4409));
AOI2BB2X1 inst_blk01_cellmath__39_I568 (.Y(N4602), .A0N(N4400), .A1N(N4630), .B0(N4164), .B1(N4640));
NAND2XL inst_blk01_cellmath__39_I569 (.Y(N4031), .A(N4640), .B(N4317));
AOI2BB2X1 inst_blk01_cellmath__39_I570 (.Y(N4185), .A0N(N4434), .A1N(N4605), .B0(N4072), .B1(N4538));
NAND2XL inst_blk01_cellmath__39_I571 (.Y(N4339), .A(N4538), .B(N4228));
AOI2BB2X1 inst_blk01_cellmath__39_I572 (.Y(N4498), .A0N(N3940), .A1N(N4501), .B0(N3977), .B1(N4447));
NAND2XL inst_blk01_cellmath__39_I573 (.Y(N3937), .A(N4447), .B(N4138));
OAI21XL inst_blk01_cellmath__39_I574 (.Y(N4405), .A0(N4585), .A1(N4111), .B0(N4422));
OAI21XL inst_blk01_cellmath__39_I575 (.Y(N4008), .A0(N4487), .A1(N4019), .B0(N4328));
NOR2XL inst_blk01_cellmath__39_I576 (.Y(N4161), .A(N4487), .B(N4175));
OAI21XL inst_blk01_cellmath__39_I577 (.Y(N4313), .A0(N4398), .A1(N3928), .B0(N4240));
NOR2XL inst_blk01_cellmath__39_I578 (.Y(N4473), .A(N4398), .B(N4082));
OAI21XL inst_blk01_cellmath__39_I579 (.Y(N4637), .A0(N4302), .A1(N4551), .B0(N4150));
NOR2XL inst_blk01_cellmath__39_I580 (.Y(N4068), .A(N4302), .B(N3991));
OAI21XL inst_blk01_cellmath__39_I581 (.Y(N4222), .A0(N4209), .A1(N4459), .B0(N4055));
NOR2XL inst_blk01_cellmath__39_I582 (.Y(N4382), .A(N4209), .B(N4628));
OAI21XL inst_blk01_cellmath__39_I583 (.Y(N4534), .A0(N4125), .A1(N4372), .B0(N3962));
NOR2XL inst_blk01_cellmath__39_I584 (.Y(N3973), .A(N4125), .B(N4525));
OAI21XL inst_blk01_cellmath__39_I585 (.Y(N4133), .A0(N4031), .A1(N4277), .B0(N4602));
NOR2XL inst_blk01_cellmath__39_I586 (.Y(N4288), .A(N4031), .B(N4431));
OAI21XL inst_blk01_cellmath__39_I587 (.Y(N4442), .A0(N3937), .A1(N4185), .B0(N4498));
NOR2XL inst_blk01_cellmath__39_I588 (.Y(N4615), .A(N3937), .B(N4339));
AOI21XL inst_blk01_cellmath__39_I589 (.Y(N4042), .A0(N4161), .A1(N4405), .B0(N4008));
AOI21XL inst_blk01_cellmath__39_I590 (.Y(N4354), .A0(N4068), .A1(N4313), .B0(N4637));
NAND2XL inst_blk01_cellmath__39_I591 (.Y(N4509), .A(N4068), .B(N4473));
AOI21XL inst_blk01_cellmath__39_I592 (.Y(N4262), .A0(N4615), .A1(N4133), .B0(N4442));
NAND2XL inst_blk01_cellmath__39_I593 (.Y(N4418), .A(N4615), .B(N4288));
OAI21XL inst_blk01_cellmath__39_I594 (.Y(N4579), .A0(N4509), .A1(N4042), .B0(N4354));
AO21XL inst_blk01_cellmath__39_I595 (.Y(N4324), .A0(N3973), .A1(N4222), .B0(N4534));
AOI31X1 inst_blk01_cellmath__39_I596 (.Y(N4484), .A0(N3973), .A1(N4382), .A2(N4579), .B0(N4324));
INVXL inst_blk01_cellmath__39_I597 (.Y(N4078), .A(N4473));
INVXL inst_blk01_cellmath__39_I598 (.Y(N4237), .A(N4313));
OAI21XL inst_blk01_cellmath__39_I599 (.Y(N4394), .A0(N4078), .A1(N4042), .B0(N4237));
INVXL inst_blk01_cellmath__39_I600 (.Y(N4048), .A(N4579));
AOI21XL inst_blk01_cellmath__39_I601 (.Y(N4299), .A0(N4382), .A1(N4579), .B0(N4222));
INVXL inst_blk01_cellmath__39_I602 (.Y(N4199), .A(N4484));
INVXL inst_blk01_cellmath__39_I603 (.Y(N4206), .A(N4288));
INVXL inst_blk01_cellmath__39_I604 (.Y(N4370), .A(N4133));
OAI21XL inst_blk01_cellmath__39_I605 (.Y(N4523), .A0(N4206), .A1(N4484), .B0(N4370));
OAI21XL inst_blk01_cellmath__39_I606 (.Y(N4122), .A0(N4418), .A1(N4484), .B0(N4262));
INVXL inst_blk01_cellmath__39_I607 (.Y(N4429), .A(N4175));
INVXL inst_blk01_cellmath__39_I608 (.Y(N4598), .A(N4019));
AOI21XL inst_blk01_cellmath__39_I609 (.Y(N4028), .A0(N4429), .A1(N4405), .B0(N4598));
INVXL inst_blk01_cellmath__39_I610 (.Y(N4362), .A(N4042));
OAI21XL inst_blk01_cellmath__39_I611 (.Y(N3934), .A0(N4082), .A1(N4042), .B0(N3928));
INVXL inst_blk01_cellmath__39_I612 (.Y(N4517), .A(N4394));
INVXL inst_blk01_cellmath__39_I613 (.Y(N4565), .A(N3991));
INVXL inst_blk01_cellmath__39_I614 (.Y(N4005), .A(N4551));
AOI21XL inst_blk01_cellmath__39_I615 (.Y(N4159), .A0(N4565), .A1(N4394), .B0(N4005));
INVXL inst_blk01_cellmath__39_I616 (.Y(N3954), .A(N4048));
OAI21XL inst_blk01_cellmath__39_I617 (.Y(N4066), .A0(N4628), .A1(N4048), .B0(N4459));
INVXL inst_blk01_cellmath__39_I618 (.Y(N4114), .A(N4299));
OAI21XL inst_blk01_cellmath__39_I619 (.Y(N3969), .A0(N4525), .A1(N4299), .B0(N4372));
INVXL inst_blk01_cellmath__39_I620 (.Y(N4268), .A(N4199));
INVXL inst_blk01_cellmath__39_I621 (.Y(N4612), .A(N4431));
INVXL inst_blk01_cellmath__39_I622 (.Y(N4040), .A(N4277));
AOI21XL inst_blk01_cellmath__39_I623 (.Y(N4192), .A0(N4612), .A1(N4199), .B0(N4040));
INVXL inst_blk01_cellmath__39_I624 (.Y(N4424), .A(N4523));
INVXL inst_blk01_cellmath__39_I625 (.Y(N4102), .A(N4339));
INVXL inst_blk01_cellmath__39_I626 (.Y(N4258), .A(N4185));
AOI21XL inst_blk01_cellmath__39_I627 (.Y(N4414), .A0(N4102), .A1(N4523), .B0(N4258));
INVXL inst_blk01_cellmath__39_I628 (.Y(N4589), .A(N4122));
OAI2BB2XL inst_blk01_cellmath__39_I629 (.Y(N4482), .A0N(N4618), .A1N(N4359), .B0(N4595), .B1(N4408));
AOI31X1 inst_blk01_cellmath__39_I630 (.Y(N3921), .A0(N4359), .A1(N4046), .A2(N4122), .B0(N4482));
INVXL inst_blk01_cellmath__39_I635 (.Y(N4367), .A(N4518));
INVXL inst_blk01_cellmath__39_I636 (.Y(N4520), .A(N4364));
OAI21XL inst_blk01_cellmath__39_I637 (.Y(N3956), .A0(N4367), .A1(N4028), .B0(N4520));
AOI21XL inst_blk01_cellmath__39_I638 (.Y(N4594), .A0(N4426), .A1(N4362), .B0(N4269));
AOI21XL inst_blk01_cellmath__39_I639 (.Y(N4492), .A0(N4332), .A1(N3934), .B0(N4178));
INVXL inst_blk01_cellmath__39_I640 (.Y(N4402), .A(N4246));
INVXL inst_blk01_cellmath__39_I641 (.Y(N4562), .A(N4086));
OAI21XL inst_blk01_cellmath__39_I642 (.Y(N4000), .A0(N4402), .A1(N4517), .B0(N4562));
INVXL inst_blk01_cellmath__39_I643 (.Y(N4633), .A(N4154));
INVXL inst_blk01_cellmath__39_I644 (.Y(N4062), .A(N3996));
OAI21XL inst_blk01_cellmath__39_I645 (.Y(N4214), .A0(N4633), .A1(N4159), .B0(N4062));
AOI21XL inst_blk01_cellmath__39_I646 (.Y(N4129), .A0(N4060), .A1(N3954), .B0(N4631));
AOI21XL inst_blk01_cellmath__39_I647 (.Y(N4037), .A0(N3966), .A1(N4066), .B0(N4530));
AOI21XL inst_blk01_cellmath__39_I648 (.Y(N3942), .A0(N4606), .A1(N4114), .B0(N4435));
AOI21XL inst_blk01_cellmath__39_I649 (.Y(N4570), .A0(N4503), .A1(N3969), .B0(N4346));
INVXL inst_blk01_cellmath__39_I650 (.Y(N4480), .A(N4409));
INVXL inst_blk01_cellmath__39_I651 (.Y(N3916), .A(N4255));
OAI21XL inst_blk01_cellmath__39_I652 (.Y(N4074), .A0(N4480), .A1(N4268), .B0(N3916));
INVXL inst_blk01_cellmath__39_I653 (.Y(N3981), .A(N4317));
INVXL inst_blk01_cellmath__39_I654 (.Y(N4140), .A(N4164));
OAI21XL inst_blk01_cellmath__39_I655 (.Y(N4293), .A0(N3981), .A1(N4192), .B0(N4140));
INVXL inst_blk01_cellmath__39_I656 (.Y(N4200), .A(N4228));
INVXL inst_blk01_cellmath__39_I657 (.Y(N4363), .A(N4072));
OAI21XL inst_blk01_cellmath__39_I658 (.Y(N4515), .A0(N4200), .A1(N4424), .B0(N4363));
INVXL inst_blk01_cellmath__39_I659 (.Y(N4423), .A(N4138));
INVXL inst_blk01_cellmath__39_I660 (.Y(N4590), .A(N3977));
OAI21XL inst_blk01_cellmath__39_I661 (.Y(N4021), .A0(N4423), .A1(N4414), .B0(N4590));
INVXL inst_blk01_cellmath__39_I662 (.Y(N3929), .A(N4046));
INVXL inst_blk01_cellmath__39_I663 (.Y(N4085), .A(N4618));
OAI21XL inst_blk01_cellmath__39_I664 (.Y(N4244), .A0(N3929), .A1(N4589), .B0(N4085));
XNOR2X1 inst_blk01_cellmath__39_I671 (.Y(N608), .A(N3956), .B(N4116));
XNOR2X1 inst_blk01_cellmath__39_I672 (.Y(N609), .A(N4362), .B(N4426));
XOR2XL inst_blk01_cellmath__39_I673 (.Y(N610), .A(N4594), .B(N4023));
XNOR2X1 inst_blk01_cellmath__39_I674 (.Y(N611), .A(N3934), .B(N4332));
XOR2XL inst_blk01_cellmath__39_I675 (.Y(N612), .A(N4492), .B(N3930));
XOR2XL inst_blk01_cellmath__39_I676 (.Y(N613), .A(N4517), .B(N4246));
XNOR2X1 inst_blk01_cellmath__39_I677 (.Y(N614), .A(N4000), .B(N4558));
XOR2XL inst_blk01_cellmath__39_I678 (.Y(N615), .A(N4159), .B(N4154));
XNOR2X1 inst_blk01_cellmath__39_I679 (.Y(N616), .A(N4214), .B(N4462));
XNOR2X1 inst_blk01_cellmath__39_I680 (.Y(N617), .A(N3954), .B(N4060));
XOR2XL inst_blk01_cellmath__39_I681 (.Y(N618), .A(N4129), .B(N4375));
XNOR2X1 inst_blk01_cellmath__39_I682 (.Y(N619), .A(N4066), .B(N3966));
XOR2XL inst_blk01_cellmath__39_I683 (.Y(N620), .A(N4037), .B(N4282));
XNOR2X1 inst_blk01_cellmath__39_I684 (.Y(N621), .A(N4114), .B(N4606));
XOR2XL inst_blk01_cellmath__39_I685 (.Y(N622), .A(N3942), .B(N4188));
XNOR2X1 inst_blk01_cellmath__39_I686 (.Y(N623), .A(N3969), .B(N4503));
XOR2XL inst_blk01_cellmath__39_I687 (.Y(N624), .A(N4570), .B(N4096));
XOR2XL inst_blk01_cellmath__39_I688 (.Y(N625), .A(N4268), .B(N4409));
XNOR2X1 inst_blk01_cellmath__39_I689 (.Y(N626), .A(N4074), .B(N4011));
XOR2XL inst_blk01_cellmath__39_I690 (.Y(N627), .A(N4192), .B(N4317));
XNOR2X1 inst_blk01_cellmath__39_I691 (.Y(N628), .A(N4293), .B(N4640));
XOR2XL inst_blk01_cellmath__39_I692 (.Y(N629), .A(N4424), .B(N4228));
XNOR2X1 inst_blk01_cellmath__39_I693 (.Y(N630), .A(N4515), .B(N4538));
XOR2XL inst_blk01_cellmath__39_I694 (.Y(N631), .A(N4414), .B(N4138));
XNOR2X1 inst_blk01_cellmath__39_I695 (.Y(N632), .A(N4021), .B(N4447));
XOR2XL inst_blk01_cellmath__39_I696 (.Y(N633), .A(N4589), .B(N4046));
XNOR2X1 inst_blk01_cellmath__39_I697 (.Y(N634), .A(N4244), .B(N4359));
XNOR2X1 inst_blk01_cellmath__39_I698 (.Y(N635), .A(N3921), .B(N4152));
OA22X1 inst_blk01_cellmath__39_I699 (.Y(N637), .A0(N4152), .A1(N3921), .B0(a_man[22]), .B1(a_man[21]));
INVXL inst_blk01_cellmath__39_I700 (.Y(N636), .A(N637));
INVXL inst_cellmath__42_0_I701 (.Y(inst_cellmath__42[0]), .A(a_exp[0]));
INVXL inst_cellmath__42_0_I702 (.Y(N5345), .A(a_exp[1]));
INVXL inst_cellmath__42_0_I703 (.Y(N5360), .A(a_exp[3]));
NAND2BXL inst_cellmath__42_0_I704 (.Y(N5349), .AN(N5345), .B(a_exp[2]));
NAND2XL inst_cellmath__42_0_I705 (.Y(N5348), .A(N5360), .B(N5349));
NOR2XL inst_cellmath__42_0_I706 (.Y(N5347), .A(a_exp[4]), .B(N5348));
INVXL inst_cellmath__42_0_I707 (.Y(inst_cellmath__42[1]), .A(N5345));
XOR2XL inst_cellmath__42_0_I710 (.Y(inst_cellmath__42[4]), .A(N5348), .B(a_exp[4]));
XNOR2X1 inst_cellmath__42_0_I711 (.Y(inst_cellmath__42[5]), .A(N5347), .B(a_exp[5]));
INVXL inst_cellmath__48_I712 (.Y(N5493), .A(inst_cellmath__42[0]));
AOI22XL inst_cellmath__48_I713 (.Y(N5410), .A0(inst_cellmath__42[0]), .A1(N609), .B0(N608), .B1(N5493));
AOI22XL inst_cellmath__48_I714 (.Y(N5456), .A0(inst_cellmath__42[0]), .A1(N610), .B0(N609), .B1(N5493));
AOI22XL inst_cellmath__48_I715 (.Y(N5502), .A0(inst_cellmath__42[0]), .A1(N611), .B0(N610), .B1(N5493));
AOI22XL inst_cellmath__48_I716 (.Y(N5549), .A0(inst_cellmath__42[0]), .A1(N612), .B0(N611), .B1(N5493));
AOI22XL inst_cellmath__48_I717 (.Y(N5383), .A0(inst_cellmath__42[0]), .A1(N613), .B0(N612), .B1(N5493));
AOI22XL inst_cellmath__48_I718 (.Y(N5429), .A0(inst_cellmath__42[0]), .A1(N614), .B0(N613), .B1(N5493));
AOI22XL inst_cellmath__48_I719 (.Y(N5474), .A0(inst_cellmath__42[0]), .A1(N615), .B0(N614), .B1(N5493));
AOI22XL inst_cellmath__48_I720 (.Y(N5521), .A0(inst_cellmath__42[0]), .A1(N616), .B0(N615), .B1(N5493));
AOI22XL inst_cellmath__48_I721 (.Y(N5567), .A0(inst_cellmath__42[0]), .A1(N617), .B0(N616), .B1(N5493));
AOI22XL inst_cellmath__48_I722 (.Y(N5402), .A0(inst_cellmath__42[0]), .A1(N618), .B0(N617), .B1(N5493));
AOI22XL inst_cellmath__48_I723 (.Y(N5449), .A0(inst_cellmath__42[0]), .A1(N619), .B0(N618), .B1(N5493));
AOI22XL inst_cellmath__48_I724 (.Y(N5495), .A0(inst_cellmath__42[0]), .A1(N620), .B0(N619), .B1(N5493));
AOI22XL inst_cellmath__48_I725 (.Y(N5542), .A0(inst_cellmath__42[0]), .A1(N621), .B0(N620), .B1(N5493));
AOI22XL inst_cellmath__48_I726 (.Y(N5375), .A0(inst_cellmath__42[0]), .A1(N622), .B0(N621), .B1(N5493));
AOI22XL inst_cellmath__48_I727 (.Y(N5422), .A0(inst_cellmath__42[0]), .A1(N623), .B0(N622), .B1(N5493));
AOI22XL inst_cellmath__48_I728 (.Y(N5468), .A0(inst_cellmath__42[0]), .A1(N624), .B0(N623), .B1(N5493));
AOI22XL inst_cellmath__48_I729 (.Y(N5516), .A0(inst_cellmath__42[0]), .A1(N625), .B0(N624), .B1(N5493));
AOI22XL inst_cellmath__48_I730 (.Y(N5561), .A0(inst_cellmath__42[0]), .A1(N626), .B0(N625), .B1(N5493));
AOI22XL inst_cellmath__48_I731 (.Y(N5395), .A0(inst_cellmath__42[0]), .A1(N627), .B0(N626), .B1(N5493));
AOI22XL inst_cellmath__48_I732 (.Y(N5443), .A0(inst_cellmath__42[0]), .A1(N628), .B0(N627), .B1(N5493));
AOI22XL inst_cellmath__48_I733 (.Y(N5486), .A0(inst_cellmath__42[0]), .A1(N629), .B0(N628), .B1(N5493));
AOI22XL inst_cellmath__48_I734 (.Y(N5534), .A0(inst_cellmath__42[0]), .A1(N630), .B0(N629), .B1(N5493));
AOI22XL inst_cellmath__48_I735 (.Y(N5581), .A0(inst_cellmath__42[0]), .A1(N631), .B0(N630), .B1(N5493));
AOI22XL inst_cellmath__48_I736 (.Y(N5415), .A0(inst_cellmath__42[0]), .A1(N632), .B0(N631), .B1(N5493));
AOI22XL inst_cellmath__48_I737 (.Y(N5460), .A0(inst_cellmath__42[0]), .A1(N633), .B0(N632), .B1(N5493));
AOI22XL inst_cellmath__48_I738 (.Y(N5506), .A0(inst_cellmath__42[0]), .A1(N634), .B0(N633), .B1(N5493));
AOI22XL inst_cellmath__48_I739 (.Y(N5553), .A0(inst_cellmath__42[0]), .A1(N635), .B0(N634), .B1(N5493));
AOI22XL inst_cellmath__48_I740 (.Y(N5386), .A0(inst_cellmath__42[0]), .A1(N636), .B0(N635), .B1(N5493));
AOI22XL inst_cellmath__48_I741 (.Y(N5434), .A0(inst_cellmath__42[0]), .A1(N637), .B0(N636), .B1(N5493));
NAND2XL inst_cellmath__48_I742 (.Y(N5478), .A(N637), .B(N5493));
INVXL inst_cellmath__48_I743 (.Y(N5540), .A(inst_cellmath__42[1]));
INVXL inst_cellmath__48_I744 (.Y(N5531), .A(N5540));
AOI22XL inst_cellmath__48_I745 (.Y(N5447), .A0(N5540), .A1(N5410), .B0(N5502), .B1(N5531));
AOI22XL inst_cellmath__48_I746 (.Y(N5494), .A0(N5540), .A1(N5456), .B0(N5549), .B1(N5531));
AOI22XL inst_cellmath__48_I747 (.Y(N5541), .A0(N5540), .A1(N5502), .B0(N5383), .B1(N5531));
AOI22XL inst_cellmath__48_I748 (.Y(N5373), .A0(N5540), .A1(N5549), .B0(N5429), .B1(N5531));
AOI22XL inst_cellmath__48_I749 (.Y(N5421), .A0(N5540), .A1(N5383), .B0(N5474), .B1(N5531));
AOI22XL inst_cellmath__48_I750 (.Y(N5467), .A0(N5540), .A1(N5429), .B0(N5521), .B1(N5531));
AOI22XL inst_cellmath__48_I751 (.Y(N5514), .A0(N5540), .A1(N5474), .B0(N5567), .B1(N5531));
AOI22XL inst_cellmath__48_I752 (.Y(N5560), .A0(N5540), .A1(N5521), .B0(N5402), .B1(N5531));
AOI22XL inst_cellmath__48_I753 (.Y(N5394), .A0(N5540), .A1(N5567), .B0(N5449), .B1(N5531));
AOI22XL inst_cellmath__48_I754 (.Y(N5441), .A0(N5540), .A1(N5402), .B0(N5495), .B1(N5531));
AOI22XL inst_cellmath__48_I755 (.Y(N5485), .A0(N5540), .A1(N5449), .B0(N5542), .B1(N5531));
AOI22XL inst_cellmath__48_I756 (.Y(N5533), .A0(N5540), .A1(N5495), .B0(N5375), .B1(N5531));
AOI22XL inst_cellmath__48_I757 (.Y(N5578), .A0(N5540), .A1(N5542), .B0(N5422), .B1(N5531));
AOI22XL inst_cellmath__48_I758 (.Y(N5414), .A0(N5540), .A1(N5375), .B0(N5468), .B1(N5531));
AOI22XL inst_cellmath__48_I759 (.Y(N5459), .A0(N5540), .A1(N5422), .B0(N5516), .B1(N5531));
AOI22XL inst_cellmath__48_I760 (.Y(N5504), .A0(N5540), .A1(N5468), .B0(N5561), .B1(N5531));
AOI22XL inst_cellmath__48_I761 (.Y(N5552), .A0(N5540), .A1(N5516), .B0(N5395), .B1(N5531));
AOI22XL inst_cellmath__48_I762 (.Y(N5385), .A0(N5540), .A1(N5561), .B0(N5443), .B1(N5531));
AOI22XL inst_cellmath__48_I763 (.Y(N5432), .A0(N5540), .A1(N5395), .B0(N5486), .B1(N5531));
AOI22XL inst_cellmath__48_I764 (.Y(N5476), .A0(N5540), .A1(N5443), .B0(N5534), .B1(N5531));
AOI22XL inst_cellmath__48_I765 (.Y(N5525), .A0(N5540), .A1(N5486), .B0(N5581), .B1(N5531));
AOI22XL inst_cellmath__48_I766 (.Y(N5570), .A0(N5540), .A1(N5534), .B0(N5415), .B1(N5531));
AOI22XL inst_cellmath__48_I767 (.Y(N5404), .A0(N5540), .A1(N5581), .B0(N5460), .B1(N5531));
AOI22XL inst_cellmath__48_I768 (.Y(N5451), .A0(N5540), .A1(N5415), .B0(N5506), .B1(N5531));
AOI22XL inst_cellmath__48_I769 (.Y(N5497), .A0(N5540), .A1(N5460), .B0(N5553), .B1(N5531));
AOI22XL inst_cellmath__48_I770 (.Y(N5544), .A0(N5540), .A1(N5506), .B0(N5386), .B1(N5531));
AOI22XL inst_cellmath__48_I771 (.Y(N5377), .A0(N5540), .A1(N5553), .B0(N5434), .B1(N5531));
AOI22XL inst_cellmath__48_I772 (.Y(N5425), .A0(N5540), .A1(N5386), .B0(N5478), .B1(N5531));
NOR2XL inst_cellmath__48_I773 (.Y(N5470), .A(N5531), .B(N5434));
NOR2XL inst_cellmath__48_I774 (.Y(N5397), .A(N5531), .B(N5478));
XOR2XL inst_cellmath__48_I8421 (.Y(N5568), .A(inst_cellmath__42[1]), .B(a_exp[2]));
INVXL inst_cellmath__48_I776 (.Y(N5562), .A(N5568));
AOI22XL inst_cellmath__48_I777 (.Y(N5527), .A0(N5562), .A1(N5421), .B0(N5447), .B1(N5568));
AOI22XL inst_cellmath__48_I778 (.Y(N5573), .A0(N5562), .A1(N5467), .B0(N5494), .B1(N5568));
AOI22XL inst_cellmath__48_I779 (.Y(N5406), .A0(N5562), .A1(N5514), .B0(N5541), .B1(N5568));
AOI22XL inst_cellmath__48_I780 (.Y(N5453), .A0(N5562), .A1(N5560), .B0(N5373), .B1(N5568));
AOI22XL inst_cellmath__48_I781 (.Y(N5499), .A0(N5562), .A1(N5394), .B0(N5421), .B1(N5568));
AOI22XL inst_cellmath__48_I782 (.Y(N5547), .A0(N5562), .A1(N5441), .B0(N5467), .B1(N5568));
AOI22XL inst_cellmath__48_I783 (.Y(N5381), .A0(N5562), .A1(N5485), .B0(N5514), .B1(N5568));
AOI22XL inst_cellmath__48_I784 (.Y(N5427), .A0(N5562), .A1(N5533), .B0(N5560), .B1(N5568));
AOI22XL inst_cellmath__48_I785 (.Y(N5472), .A0(N5562), .A1(N5578), .B0(N5394), .B1(N5568));
AOI22XL inst_cellmath__48_I786 (.Y(N5519), .A0(N5562), .A1(N5414), .B0(N5441), .B1(N5568));
AOI22XL inst_cellmath__48_I787 (.Y(N5565), .A0(N5562), .A1(N5459), .B0(N5485), .B1(N5568));
AOI22XL inst_cellmath__48_I788 (.Y(N5399), .A0(N5562), .A1(N5504), .B0(N5533), .B1(N5568));
AOI22XL inst_cellmath__48_I789 (.Y(N5446), .A0(N5562), .A1(N5552), .B0(N5578), .B1(N5568));
AOI22XL inst_cellmath__48_I790 (.Y(N5492), .A0(N5562), .A1(N5385), .B0(N5414), .B1(N5568));
AOI22XL inst_cellmath__48_I791 (.Y(N5539), .A0(N5562), .A1(N5432), .B0(N5459), .B1(N5568));
AOI22XL inst_cellmath__48_I792 (.Y(N5586), .A0(N5562), .A1(N5476), .B0(N5504), .B1(N5568));
AOI22XL inst_cellmath__48_I793 (.Y(N5420), .A0(N5562), .A1(N5525), .B0(N5552), .B1(N5568));
AOI22XL inst_cellmath__48_I794 (.Y(N5465), .A0(N5562), .A1(N5570), .B0(N5385), .B1(N5568));
AOI22XL inst_cellmath__48_I795 (.Y(N5511), .A0(N5562), .A1(N5404), .B0(N5432), .B1(N5568));
AOI22XL inst_cellmath__48_I796 (.Y(N5558), .A0(N5562), .A1(N5451), .B0(N5476), .B1(N5568));
AOI22XL inst_cellmath__48_I797 (.Y(N5392), .A0(N5562), .A1(N5497), .B0(N5525), .B1(N5568));
AOI22XL inst_cellmath__48_I798 (.Y(N5439), .A0(N5562), .A1(N5544), .B0(N5570), .B1(N5568));
AOI22XL inst_cellmath__48_I799 (.Y(N5483), .A0(N5562), .A1(N5377), .B0(N5404), .B1(N5568));
AOI22XL inst_cellmath__48_I800 (.Y(N5530), .A0(N5562), .A1(N5425), .B0(N5451), .B1(N5568));
AOI22XL inst_cellmath__48_I801 (.Y(N5576), .A0(N5562), .A1(N5470), .B0(N5497), .B1(N5568));
AOI22XL inst_cellmath__48_I802 (.Y(N5411), .A0(N5562), .A1(N5397), .B0(N5544), .B1(N5568));
NAND2XL inst_cellmath__48_I803 (.Y(N5457), .A(N5377), .B(N5568));
NAND2XL inst_cellmath__48_I804 (.Y(N5550), .A(N5425), .B(N5568));
NAND2XL inst_cellmath__48_I805 (.Y(N5430), .A(N5470), .B(N5568));
NAND2XL inst_cellmath__48_I806 (.Y(N5522), .A(N5397), .B(N5568));
XNOR2X1 inst_cellmath__48_I8422 (.Y(N5545), .A(N5349), .B(N5360));
INVXL inst_cellmath__48_I808 (.Y(N5379), .A(N5545));
AOI22XL inst_cellmath__48_I809 (.Y(N5490), .A0(N5545), .A1(N5527), .B0(N5472), .B1(N5379));
AOI22XL inst_cellmath__48_I810 (.Y(N5537), .A0(N5545), .A1(N5573), .B0(N5519), .B1(N5379));
AOI22XL inst_cellmath__48_I811 (.Y(N5584), .A0(N5545), .A1(N5406), .B0(N5565), .B1(N5379));
AOI22XL inst_cellmath__48_I812 (.Y(N5418), .A0(N5545), .A1(N5453), .B0(N5399), .B1(N5379));
AOI22XL inst_cellmath__48_I813 (.Y(N5463), .A0(N5545), .A1(N5499), .B0(N5446), .B1(N5379));
AOI22XL inst_cellmath__48_I814 (.Y(N5509), .A0(N5545), .A1(N5547), .B0(N5492), .B1(N5379));
AOI22XL inst_cellmath__48_I815 (.Y(N5556), .A0(N5545), .A1(N5381), .B0(N5539), .B1(N5379));
AOI22XL inst_cellmath__48_I816 (.Y(N5390), .A0(N5545), .A1(N5427), .B0(N5586), .B1(N5379));
AOI22XL inst_cellmath__48_I817 (.Y(N5437), .A0(N5545), .A1(N5472), .B0(N5420), .B1(N5379));
AOI22XL inst_cellmath__48_I818 (.Y(N5481), .A0(N5545), .A1(N5519), .B0(N5465), .B1(N5379));
AOI22XL inst_cellmath__48_I819 (.Y(N5529), .A0(N5545), .A1(N5565), .B0(N5511), .B1(N5379));
AOI22XL inst_cellmath__48_I820 (.Y(N5575), .A0(N5545), .A1(N5399), .B0(N5558), .B1(N5379));
AOI22XL inst_cellmath__48_I821 (.Y(N5408), .A0(N5545), .A1(N5446), .B0(N5392), .B1(N5379));
AOI22XL inst_cellmath__48_I822 (.Y(N5455), .A0(N5545), .A1(N5492), .B0(N5439), .B1(N5379));
AOI22XL inst_cellmath__48_I823 (.Y(N5501), .A0(N5545), .A1(N5539), .B0(N5483), .B1(N5379));
AOI22XL inst_cellmath__48_I824 (.Y(N5548), .A0(N5545), .A1(N5586), .B0(N5530), .B1(N5379));
AOI22XL inst_cellmath__48_I825 (.Y(N5382), .A0(N5545), .A1(N5420), .B0(N5576), .B1(N5379));
AOI22XL inst_cellmath__48_I826 (.Y(N5428), .A0(N5545), .A1(N5465), .B0(N5411), .B1(N5379));
AOI22XL inst_cellmath__48_I827 (.Y(N5473), .A0(N5545), .A1(N5511), .B0(N5457), .B1(N5379));
AOI22XL inst_cellmath__48_I828 (.Y(N5520), .A0(N5545), .A1(N5558), .B0(N5550), .B1(N5379));
AOI22XL inst_cellmath__48_I829 (.Y(N5566), .A0(N5545), .A1(N5392), .B0(N5430), .B1(N5379));
AOI22XL inst_cellmath__48_I830 (.Y(N5401), .A0(N5545), .A1(N5439), .B0(N5522), .B1(N5379));
NOR2XL inst_cellmath__48_I831 (.Y(N5448), .A(N5379), .B(N5483));
NOR2XL inst_cellmath__48_I832 (.Y(N5374), .A(N5379), .B(N5530));
NOR2XL inst_cellmath__48_I833 (.Y(N5515), .A(N5379), .B(N5576));
NOR2XL inst_cellmath__48_I834 (.Y(N5442), .A(N5379), .B(N5411));
NOR2XL inst_cellmath__48_I835 (.Y(N5579), .A(N5379), .B(N5457));
NOR2XL inst_cellmath__48_I836 (.Y(N5505), .A(N5379), .B(N5550));
NOR2XL inst_cellmath__48_I837 (.Y(N5433), .A(N5379), .B(N5430));
NOR2XL inst_cellmath__48_I838 (.Y(N5571), .A(N5379), .B(N5522));
INVXL inst_cellmath__48_I839 (.Y(N5409), .A(inst_cellmath__42[4]));
AOI22XL inst_cellmath__48_I840 (.Y(N5488), .A0(inst_cellmath__42[4]), .A1(N5382), .B0(N5490), .B1(N5409));
AOI22XL inst_cellmath__48_I841 (.Y(N5536), .A0(inst_cellmath__42[4]), .A1(N5428), .B0(N5537), .B1(N5409));
AOI22XL inst_cellmath__48_I842 (.Y(N5583), .A0(inst_cellmath__42[4]), .A1(N5473), .B0(N5584), .B1(N5409));
AOI22XL inst_cellmath__48_I843 (.Y(N5417), .A0(inst_cellmath__42[4]), .A1(N5520), .B0(N5418), .B1(N5409));
AOI22XL inst_cellmath__48_I844 (.Y(N5462), .A0(inst_cellmath__42[4]), .A1(N5566), .B0(N5463), .B1(N5409));
AOI22XL inst_cellmath__48_I845 (.Y(N5508), .A0(inst_cellmath__42[4]), .A1(N5401), .B0(N5509), .B1(N5409));
AOI22XL inst_cellmath__48_I846 (.Y(N5555), .A0(inst_cellmath__42[4]), .A1(N5448), .B0(N5556), .B1(N5409));
AOI22XL inst_cellmath__48_I847 (.Y(N5388), .A0(inst_cellmath__42[4]), .A1(N5374), .B0(N5390), .B1(N5409));
AOI22XL inst_cellmath__48_I848 (.Y(N5436), .A0(inst_cellmath__42[4]), .A1(N5515), .B0(N5437), .B1(N5409));
AOI22XL inst_cellmath__48_I849 (.Y(N5480), .A0(inst_cellmath__42[4]), .A1(N5442), .B0(N5481), .B1(N5409));
AOI22XL inst_cellmath__48_I850 (.Y(N5528), .A0(inst_cellmath__42[4]), .A1(N5579), .B0(N5529), .B1(N5409));
AOI22XL inst_cellmath__48_I851 (.Y(N5574), .A0(inst_cellmath__42[4]), .A1(N5505), .B0(N5575), .B1(N5409));
AOI22XL inst_cellmath__48_I852 (.Y(N5407), .A0(inst_cellmath__42[4]), .A1(N5433), .B0(N5408), .B1(N5409));
AOI22XL inst_cellmath__48_I853 (.Y(N5454), .A0(inst_cellmath__42[4]), .A1(N5571), .B0(N5455), .B1(N5409));
NOR2XL inst_cellmath__48_I854 (.Y(N733), .A(inst_cellmath__42[5]), .B(N5488));
NOR2XL inst_cellmath__48_I855 (.Y(N734), .A(inst_cellmath__42[5]), .B(N5536));
NOR2XL inst_cellmath__48_I856 (.Y(N735), .A(inst_cellmath__42[5]), .B(N5583));
NOR2XL inst_cellmath__48_I857 (.Y(N736), .A(inst_cellmath__42[5]), .B(N5417));
NOR2XL inst_cellmath__48_I858 (.Y(N737), .A(inst_cellmath__42[5]), .B(N5462));
NOR2XL inst_cellmath__48_I859 (.Y(N738), .A(inst_cellmath__42[5]), .B(N5508));
NOR2XL inst_cellmath__48_I860 (.Y(N739), .A(inst_cellmath__42[5]), .B(N5555));
NOR2XL inst_cellmath__48_I861 (.Y(N740), .A(inst_cellmath__42[5]), .B(N5388));
NOR2XL inst_cellmath__48_I862 (.Y(N741), .A(inst_cellmath__42[5]), .B(N5436));
NOR2XL inst_cellmath__48_I863 (.Y(N742), .A(inst_cellmath__42[5]), .B(N5480));
NOR2XL inst_cellmath__48_I864 (.Y(N743), .A(inst_cellmath__42[5]), .B(N5528));
NOR2XL inst_cellmath__48_I865 (.Y(N744), .A(inst_cellmath__42[5]), .B(N5574));
NOR2XL inst_cellmath__48_I866 (.Y(N745), .A(inst_cellmath__42[5]), .B(N5407));
NOR2XL inst_cellmath__48_I867 (.Y(N746), .A(inst_cellmath__42[5]), .B(N5454));
NAND2XL inst_cellmath__48_I868 (.Y(N5580), .A(N5501), .B(N5409));
NOR2XL inst_cellmath__48_I869 (.Y(N747), .A(inst_cellmath__42[5]), .B(N5580));
NAND2XL inst_cellmath__48_I870 (.Y(N5477), .A(N5548), .B(N5409));
NOR2XL inst_cellmath__48_I871 (.Y(N748), .A(inst_cellmath__42[5]), .B(N5477));
NAND2XL inst_cellmath__48_I872 (.Y(N5378), .A(N5382), .B(N5409));
NOR2XL inst_cellmath__48_I873 (.Y(N749), .A(inst_cellmath__42[5]), .B(N5378));
NAND2XL inst_cellmath__48_I874 (.Y(N5489), .A(N5428), .B(N5409));
NOR2XL inst_cellmath__48_I875 (.Y(N750), .A(inst_cellmath__42[5]), .B(N5489));
NAND2XL inst_cellmath__48_I876 (.Y(N5389), .A(N5473), .B(N5409));
NOR2XL inst_cellmath__48_I877 (.Y(N751), .A(inst_cellmath__42[5]), .B(N5389));
NAND2XL inst_cellmath__48_I878 (.Y(N5500), .A(N5520), .B(N5409));
NOR2XL inst_cellmath__48_I879 (.Y(N752), .A(inst_cellmath__42[5]), .B(N5500));
NAND2XL inst_cellmath__48_I880 (.Y(N5400), .A(N5566), .B(N5409));
NOR2XL inst_cellmath__48_I881 (.Y(N753), .A(inst_cellmath__42[5]), .B(N5400));
NAND2XL inst_cellmath__48_I882 (.Y(N5513), .A(N5401), .B(N5409));
NOR2XL inst_cellmath__48_I883 (.Y(N754), .A(inst_cellmath__42[5]), .B(N5513));
NAND2XL inst_cellmath__48_I884 (.Y(N5413), .A(N5448), .B(N5409));
NOR2XL inst_cellmath__48_I885 (.Y(N755), .A(inst_cellmath__42[5]), .B(N5413));
NAND2XL inst_cellmath__48_I886 (.Y(N5524), .A(N5374), .B(N5409));
NAND2XL inst_cellmath__48_I888 (.Y(N5424), .A(N5515), .B(N5409));
NOR2XL inst_cellmath__48_I889 (.Y(N757), .A(inst_cellmath__42[5]), .B(N5424));
OR2XL inst_cellmath__61_0_I8423 (.Y(N5778), .A(inst_cellmath__42[5]), .B(N5524));
XNOR2X1 inst_cellmath__61_0_I892 (.Y(inst_cellmath__61[1]), .A(N734), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I893 (.Y(inst_cellmath__61[2]), .A(N735), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I894 (.Y(inst_cellmath__61[3]), .A(N736), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I895 (.Y(inst_cellmath__61[4]), .A(N737), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I896 (.Y(inst_cellmath__61[5]), .A(N738), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I897 (.Y(inst_cellmath__61[6]), .A(N739), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I898 (.Y(inst_cellmath__61[7]), .A(N740), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I899 (.Y(inst_cellmath__61[8]), .A(N741), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I900 (.Y(inst_cellmath__61[9]), .A(N742), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I901 (.Y(inst_cellmath__61[10]), .A(N743), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I902 (.Y(inst_cellmath__61[11]), .A(N744), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I903 (.Y(inst_cellmath__61[12]), .A(N745), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I904 (.Y(inst_cellmath__61[13]), .A(N746), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I905 (.Y(inst_cellmath__61[14]), .A(N747), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I906 (.Y(inst_cellmath__61[15]), .A(N748), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I908 (.Y(inst_cellmath__61[17]), .A(N750), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I909 (.Y(inst_cellmath__61[18]), .A(N751), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I910 (.Y(inst_cellmath__61[19]), .A(N752), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I911 (.Y(inst_cellmath__61[20]), .A(N753), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I912 (.Y(inst_cellmath__61[21]), .A(N754), .B(N5778));
XNOR2X1 inst_cellmath__61_0_I913 (.Y(inst_cellmath__61[22]), .A(N755), .B(N5778));
XOR2XL cynw_cm_float_sin_I8424 (.Y(inst_cellmath__115__W1[0]), .A(N749), .B(N5778));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I914 (.Y(N6300), .A(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I915 (.Y(N6574), .A(inst_cellmath__61[20]), .B(inst_cellmath__61[21]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I916 (.Y(N6329), .A(N6574), .B(N6300));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I917 (.Y(N6008), .A(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I918 (.Y(N6299), .A(inst_cellmath__61[17]), .B(inst_cellmath__61[18]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I919 (.Y(N5840), .A(N6299), .B(N6008));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I920 (.Y(N6653), .A(N5840), .B(N6329));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I921 (.Y(N6006), .A(inst_cellmath__61[17]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I922 (.Y(N6187), .A(N6006), .B(inst_cellmath__61[18]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I923 (.Y(N6215), .A(N6187), .B(N6008));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I924 (.Y(N6540), .A(N6215), .B(N6329));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I925 (.Y(N5891), .A(inst_cellmath__61[18]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I926 (.Y(N6076), .A(inst_cellmath__61[17]), .B(N5891));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I927 (.Y(N6568), .A(N6076), .B(N6008));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I928 (.Y(N6442), .A(N6568), .B(N6329));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I929 (.Y(N6621), .A(N6006), .B(N5891));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I930 (.Y(N6106), .A(N6621), .B(N6008));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I931 (.Y(N6159), .A(N6106), .B(N6329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I932 (.Y(N6466), .A(N6299), .B(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I933 (.Y(N6511), .A(N6466), .B(N6329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I934 (.Y(N6002), .A(N6187), .B(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I935 (.Y(N6047), .A(N6002), .B(N6329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I936 (.Y(N6365), .A(N6076), .B(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I937 (.Y(N6406), .A(N6365), .B(N6329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I938 (.Y(N5885), .A(N6621), .B(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I939 (.Y(N5944), .A(N5885), .B(N6329));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I940 (.Y(N6130), .A(inst_cellmath__61[20]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I941 (.Y(N6317), .A(N6130), .B(inst_cellmath__61[21]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I942 (.Y(N6264), .A(N6317), .B(N6300));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I943 (.Y(N6670), .A(N5840), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I944 (.Y(N6022), .A(N6215), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I945 (.Y(N6200), .A(N6568), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I946 (.Y(N6380), .A(N6106), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I947 (.Y(N6555), .A(N6466), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I948 (.Y(N5905), .A(N6002), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I949 (.Y(N6093), .A(N6365), .B(N6264));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I950 (.Y(N6284), .A(N5885), .B(N6264));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I951 (.Y(N6456), .A(inst_cellmath__61[21]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I952 (.Y(N6634), .A(inst_cellmath__61[20]), .B(N6456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I953 (.Y(N6614), .A(N6634), .B(N6300));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I954 (.Y(N6172), .A(N5840), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I955 (.Y(N6152), .A(N6215), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I956 (.Y(N6523), .A(N6568), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I957 (.Y(N6503), .A(N6106), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I958 (.Y(N6042), .A(N6466), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I959 (.Y(N6402), .A(N6002), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I960 (.Y(N6422), .A(N6365), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I961 (.Y(N6605), .A(N5885), .B(N6614));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I962 (.Y(N5957), .A(N6130), .B(N6456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I963 (.Y(N5939), .A(N5957), .B(N6300));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I964 (.Y(N6332), .A(N5840), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I965 (.Y(N6496), .A(N6215), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I966 (.Y(N5842), .A(N6568), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I967 (.Y(N6031), .A(N6106), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I968 (.Y(N6217), .A(N6466), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I969 (.Y(N6389), .A(N6002), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I970 (.Y(N6310), .A(N6365), .B(N5939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I971 (.Y(N5923), .A(N5885), .B(N5939));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I972 (.Y(N6662), .A(N6574), .B(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I973 (.Y(N6295), .A(N5840), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I974 (.Y(N6193), .A(N6215), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I975 (.Y(N6649), .A(N6568), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I976 (.Y(N6004), .A(N6106), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I977 (.Y(N6185), .A(N6466), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I978 (.Y(N6366), .A(N6002), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I979 (.Y(N6547), .A(N6365), .B(N6662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I980 (.Y(N5888), .A(N5885), .B(N6662));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I981 (.Y(N6087), .A(N6317), .B(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I982 (.Y(N6266), .A(N5840), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I983 (.Y(N6437), .A(N6215), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I984 (.Y(N6616), .A(N6568), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I985 (.Y(N5974), .A(N6106), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I986 (.Y(N6154), .A(N6466), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I987 (.Y(N6343), .A(N6002), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I988 (.Y(N6451), .A(N6365), .B(N6087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I989 (.Y(N5855), .A(N5885), .B(N6087));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I990 (.Y(N5988), .A(N6634), .B(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I991 (.Y(N6233), .A(N5840), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I992 (.Y(N6403), .A(N6215), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I993 (.Y(N6589), .A(N6568), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I994 (.Y(N6352), .A(N6106), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I995 (.Y(N6124), .A(N6466), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I996 (.Y(N6312), .A(N6002), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I997 (.Y(N6481), .A(N6365), .B(N5988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I998 (.Y(N6663), .A(N5885), .B(N5988));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I999 (.Y(N5868), .A(N5957), .B(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1000 (.Y(N6195), .A(N5840), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1001 (.Y(N6375), .A(N6215), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1002 (.Y(N6550), .A(N6568), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1003 (.Y(N5902), .A(N6106), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1004 (.Y(N6089), .A(N6466), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1005 (.Y(N6280), .A(N6002), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1006 (.Y(N6453), .A(N6365), .B(N5868));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1007 (.Y(N6630), .A(N5885), .B(N5868));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1008 (.Y(N6571), .A(N6653));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1009 (.Y(N5925), .A(N6540));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1010 (.Y(N6245), .A(N6540), .B(N6653));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1011 (.Y(N6470), .A(N6442));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1012 (.Y(N6650), .A(N6159));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1013 (.Y(N6598), .A(N6159), .B(N6442));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1014 (.Y(N6136), .A(N6047), .B(N6511));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1015 (.Y(N5889), .A(N6047));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1016 (.Y(N6072), .A(N6511));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1017 (.Y(N6268), .A(N6406));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1018 (.Y(N6439), .A(N5944));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1019 (.Y(N6490), .A(N5944), .B(N6406));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1020 (.Y(N6027), .A(N6022), .B(N6670));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1021 (.Y(N6507), .A(N6670));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1022 (.Y(N5856), .A(N6022));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1023 (.Y(N6386), .A(N6380), .B(N6200));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1024 (.Y(N6404), .A(N6380));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1025 (.Y(N6590), .A(N6200));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1026 (.Y(N5943), .A(N5905));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1027 (.Y(N6126), .A(N6555));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1028 (.Y(N5916), .A(N5905), .B(N6555));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1029 (.Y(N6665), .A(N6093));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1030 (.Y(N6291), .A(N6284), .B(N6093));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1031 (.Y(N6376), .A(N6284));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1032 (.Y(N6551), .A(N6172));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1033 (.Y(N6643), .A(N6152), .B(N6172));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1034 (.Y(N6281), .A(N6152));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1035 (.Y(N6455), .A(N6503));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1036 (.Y(N6180), .A(N6503), .B(N6523));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1037 (.Y(N6054), .A(N6523));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1038 (.Y(N6533), .A(N6402), .B(N6042));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1039 (.Y(N6600), .A(N6042));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1040 (.Y(N5954), .A(N6402));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1041 (.Y(N6138), .A(N6605));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1042 (.Y(N6326), .A(N6422));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1043 (.Y(N6070), .A(N6605), .B(N6422));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1044 (.Y(N6029), .A(N6496));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1045 (.Y(N6214), .A(N6332));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1046 (.Y(N6432), .A(N6496), .B(N6332));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1047 (.Y(N5920), .A(N6031));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1048 (.Y(N5969), .A(N6031), .B(N5842));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1049 (.Y(N6262), .A(N5842));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1050 (.Y(N6338), .A(N6389), .B(N6217));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1051 (.Y(N5971), .A(N6389));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1052 (.Y(N6151), .A(N6217));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1053 (.Y(N5850), .A(N5923), .B(N6310));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1054 (.Y(N5938), .A(N6310));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1055 (.Y(N6120), .A(N5923));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1056 (.Y(N6225), .A(N6193), .B(N6295));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1057 (.Y(N6660), .A(N6295));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1058 (.Y(N6014), .A(N6193));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1059 (.Y(N6192), .A(N6004));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1060 (.Y(N6372), .A(N6649));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1061 (.Y(N6583), .A(N6004), .B(N6649));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1062 (.Y(N6086), .A(N6185));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1063 (.Y(N6115), .A(N6366), .B(N6185));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1064 (.Y(N6518), .A(N6366));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1065 (.Y(N6476), .A(N5888), .B(N6547));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1066 (.Y(N6244), .A(N5888));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1067 (.Y(N6416), .A(N6547));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1068 (.Y(N6597), .A(N6266));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1069 (.Y(N6208), .A(N6437), .B(N6266));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1070 (.Y(N6383), .A(N6437));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1071 (.Y(N6563), .A(N5974));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1072 (.Y(N5914), .A(N6616));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1073 (.Y(N6370), .A(N5974), .B(N6616));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1074 (.Y(N6461), .A(N6154));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1075 (.Y(N6641), .A(N6343));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1076 (.Y(N5897), .A(N6343), .B(N6154));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1077 (.Y(N6430), .A(N5855));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1078 (.Y(N6275), .A(N5855), .B(N6451));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1079 (.Y(N6147), .A(N6451));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1080 (.Y(N6336), .A(N6403));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1081 (.Y(N6626), .A(N6403), .B(N6233));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1082 (.Y(N6039), .A(N6233));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1083 (.Y(N6164), .A(N6352), .B(N6589));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1084 (.Y(N6580), .A(N6352));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1085 (.Y(N5932), .A(N6589));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1086 (.Y(N6545), .A(N6312), .B(N6124));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1087 (.Y(N5894), .A(N6124));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1088 (.Y(N6080), .A(N6312));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1089 (.Y(N6050), .A(N6663), .B(N6481));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1090 (.Y(N6623), .A(N6663));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1091 (.Y(N5981), .A(N6481));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1092 (.Y(N6162), .A(N6195));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1093 (.Y(N6411), .A(N6375), .B(N6195));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1094 (.Y(N5863), .A(N6375));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1095 (.Y(N6487), .A(N5902), .B(N6550));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1096 (.Y(N6674), .A(N6550));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1097 (.Y(N6024), .A(N5902));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1098 (.Y(N6202), .A(N6280));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1099 (.Y(N6321), .A(N6280), .B(N6089));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1100 (.Y(N5909), .A(N6089));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1101 (.Y(N6096), .A(N6630));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1102 (.Y(N6676), .A(N6630), .B(N6453));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1103 (.Y(N5875), .A(N6453));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1104 (.Y(N6041), .A(N6461), .B(N6597), .C(N6470), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1105 (.Y(N6229), .A(N6192), .B(N6563), .C(N6138), .D(N6202));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1106 (.Y(N6401), .A(N6086), .B(N6551), .C(N6571));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1107 (.Y(N6585), .A(N6401), .B(N6336), .C(N6029), .D(N5920));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1108 (.Y(N5937), .A(N6386), .B(N6050), .C(N6487), .D(N5850));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1109 (.Y(N6119), .A(N6533), .B(N6164), .C(N6136), .D(N6027));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1110 (.Y(N6307), .A(N6225));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1111 (.Y(N6479), .A(N6307), .B(N6041), .C(N6229), .D(N5937));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1114 (.Y(N5987), .A(N6660), .B(N6551));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1115 (.Y(N6449), .A(N6600), .B(N6214), .C(N6162), .D(N6507));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1116 (.Y(N6628), .A(N6268), .B(N6563), .C(N6138), .D(N6650));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1117 (.Y(N6167), .A(N5987), .B(N6202), .C(N6641), .D(N6455));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1118 (.Y(N6517), .A(N6291));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1119 (.Y(N6053), .AN(N6338), .B(N6031), .C(N6449), .D(N6517));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1120 (.Y(N6243), .A(N6487), .B(N5850), .C(N6476), .D(N6545));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1121 (.Y(N6064), .A(N6208));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1122 (.Y(N6255), .A(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1123 (.Y(N5952), .A(N6064), .B(N6255), .C(N6628), .D(N6243));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1125 (.Y(N6562), .A(N5914), .B(N6192), .C(N6404), .D(N6650));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1126 (.Y(N5913), .A(N6623), .B(N6439), .C(N6244), .D(N6321));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1127 (.Y(N6289), .A(N5938), .B(N6338), .C(N6487), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1128 (.Y(N6460), .A(N6411), .B(N6533), .C(N6643), .D(N6027));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1129 (.Y(N6640), .A(N6208), .B(N6180), .C(N6115), .D(N6432));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1130 (.Y(N6425), .A(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1131 (.Y(N6178), .A(N6425), .B(N6562), .C(N5913), .D(N6460));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1134 (.Y(N6611), .A(N6162), .B(N6372), .C(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1135 (.Y(N6146), .A(N6563), .B(N6138), .C(N6623), .D(N6202));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1136 (.Y(N6335), .A(N6096), .B(N6430), .C(N5971), .D(N6641));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1137 (.Y(N6500), .A(N6244), .B(N5954), .C(N6281), .D(N5889));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1138 (.Y(N5847), .A(N6014), .B(N6518), .C(N6336), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1139 (.Y(N6038), .A(N6386), .B(N6487), .C(N6545), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1140 (.Y(N6222), .A(N6611), .B(N6335), .C(N5847), .D(N6500));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1143 (.Y(N6544), .A(N6597), .B(N6262), .C(N5981), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1144 (.Y(N5893), .A(N6563), .B(N5943), .C(N5954), .D(N6336));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1145 (.Y(N6079), .A(N6072), .B(N6151), .C(N6507));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1146 (.Y(N6272), .A(N6079), .B(N5850), .C(N6490), .D(N5897));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1147 (.Y(N6606), .A(N6432));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1149 (.Y(N6409), .A(N5894), .B(N6126));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1150 (.Y(N6239), .A(N6507), .B(N5981), .C(N5914), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1151 (.Y(N6592), .A(N6665), .B(N6409), .C(N6192), .D(N6641));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1152 (.Y(N5947), .A(N5863), .B(N6580), .C(N5889), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1153 (.Y(N6133), .A(N6676), .B(N6338), .C(N6476), .D(N6643));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1154 (.Y(N5961), .A(N6180));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1155 (.Y(N6486), .A(N5961), .B(N6239), .C(N5947), .D(N6592));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1156 (.Y(N6672), .A(N6133));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1158 (.Y(N5908), .A(N6072), .B(N5894), .C(N6162), .D(N6151));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1159 (.Y(N6636), .A(N6200), .B(N6547), .C(N6649), .D(N6653));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1160 (.Y(N5995), .A(N5914), .B(N6650), .C(N6096), .D(N6430));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1161 (.Y(N6175), .A(N6024), .B(N6120), .C(N6641), .D(N5954));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1162 (.Y(N6359), .A(N6014), .B(N6383), .C(N6336), .D(N5920));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1163 (.Y(N6527), .A(N5916), .B(N6291), .C(N6490), .D(N6643));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1164 (.Y(N5874), .A(N5908));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1165 (.Y(N6062), .A(N5995));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1166 (.Y(N6254), .A(N6180), .B(N5874), .C(N6062), .D(N6636));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1168 (.Y(N5843), .A(N6674), .B(N6563), .C(N6376), .D(N6641));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1169 (.Y(N6034), .A(N5889), .B(N6583), .C(N6386), .D(N5916));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1170 (.Y(N6219), .A(N6571), .B(N6262), .C(N6470));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1171 (.Y(N6392), .A(N6676), .B(N6275), .C(N6219), .D(N6338));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1172 (.Y(N6573), .A(N5850), .B(N6476), .C(N6545), .D(N6643));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1173 (.Y(N5928), .A(N6027), .B(N6225), .C(N6180), .D(N6115));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1174 (.Y(N6298), .A(N6606), .B(N6034), .C(N5843), .D(N5928));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1177 (.Y(N5978), .A(N6072), .B(N6162));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1178 (.Y(N6075), .A(N6597), .B(N6326), .C(N6470), .D(N6372));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1179 (.Y(N6269), .A(N5914), .B(N6674), .C(N5925), .D(N5943));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1180 (.Y(N6441), .A(N6202), .B(N6430), .C(N6641), .D(N5856));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1181 (.Y(N6619), .A(N6014), .B(N6518), .C(N6336), .D(N6050));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1182 (.Y(N6157), .A(N6676), .B(N6291), .C(N5978), .D(N6338));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1183 (.Y(N6345), .A(N5850), .B(N6476), .C(N6545), .D(N6533));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1184 (.Y(N5858), .A(N5961), .B(N6075), .C(N6269), .D(N6619));
NOR4BX1 inst_cellmath__203_0_I23855 (.Y(N9277), .AN(N5858), .B(N6441), .C(N6345), .D(N6157));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1189 (.Y(N6128), .A(N6660), .B(N6214), .C(N6162), .D(N6054));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1190 (.Y(N6315), .A(N6147), .B(N6470), .C(N6372), .D(N5938));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1191 (.Y(N6484), .A(N5914), .B(N6376), .C(N5971), .D(N6439));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1192 (.Y(N6668), .A(N6244), .B(N5889), .C(N5856), .D(N6383));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1193 (.Y(N6020), .A(N6518), .B(N5920), .C(N6386), .D(N6245));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1194 (.Y(N6199), .A(N6070), .B(N5916), .C(N6487), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1195 (.Y(N6378), .A(N6545), .B(N6164), .C(N6643), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1196 (.Y(N6554), .A(N6128), .B(N6315), .C(N6484), .D(N6668));
NOR4BX1 inst_cellmath__203_0_I23856 (.Y(N9670), .AN(N6554), .B(N6020), .C(N6378), .D(N6199));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1201 (.Y(N6522), .A(N5981), .B(N6665), .C(N6461), .D(N6192));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1202 (.Y(N5870), .A(N6404), .B(N5943), .C(N6650), .D(N6202));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1203 (.Y(N6058), .A(N6096), .B(N6244), .C(N5863), .D(N5954));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1204 (.Y(N6250), .A(N6580), .B(N6014), .C(N6383), .D(N6455));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1205 (.Y(N6420), .A(N6518), .B(N6029), .C(N5920), .D(N6370));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1206 (.Y(N6603), .A(N6275), .B(N6338), .C(N6545), .D(N6136));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1207 (.Y(N5956), .A(N6027));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1208 (.Y(N6140), .A(N5956), .B(N6522), .C(N5870), .D(N6058));
NOR4BX1 inst_cellmath__203_0_I23857 (.Y(N10038), .AN(N6140), .B(N6250), .C(N6603), .D(N6420));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1213 (.Y(N5922), .A(N6660), .B(N6126), .C(N6039), .D(N6507));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1214 (.Y(N6107), .A(N6326), .B(N6590), .C(N6470), .D(N5925));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1215 (.Y(N6293), .A(N6024), .B(N6120), .C(N6439), .D(N6641));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1216 (.Y(N6468), .A(N6244), .B(N5863), .C(N5889), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1217 (.Y(N6647), .A(N5920), .B(N6583), .C(N6370), .D(N6050));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1218 (.Y(N6003), .A(N6676), .B(N6275), .C(N6291), .D(N6545));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1219 (.Y(N6184), .A(N6533), .B(N6164), .C(N6208), .D(N6180));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1220 (.Y(N6142), .A(N6115));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1221 (.Y(N6536), .A(N6142), .B(N5922), .C(N6107), .D(N6468));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1222 (.Y(N5887), .A(N6293), .B(N6647), .C(N6184), .D(N6003));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1224 (.Y(N5853), .A(N6072), .B(N5894));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1225 (.Y(N6153), .A(N6151), .B(N5932), .C(N6590), .D(N6416));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1226 (.Y(N6342), .A(N5981), .B(N6665), .C(N6192), .D(N6563));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1227 (.Y(N6505), .A(N5925), .B(N6650), .C(N6383), .D(N6455));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1228 (.Y(N6043), .A(N5853), .B(N5920), .C(N6321), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1229 (.Y(N6232), .A(N5850), .B(N6411), .C(N6643), .D(N6225));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1230 (.Y(N6587), .A(N6606), .B(N6153), .C(N6505), .D(N6342));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1233 (.Y(N6016), .A(N6039), .B(N6072), .C(N5894));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1234 (.Y(N6373), .A(N6126), .B(N6461), .C(N6597), .D(N6054));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1235 (.Y(N6548), .A(N6147), .B(N6470), .C(N6563), .D(N5925));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1236 (.Y(N5901), .A(N6138), .B(N6623), .C(N6376), .D(N6120));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1237 (.Y(N5990), .A(N5920), .B(N6338), .C(N6490), .D(N6476));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1238 (.Y(N6169), .A(N6373));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1239 (.Y(N6353), .A(N6411), .B(N6169), .C(N6643), .D(N6027));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1240 (.Y(N6247), .A(N6352), .B(N6402), .C(N6193), .D(N6016));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1241 (.Y(N6418), .A(N5901), .B(N6548), .C(N6606), .D(N6142));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1243 (.Y(N6492), .A(N6571), .B(N5909), .C(N6214), .D(N6126));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1244 (.Y(N5838), .A(N6151), .B(N5932), .C(N6326), .D(N5875));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1245 (.Y(N6028), .A(N5914), .B(N6674), .C(N6404), .D(N6623));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1246 (.Y(N6212), .A(N6439), .B(N5863), .C(N5954), .D(N5856));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1247 (.Y(N6387), .A(N6492));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1248 (.Y(N6566), .A(N6583), .B(N6275), .C(N6387), .D(N5850));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1249 (.Y(N5918), .A(N5838));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1250 (.Y(N6102), .A(N6476), .B(N5918), .C(N6545), .D(N6136));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1251 (.Y(N6000), .A(N6028), .B(N6212), .C(N6064), .D(N6142));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1253 (.Y(N5970), .A(N5981), .B(N6376), .C(N5971), .D(N5863));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1254 (.Y(N6149), .A(N6281), .B(N5856), .C(N6455), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1255 (.Y(N6339), .A(N5916), .B(N6676), .C(N6275), .D(N6487));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1256 (.Y(N6502), .A(N6326), .B(N6268), .C(N6590));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1257 (.Y(N5851), .A(N5850), .B(N6502), .C(N6545), .D(N6136));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1258 (.Y(N6227), .A(N6255), .B(N5970), .C(N6149), .D(N6339));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1260 (.Y(N6117), .A(N6660), .B(N6086), .C(N5894), .D(N6214));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1261 (.Y(N6305), .A(N6507), .B(N6461), .C(N6597), .D(N5875));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1262 (.Y(N6477), .A(N6054), .B(N6416), .C(N5981), .D(N6372));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1263 (.Y(N6659), .A(N5914), .B(N6665), .C(N6202), .D(N6430));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1264 (.Y(N6012), .A(N5971), .B(N6024), .C(N6120), .D(N5954));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1265 (.Y(N5898), .A(N6352), .B(N6152), .C(N6403), .D(N6117));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1266 (.Y(N6084), .A(N5920), .B(N5916), .C(N6490), .D(N6411));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1267 (.Y(N6276), .A(N6136));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1268 (.Y(N6448), .A(N6276), .B(N6305), .C(N6477), .D(N6659));
NOR4BBX1 inst_cellmath__203_0_I23851 (.Y(N8842), .AN(N5898), .BN(N6448), .C(N6012), .D(N6084));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1272 (.Y(N6414), .A(N6551), .B(N6151), .C(N6039), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1273 (.Y(N6595), .A(N6202), .B(N6430), .C(N6120), .D(N5863));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1274 (.Y(N5951), .A(N5954), .B(N6580), .C(N5920), .D(N6245));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1275 (.Y(N6135), .A(N6070), .B(N5916), .C(N6598), .D(N6050));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1276 (.Y(N6322), .A(N6291), .B(N5897), .C(N6225), .D(N6208));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1277 (.Y(N6678), .A(N6142), .B(N6414), .C(N6322), .D(N6595));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1280 (.Y(N5878), .A(N5863), .B(N6580), .C(N5920), .D(N5916));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1281 (.Y(N6066), .A(N6291), .B(N6338), .C(N6487), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1282 (.Y(N6257), .A(N6476), .B(N6545), .C(N6643), .D(N6180));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1283 (.Y(N6610), .A(N6089), .B(N6042), .C(N6451), .D(N6310));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1284 (.Y(N5964), .A(N6142), .B(N6610), .C(N6066), .D(N5878));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1286 (.Y(N6396), .A(N6162), .B(N6262), .C(N6580), .D(N6370));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1287 (.Y(N6576), .A(N6070), .B(N5916), .C(N6050), .D(N6291));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1288 (.Y(N5931), .A(N6476), .B(N6545), .C(N6533), .D(N6643));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1290 (.Y(N6542), .A(N5932), .B(N6386));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1291 (.Y(N6078), .A(N6370), .B(N6245), .C(N6598), .D(N6275));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1292 (.Y(N6270), .A(N6490), .B(N5897), .C(N6476), .D(N6136));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1293 (.Y(N6443), .A(N6027), .B(N6208), .C(N6115), .D(N6626));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1295 (.Y(N5861), .A(N6583), .B(N6386));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1296 (.Y(N6237), .A(N6245), .B(N6070), .C(N5916), .D(N6598));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1297 (.Y(N6407), .A(N6291), .B(N6338), .C(N5850), .D(N6490));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1298 (.Y(N6591), .A(N6533), .B(N6643), .C(N6136), .D(N6027));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1299 (.Y(N5945), .A(N6225), .B(N6180), .C(N6432), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1300 (.Y(N6131), .A(N5861), .B(N6237), .C(N6407), .D(N5945));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1302 (.Y(N5993), .A(N6086), .B(N6551), .C(N6126), .D(N6597));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1303 (.Y(N6173), .A(N6268), .B(N6372), .C(N5914), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1304 (.Y(N6358), .A(N6665), .B(N6430), .C(N6120), .D(N6244));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1305 (.Y(N6524), .A(N5954), .B(N5856), .C(N6336), .D(N6029));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1306 (.Y(N5873), .A(N5993));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1307 (.Y(N6061), .A(N5873), .B(N5920), .C(N6070), .D(N6050));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1308 (.Y(N6252), .A(N6676), .B(N6338), .C(N5897), .D(N6545));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1309 (.Y(N6424), .A(N6164));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1310 (.Y(N5958), .A(N6173), .B(N6358), .C(N6524), .D(N6424));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1312 (.Y(N5926), .A(N6039), .B(N6600));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1313 (.Y(N6572), .A(N6162), .B(N6507), .C(N6461), .D(N6147));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1314 (.Y(N6110), .A(N6416), .B(N5938), .C(N5926), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1315 (.Y(N6296), .A(N6665), .B(N5925), .C(N6623), .D(N6096));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1316 (.Y(N6471), .A(N6080), .B(N6014), .C(N6518), .D(N6386));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1317 (.Y(N6651), .A(N6370), .B(N5916), .C(N6598), .D(N6180));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1318 (.Y(N6186), .A(N6606), .B(N6572), .C(N6110), .D(N6471));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1321 (.Y(N5976), .A(N6072), .B(N6600), .C(N5894));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1322 (.Y(N6344), .A(N6214), .B(N6262), .C(N6590), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1323 (.Y(N6508), .A(N6138), .B(N5971), .C(N6244), .D(N6580));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1324 (.Y(N5857), .A(N6014), .B(N6383), .C(N6455), .D(N6321));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1325 (.Y(N6045), .A(N6291), .B(N5897), .C(N6027), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1326 (.Y(N6234), .A(N5976), .B(N6344), .C(N6508), .D(N5857));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1328 (.Y(N6314), .A(N5894), .B(N6151));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1329 (.Y(N6666), .A(N5875), .B(N6054), .C(N6416), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1330 (.Y(N6019), .A(N6138), .B(N6650), .C(N6623), .D(N6120));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1331 (.Y(N6196), .A(N6439), .B(N5863), .C(N6580), .D(N5889));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1332 (.Y(N6377), .A(N6014), .B(N6518), .C(N6583), .D(N6386));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1333 (.Y(N6553), .A(N6314));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1334 (.Y(N5903), .A(N6487), .B(N6553), .C(N6643), .D(N6432));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1335 (.Y(N6282), .A(N6425), .B(N6019), .C(N6666), .D(N6377));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1338 (.Y(N6056), .A(N5909), .B(N6214), .C(N6326), .D(N5914));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1339 (.Y(N6419), .A(N6600), .B(N6674), .C(N6376), .D(N5971));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1340 (.Y(N6601), .A(N6120), .B(N6244), .C(N6281), .D(N5889));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1341 (.Y(N5955), .A(N6014), .B(N6383), .C(N6518), .D(N6336));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1342 (.Y(N6139), .A(N6583), .B(N5916), .C(N6598), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1343 (.Y(N6328), .A(N6545), .B(N6411), .C(N6164), .D(N6027));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1344 (.Y(N6030), .A(N6419), .B(N6056), .C(N6601), .D(N6425));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1346 (.Y(N6105), .A(N6660), .B(N6600));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1347 (.Y(N6465), .A(N6126), .B(N6268), .C(N6147), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1348 (.Y(N6646), .A(N6138), .B(N6650), .C(N6623), .D(N6641));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1349 (.Y(N6535), .A(N6375), .B(N6047), .C(N6503), .D(N6105));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1350 (.Y(N5884), .A(N6336), .B(N6029), .C(N5920), .D(N6583));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1351 (.Y(N6071), .A(N6321), .B(N5850), .C(N6027), .D(N6208));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1352 (.Y(N6435), .A(N6142), .B(N6646), .C(N6465), .D(N6071));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1354 (.Y(N6230), .A(N6126), .B(N6416), .C(N5981), .D(N6404));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1355 (.Y(N6586), .A(N6086), .B(N6376), .C(N5863), .D(N5954));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1356 (.Y(N5940), .A(N6281), .B(N5889), .C(N6014), .D(N6383));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1357 (.Y(N6121), .A(N6029), .B(N6275), .C(N6338), .D(N6487));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1358 (.Y(N6309), .A(N5850), .B(N5897), .C(N6545), .D(N6164));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1359 (.Y(N6661), .A(N5961), .B(N6230), .C(N6586), .D(N5940));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1362 (.Y(N6279), .A(N5909), .B(N6126), .C(N6507));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1363 (.Y(N6629), .A(N5932), .B(N6326), .C(N6054), .D(N5981));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1364 (.Y(N5989), .A(N6192), .B(N6563), .C(N6096), .D(N6024));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1365 (.Y(N6168), .A(N6244), .B(N6080), .C(N6383), .D(N6336));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1366 (.Y(N6351), .A(N6275), .B(N6291), .C(N6490), .D(N6533));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1367 (.Y(N6519), .A(N6643), .B(N6136), .C(N6225), .D(N6432));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1368 (.Y(N5867), .A(N6279), .B(N6629), .C(N5989), .D(N6168));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1371 (.Y(N6324), .A(N6660), .B(N5894), .C(N6151), .D(N6054));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1372 (.Y(N6491), .A(N5981), .B(N6372), .C(N5914), .D(N6430));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1373 (.Y(N5837), .A(N6120), .B(N6439), .C(N5863), .D(N6580));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1374 (.Y(N6026), .A(N6281), .B(N6336), .C(N6029), .D(N5920));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1375 (.Y(N6211), .A(N6245), .B(N6598), .C(N6676), .D(N6291));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1376 (.Y(N6385), .A(N5897), .B(N6533), .C(N6136), .D(N6115));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1377 (.Y(N6565), .A(N6324), .B(N6491), .C(N5837), .D(N6211));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1380 (.Y(N6181), .A(N6660), .B(N6086), .C(N6597), .D(N6262));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1381 (.Y(N6364), .A(N5875), .B(N6268), .C(N6054), .D(N6147));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1382 (.Y(N6532), .A(N6665), .B(N6563), .C(N5925), .D(N5943));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1383 (.Y(N5881), .A(N6650), .B(N5971), .C(N6120), .D(N5954));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1384 (.Y(N6069), .A(N6281), .B(N5889), .C(N6583), .D(N6070));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1385 (.Y(N6260), .A(N6321), .B(N6164), .C(N6626), .D(N6432));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1386 (.Y(N6433), .A(N6181), .B(N6364), .C(N6069), .D(N5881));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1389 (.Y(N6040), .A(N6551), .B(N6162), .C(N6126), .D(N6507));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1390 (.Y(N6226), .A(N6461), .B(N6268), .C(N6590), .D(N5981));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1391 (.Y(N6399), .A(N6138), .B(N6202), .C(N6244), .D(N6580));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1392 (.Y(N6582), .A(N6455), .B(N6518), .C(N6029), .D(N6598));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1393 (.Y(N5935), .A(N6275), .B(N6291), .C(N6338), .D(N6545));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1394 (.Y(N6114), .A(N6533), .B(N6225), .C(N6626), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1395 (.Y(N6304), .A(N6040), .B(N6226), .C(N6399), .D(N6582));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1398 (.Y(N6165), .A(N6660), .B(N6086));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1399 (.Y(N6082), .A(N6551), .B(N6600), .C(N5909), .D(N6214));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1400 (.Y(N6274), .A(N6162), .B(N6461), .C(N5932), .D(N6268));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1401 (.Y(N6446), .A(N6590), .B(N6054), .C(N6372), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1402 (.Y(N6625), .A(N6665), .B(N6138), .C(N5943), .D(N6623));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1403 (.Y(N5984), .A(N6430), .B(N6244), .C(N5856), .D(N6336));
NAND3XL hyperpropagate_4_1_A_I23860 (.Y(N37704), .A(N6370), .B(N6165), .C(N5850));
NOR2XL hyperpropagate_4_1_A_I23861 (.Y(N5950), .A(N6082), .B(N37704));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1406 (.Y(N6241), .A(N6276), .B(N6064), .C(N6274), .D(N6446));
NOR4BBX1 inst_cellmath__203_0_I23852 (.Y(N9284), .AN(N5950), .BN(N6241), .C(N6625), .D(N5984));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1411 (.Y(N5911), .A(N6551), .B(N6600));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1412 (.Y(N6206), .A(N6461), .B(N6590), .C(N6623), .D(N6376));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1413 (.Y(N6382), .A(N5971), .B(N6120), .C(N6439), .D(N6244));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1414 (.Y(N6560), .A(N6080), .B(N6580), .C(N6455), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1415 (.Y(N6098), .A(N5911), .B(N5920), .C(N6583), .D(N6370));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1416 (.Y(N6287), .A(N6070), .B(N6487), .C(N6027), .D(N6208));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1417 (.Y(N6638), .A(N6255), .B(N6206), .C(N6382), .D(N6560));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1420 (.Y(N6428), .A(N6600), .B(N6597), .C(N5932), .D(N6590));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1421 (.Y(N6608), .A(N5981), .B(N5914), .C(N6192), .D(N6430));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1422 (.Y(N5963), .A(N6080), .B(N6281), .C(N6518), .D(N6336));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1423 (.Y(N6144), .A(N6245), .B(N6598), .C(N6321), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1424 (.Y(N6498), .A(N6660), .B(N6338), .C(N6487), .D(N6490));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1425 (.Y(N5845), .A(N5897), .B(N6136), .C(N6027), .D(N6180));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1426 (.Y(N6220), .A(N6606), .B(N6428), .C(N6608), .D(N6144));
NOR4BX1 inst_cellmath__203_0_I23858 (.Y(N10044), .AN(N6220), .B(N5963), .C(N6498), .D(N5845));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1431 (.Y(N6007), .A(N6039), .B(N6086), .C(N6072), .D(N6214));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1432 (.Y(N6188), .A(N6507), .B(N6326), .C(N6268), .D(N6470));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1433 (.Y(N6541), .A(N5938), .B(N6571), .C(N6192), .D(N5943));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1434 (.Y(N5892), .A(N6430), .B(N6376), .C(N5971), .D(N6244));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1435 (.Y(N5979), .A(N5920), .B(N6386), .C(N6370), .D(N6050));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1436 (.Y(N6512), .AN(N6411), .B(N6188), .C(N6307), .D(N6541));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1437 (.Y(N5860), .A(N6312), .B(N6152), .C(N6503), .D(N6007));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1438 (.Y(N6236), .AN(N6512), .B(N5892), .C(N5979), .D(N5860));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1440 (.Y(N6671), .A(N6054), .B(N6372), .C(N6665), .D(N5943));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1441 (.Y(N6556), .A(N5855), .B(N5888), .C(N6152), .D(N6314));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1442 (.Y(N5906), .A(N5920), .B(N6245), .C(N6070), .D(N6164));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1443 (.Y(N6094), .A(N6136), .B(N6027), .C(N6225), .D(N6208));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1444 (.Y(N6457), .A(N6255), .B(N6671), .C(N6094), .D(N5906));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1446 (.Y(N5872), .A(N6126), .B(N6147), .C(N6244), .D(N6281));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1447 (.Y(N6060), .A(N5920), .B(N6386), .C(N6370), .D(N6245));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1448 (.Y(N6251), .A(N6598), .B(N6338), .C(N5850), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1449 (.Y(N6423), .A(N6533), .B(N6027), .C(N6208), .D(N6180));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1451 (.Y(N6497), .A(N6262), .B(N6244), .C(N6281));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1452 (.Y(N6032), .A(N6370), .B(N6245), .C(N6070), .D(N6598));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1453 (.Y(N6218), .A(N6050), .B(N6321), .C(N6676), .D(N6275));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1454 (.Y(N6390), .A(N6487), .B(N6490), .C(N5897), .D(N6545));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1455 (.Y(N6570), .A(N6411), .B(N6533), .C(N6164), .D(N6136));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1456 (.Y(N5924), .A(N6208), .B(N6180), .C(N6626), .D(N6432));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1457 (.Y(N6109), .A(N6032), .B(N6218), .C(N6570), .D(N6497));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1460 (.Y(N6537), .A(N6551), .B(N6244));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1461 (.Y(N6073), .A(N6386), .B(N6370), .C(N6245), .D(N5916));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1462 (.Y(N6267), .A(N6598), .B(N6050), .C(N6321), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1463 (.Y(N6438), .A(N6275), .B(N6291), .C(N6487), .D(N6490));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1464 (.Y(N6617), .A(N5897), .B(N6545), .C(N6411), .D(N6164));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1465 (.Y(N5975), .A(N6136), .B(N6027), .C(N6208), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1466 (.Y(N6155), .A(N6073), .B(N6267), .C(N6438), .D(N6537));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1469 (.Y(N5942), .A(N6416), .B(N6583), .C(N6386), .D(N6245));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1470 (.Y(N6125), .A(N6070), .B(N5916), .C(N6598), .D(N6291));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1471 (.Y(N6313), .A(N6338), .B(N5850), .C(N6490), .D(N6533));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1472 (.Y(N6482), .A(N6643), .B(N6136), .C(N6027), .D(N6225));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1473 (.Y(N6664), .A(N6180), .B(N6115), .C(N6432), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1474 (.Y(N6017), .A(N5942), .B(N6125), .C(N6313), .D(N6664));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1476 (.Y(N6090), .A(N6162), .B(N6126), .C(N6461));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1477 (.Y(N6454), .A(N6326), .B(N5981), .C(N5938), .D(N6404));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1478 (.Y(N6631), .A(N6563), .B(N5925), .C(N6096), .D(N6580));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1479 (.Y(N5992), .A(N6281), .B(N5889), .C(N5920), .D(N6583));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1480 (.Y(N6170), .A(N6598), .B(N6321), .C(N6291), .D(N6338));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1481 (.Y(N6354), .A(N6487), .B(N6490), .C(N6533), .D(N6027));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1482 (.Y(N6520), .A(N6090), .B(N6454), .C(N6631), .D(N6170));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1483 (.Y(N6055), .A(N5992));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1484 (.Y(inst_cellmath__195[0]), .AN(N6354), .B(N6055), .C(N6520));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1485 (.Y(N6327), .A(N6214), .B(N6151), .C(N6326), .D(N5914));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1486 (.Y(N6494), .A(N5925), .B(N6202), .C(N6439), .D(N6281));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1487 (.Y(N5839), .A(N6383), .B(N6518), .C(N6583), .D(N6386));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1488 (.Y(N6213), .A(N6598));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1489 (.Y(N6388), .A(N6050));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1490 (.Y(N6567), .AN(N5916), .B(N6388), .C(N6124), .D(N6213));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1491 (.Y(N5919), .A(N6487), .B(N6476), .C(N6411), .D(N6533));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1492 (.Y(N6104), .A(N6164), .B(N6136), .C(N6027), .D(N6225));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1493 (.Y(N6464), .A(N6425), .B(N6327), .C(N5839), .D(N6494));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1494 (.Y(N6645), .A(N5919));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1495 (.Y(N6001), .A(N6104));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1496 (.Y(inst_cellmath__195[1]), .A(N6645), .B(N6567), .C(N6001), .D(N6464));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1497 (.Y(N5883), .A(N6551), .B(N6162), .C(N6470));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1498 (.Y(N6263), .A(N6665), .B(N5925), .C(N6096), .D(N6439));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1499 (.Y(N6434), .A(N5954), .B(N5889), .C(N6014), .D(N6455));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1500 (.Y(N6613), .A(N6029), .B(N5920), .C(N6583), .D(N6386));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1501 (.Y(N5972), .A(N6370), .B(N6050), .C(N6338), .D(N5850));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1502 (.Y(N6150), .A(N6476), .B(N6164), .C(N6208), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1503 (.Y(N6341), .A(N5883), .B(N6434), .C(N6263), .D(N6150));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1504 (.Y(N5852), .A(N6613));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1505 (.Y(inst_cellmath__195[2]), .AN(N5972), .B(N5852), .C(N6341));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1506 (.Y(N6118), .A(N6470), .B(N5981), .C(N6665), .D(N6192));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1507 (.Y(N6308), .A(N5925), .B(N6096), .C(N6024), .D(N6080));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1508 (.Y(N6480), .A(N5863), .B(N5954), .C(N6281), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1509 (.Y(N6015), .A(N6416), .B(N6386), .C(N6370), .D(N6070));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1510 (.Y(N6191), .A(N6321), .B(N6275), .C(N5850), .D(N6490));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1511 (.Y(N6371), .A(N5897), .B(N6225), .C(N6208), .D(N6180));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1512 (.Y(N5899), .A(N6142), .B(N6308), .C(N6118), .D(N6480));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1513 (.Y(N6085), .A(N6015));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1514 (.Y(N6278), .A(N6191));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1515 (.Y(N6450), .A(N6371));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1516 (.Y(inst_cellmath__195[3]), .A(N6085), .B(N6278), .C(N6450), .D(N5899));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1517 (.Y(N5866), .A(N6072), .B(N6600), .C(N5894), .D(N5909));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1518 (.Y(N6052), .A(N6214), .B(N6151), .C(N6326), .D(N6268));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1519 (.Y(N6415), .A(N5938), .B(N6571), .C(N6192), .D(N6404));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1520 (.Y(N6596), .A(N6623), .B(N6024), .C(N6014), .D(N6291));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1521 (.Y(N6323), .AN(N6476), .B(N6052), .C(N6424), .D(N5866));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1522 (.Y(N6209), .A(N5956), .B(N6064), .C(N5961), .D(N6415));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1523 (.Y(inst_cellmath__195[4]), .AN(N6596), .B(N6323), .C(N6209));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1524 (.Y(N5998), .A(N6214), .B(N5938), .C(N6404), .D(N5925));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1525 (.Y(N6362), .A(N6376), .B(N6439), .C(N5909), .D(N6244));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1526 (.Y(N6530), .A(N5856), .B(N6518), .C(N6050), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1527 (.Y(N5879), .A(N6275), .B(N6338), .C(N6487), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1528 (.Y(N6067), .A(N6643), .B(N6136), .C(N6225), .D(N6208));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1529 (.Y(N6429), .A(N6425), .B(N5998), .C(N6530), .D(N6362));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1530 (.Y(N5966), .A(N5879));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1531 (.Y(inst_cellmath__195[5]), .AN(N6067), .B(N5966), .C(N6429));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1532 (.Y(N5848), .A(N6551), .B(N6600), .C(N6262), .D(N5875));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1533 (.Y(N6037), .A(N6416), .B(N6470), .C(N6372), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1534 (.Y(N6223), .A(N6138), .B(N6080), .C(N6580), .D(N5856));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1535 (.Y(N6397), .A(N6383), .B(N6029), .C(N6370), .D(N5916));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1536 (.Y(N6578), .A(N6050), .B(N6321), .C(N6275), .D(N6487));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1537 (.Y(N5933), .A(N5850), .B(N6490), .C(N5897), .D(N6411));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1538 (.Y(N6112), .A(N6136), .B(N6180), .C(N6115), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1539 (.Y(N6302), .A(N5848), .B(N6223), .C(N6037), .D(N6397));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1540 (.Y(N6474), .A(N6578));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1541 (.Y(N6655), .A(N5933));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1542 (.Y(N6010), .A(N6112));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1543 (.Y(inst_cellmath__195[6]), .A(N6474), .B(N6655), .C(N6010), .D(N6302));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1544 (.Y(N5895), .A(N5894), .B(N6126), .C(N5932));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1545 (.Y(N6271), .A(N5875), .B(N6054), .C(N6416), .D(N6470));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1546 (.Y(N6444), .A(N5981), .B(N6372), .C(N5914), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1547 (.Y(N6622), .A(N6439), .B(N6641), .C(N5856), .D(N6518));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1548 (.Y(N5982), .A(N5920), .B(N6245), .C(N6070), .D(N6321));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1549 (.Y(N6161), .A(N6275), .B(N6487), .C(N6225), .D(N6626));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1550 (.Y(N6514), .A(N5895), .B(N6271), .C(N6622), .D(N6444));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1551 (.Y(inst_cellmath__195[7]), .A(N6514), .B(N5982), .C(N6161));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1552 (.Y(N5948), .A(N6072), .B(N5909), .C(N6214));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1553 (.Y(N6319), .A(N6162), .B(N6597), .C(N6262), .D(N5875));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1554 (.Y(N6488), .A(N6268), .B(N6416), .C(N6470), .D(N5981));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1555 (.Y(N6673), .A(N6372), .B(N5938), .C(N6024), .D(N6641));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1556 (.Y(N6023), .A(N6580), .B(N5856), .C(N6291), .D(N6338));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1557 (.Y(N6203), .A(N6545), .B(N6533), .C(N6180), .D(N6115));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1558 (.Y(N6558), .A(N5948), .B(N6319), .C(N6673), .D(N6488));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1559 (.Y(inst_cellmath__195[8]), .A(N6558), .B(N6023), .C(N6203));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1560 (.Y(N6526), .A(N6268), .B(N6138), .C(N5943), .D(N6202));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1561 (.Y(N5876), .A(N6580), .B(N5856), .C(N6014), .D(N6383));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1562 (.Y(N6063), .A(N6461), .B(N6551), .C(N6571));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1563 (.Y(N6253), .A(N6455), .B(N6063), .C(N5920), .D(N6275));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1564 (.Y(N6426), .A(N6487), .B(N5850), .C(N6476), .D(N6411));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1565 (.Y(N5960), .A(N6606), .B(N6526), .C(N5876), .D(N6253));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1566 (.Y(inst_cellmath__195[9]), .AN(N6426), .B(N5960));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1567 (.Y(N6393), .A(N6461), .B(N6147), .C(N6416), .D(N5981));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1568 (.Y(N5929), .A(N5938), .B(N5914), .C(N5909), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1569 (.Y(N6111), .A(N6404), .B(N5971), .C(N6439), .D(N5856));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1570 (.Y(N6297), .A(N6014), .B(N6455), .C(N6518), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1571 (.Y(N6472), .A(N6245), .B(N6598), .C(N6676), .D(N6164));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1572 (.Y(N6005), .A(N6255), .B(N6111), .C(N6393), .D(N6297));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1573 (.Y(N6367), .A(N6472));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1574 (.Y(inst_cellmath__195[10]), .AN(N5929), .B(N6367), .C(N6005));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1575 (.Y(N6620), .A(N6151), .B(N6590), .C(N6054), .D(N6147));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1576 (.Y(N5977), .A(N6470), .B(N6372), .C(N6563), .D(N6138));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1577 (.Y(N6158), .A(N6202), .B(N6024), .C(N5889), .D(N6336));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1578 (.Y(N6346), .A(N6245), .B(N6291), .C(N6490), .D(N6533));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1579 (.Y(N6510), .A(N6643), .B(N6225), .C(N6208), .D(N6115));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1580 (.Y(N5859), .A(N6620), .B(N5977), .C(N6158), .D(N6346));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1581 (.Y(inst_cellmath__195[11]), .AN(N6510), .B(N5859));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1582 (.Y(N6129), .A(N6126), .B(N6507), .C(N6461), .D(N6268));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1583 (.Y(N6316), .A(N6590), .B(N6372), .C(N5914), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1584 (.Y(N6669), .A(N5909), .B(N6665), .C(N6138), .D(N6650));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1585 (.Y(N6021), .A(N6244), .B(N5889), .C(N6455), .D(N6336));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1586 (.Y(N6198), .A(N5850), .B(N6545), .C(N6411), .D(N6533));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1587 (.Y(N6379), .A(N6164), .B(N6208), .C(N6115), .D(N6432));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1588 (.Y(N6092), .A(N6129), .B(N6669), .C(N6316), .D(N6425));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1589 (.Y(inst_cellmath__195[12]), .A(N6021), .B(N6092), .C(N6379), .D(N6198));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1590 (.Y(N6356), .A(N6551), .B(N6597), .C(N6326), .D(N5875));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1591 (.Y(N5871), .A(N6039), .B(N6590), .C(N5981), .D(N5943));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1592 (.Y(N6059), .A(N6202), .B(N6641), .C(N5954), .D(N6580));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1593 (.Y(N6249), .A(N5856), .B(N6455), .C(N6518), .D(N6598));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1594 (.Y(N6421), .A(N6291), .B(N6487), .C(N5850), .D(N6490));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1595 (.Y(N6604), .A(N6545), .B(N6411), .C(N6136), .D(N6432));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1596 (.Y(N6331), .A(N6356), .B(N5871), .C(N6059), .D(N6425));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1597 (.Y(inst_cellmath__195[13]), .A(N6331), .B(N6249), .C(N6421), .D(N6604));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1598 (.Y(N6216), .A(N6214), .B(N6507));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1599 (.Y(N6569), .A(N6597), .B(N6326), .C(N6372), .D(N5938));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1600 (.Y(N5921), .A(N5914), .B(N6674), .C(N6665), .D(N6404));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1601 (.Y(N6108), .A(N5943), .B(N6623), .C(N6439), .D(N6641));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1602 (.Y(N6294), .A(N6080), .B(N5863), .C(N5954), .D(N6281));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1603 (.Y(N6467), .A(N6014), .B(N6518), .C(N6336), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1604 (.Y(N6648), .A(N6275), .B(N6164), .C(N6136), .D(N6180));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1605 (.Y(N6183), .A(N6216), .B(N6108), .C(N6569), .D(N6294));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1606 (.Y(inst_cellmath__195[14]), .A(N5921), .B(N6183), .C(N6467), .D(N6648));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1607 (.Y(N5886), .A(N6039), .B(N5909));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1608 (.Y(N6265), .A(N6151), .B(N6590), .C(N6416), .D(N5938));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1609 (.Y(N6436), .A(N6674), .B(N6563), .C(N5943), .D(N6376));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1610 (.Y(N6615), .A(N6641), .B(N5863), .C(N5954), .D(N6281));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1611 (.Y(N5973), .A(N5856), .B(N6383), .C(N6583), .D(N6070));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1612 (.Y(N6504), .A(N6676));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1613 (.Y(N5854), .A(N6213), .B(N6388), .C(N6504), .D(N5886));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1614 (.Y(N6044), .A(N6275), .B(N6490), .C(N6545), .D(N6164));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1615 (.Y(N6231), .A(N6136), .B(N6225), .C(N6115), .D(N6432));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1616 (.Y(N6588), .A(N6425), .B(N6265), .C(N6436), .D(N5973));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1617 (.Y(N5941), .A(N6615));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1618 (.Y(N6123), .A(N6044));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1619 (.Y(N6311), .A(N5941), .B(N6123), .C(N6588), .D(N5854));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1620 (.Y(inst_cellmath__195[15]), .A(N6231), .B(N6311));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1621 (.Y(N6374), .A(N6086), .B(N6551), .C(N6072), .D(N5894));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1622 (.Y(N6549), .A(N6597), .B(N6147), .C(N6372), .D(N5943));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1623 (.Y(N5900), .A(N6650), .B(N6376), .C(N5971), .D(N5954));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1624 (.Y(N6088), .A(N6014), .B(N6455), .C(N6336), .D(N6029));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1625 (.Y(N6452), .A(N6321), .B(N5897), .C(N6411), .D(N6027));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1626 (.Y(N5991), .A(N6374), .B(N6549), .C(N5900), .D(N6088));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1627 (.Y(inst_cellmath__195[16]), .A(N5991), .B(N6452), .C(N6060));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1628 (.Y(N6417), .A(N5909), .B(N6054), .C(N5914), .D(N6674));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1629 (.Y(N6599), .A(N5925), .B(N6096), .C(N6376), .D(N6580));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1630 (.Y(N5953), .A(N6386), .B(N6070), .C(N6275), .D(N5850));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1631 (.Y(N6137), .A(N6490), .B(N5897), .C(N6476), .D(N6545));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1632 (.Y(N6325), .A(N6411), .B(N6643), .C(N6225), .D(N6115));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1633 (.Y(N6493), .A(N6417), .B(N6599), .C(N6325), .D(N5953));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1634 (.Y(inst_cellmath__195[17]), .AN(N6137), .B(N6493));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1635 (.Y(N5917), .A(N5894), .B(N6126), .C(N6461), .D(N5932));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1636 (.Y(N6103), .A(N6590), .B(N6147), .C(N5938), .D(N6665));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1637 (.Y(N6292), .A(N6138), .B(N6024), .C(N6439), .D(N5863));
NAND3XL hyperpropagate_4_1_A_I23862 (.Y(N37712), .A(N5920), .B(N6598), .C(N6050));
NOR2XL hyperpropagate_4_1_A_I23863 (.Y(N5882), .A(N6105), .B(N37712));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1640 (.Y(N6182), .A(N6136), .B(N6208), .C(N6115), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1641 (.Y(N6534), .A(N6606), .B(N5917), .C(N6292), .D(N6103));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1643 (.Y(N6261), .A(N6182));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1644 (.Y(inst_cellmath__195[18]), .A(N5882), .B(N6672), .C(N6261), .D(N6534));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1645 (.Y(N6340), .A(N6461), .B(N6268), .C(N6590), .D(N6147));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1646 (.Y(N6228), .A(N6547), .B(N6310), .C(N6616), .D(N6295));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1647 (.Y(N6400), .A(N6665), .B(N6192), .C(N6623), .D(N6096));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1648 (.Y(N6584), .A(N5856), .B(N6383), .C(N6455), .D(N6518));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1649 (.Y(N5936), .A(N6029), .B(N5920), .C(N6245), .D(N6598));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1650 (.Y(N6116), .A(N6487), .B(N6411), .C(N6533), .D(N6136));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1651 (.Y(N6306), .A(N6340));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1652 (.Y(N6478), .A(N6584));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1653 (.Y(N6658), .A(N6626), .B(N6306), .C(N6478), .D(N6228));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1654 (.Y(inst_cellmath__195[19]), .A(N6400), .B(N5936), .C(N6116), .D(N6658));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1655 (.Y(N6083), .A(N6551), .B(N5894), .C(N6151), .D(N6326));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1656 (.Y(N6277), .A(N6416), .B(N6404), .C(N6563), .D(N5925));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1657 (.Y(N6447), .A(N6650), .B(N6623), .C(N6430), .D(N6024));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1658 (.Y(N5986), .A(N6120), .B(N6086), .C(N6439), .D(N5889));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1659 (.Y(N6166), .A(N6383), .B(N6336), .C(N5920), .D(N6583));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1660 (.Y(N6350), .A(N5916), .B(N6676), .C(N6533), .D(N6180));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1661 (.Y(N5865), .A(N6606), .B(N6083), .C(N6447), .D(N6277));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1662 (.Y(N6051), .A(N5986));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1663 (.Y(N6242), .A(N6350));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1664 (.Y(N6413), .A(N6166));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1665 (.Y(inst_cellmath__195[20]), .A(N6051), .B(N6242), .C(N6413), .D(N5865));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1666 (.Y(N6677), .A(N6674), .B(N6138), .C(N6202), .D(N6120));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1667 (.Y(N5912), .A(N5920), .B(N6583), .C(N6598), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1668 (.Y(N6099), .A(N6338), .B(N6490), .C(N6545), .D(N6411));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1669 (.Y(N6288), .A(N6643), .B(N6208), .C(N6115), .D(N6626));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1670 (.Y(N6639), .A(N6451), .B(N6402), .C(N6193), .D(N6503));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1671 (.Y(N5997), .A(N6606), .B(N6677), .C(N6639), .D(N5912));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1672 (.Y(N6361), .A(N6099));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1673 (.Y(inst_cellmath__195[21]), .AN(N6288), .B(N6361), .C(N5997));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1674 (.Y(N6258), .A(N6600), .B(N6162), .C(N6461));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1675 (.Y(N6609), .A(N5981), .B(N5914), .C(N6674), .D(N6138));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1676 (.Y(N5965), .A(N6430), .B(N5971), .C(N6383), .D(N6455));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1677 (.Y(N6145), .A(N6029), .B(N6583), .C(N6386), .D(N6245));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1678 (.Y(N6334), .A(N5916), .B(N6598), .C(N6321), .D(N6676));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1679 (.Y(N6499), .A(N6291), .B(N6476), .C(N6545), .D(N6027));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1680 (.Y(N5846), .A(N6225), .B(N6115), .C(N6626), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1681 (.Y(N6036), .A(N6258), .B(N5965), .C(N6609), .D(N6145));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1682 (.Y(N6221), .A(N6334));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1683 (.Y(N6395), .A(N5846));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1684 (.Y(N6577), .A(N6499));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1685 (.Y(inst_cellmath__195[22]), .A(N6221), .B(N6395), .C(N6577), .D(N6036));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1686 (.Y(N6301), .A(N6571), .B(N6600), .C(N6162), .D(N6597));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1687 (.Y(N6473), .A(N5932), .B(N6470), .C(N6404), .D(N5943));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1688 (.Y(N6654), .A(N6623), .B(N6430), .C(N6376), .D(N6024));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1689 (.Y(N6009), .A(N6439), .B(N6080), .C(N6281), .D(N5889));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1690 (.Y(N6189), .A(N5856), .B(N6336), .C(N6583), .D(N6070));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1691 (.Y(N6368), .A(N6321), .B(N6676), .C(N5850), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1692 (.Y(N6543), .A(N6476), .B(N6225), .C(N6115), .D(N5969));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1693 (.Y(N6077), .A(N6473), .B(N6301), .C(N6654), .D(N6009));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1694 (.Y(inst_cellmath__195[23]), .A(N6077), .B(N6189), .C(N6543), .D(N6368));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1695 (.Y(N5980), .A(N6660), .B(N6086), .C(N6551), .D(N6072));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1696 (.Y(N6160), .A(N6126), .B(N6507), .C(N6151), .D(N6597));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1697 (.Y(N6347), .A(N6326), .B(N6416), .C(N6372), .D(N5938));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1698 (.Y(N6513), .A(N5914), .B(N6404), .C(N6376), .D(N6439));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1699 (.Y(N5862), .A(N6641), .B(N5863), .C(N6580), .D(N6455));
NAND3XL hyperpropagate_4_1_A_I23864 (.Y(N37720), .A(N6029), .B(N5920), .C(N6598));
NOR2XL hyperpropagate_4_1_A_I23865 (.Y(N6318), .A(N5980), .B(N37720));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1702 (.Y(N6408), .A(N6321), .B(N6676), .C(N6487), .D(N6545));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1703 (.Y(N5946), .A(N6255), .B(N6160), .C(N6347), .D(N5862));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1704 (.Y(N6132), .A(N6513));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1706 (.Y(N6485), .A(N6408));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1707 (.Y(inst_cellmath__195[24]), .A(N6132), .B(N6318), .C(N6485), .D(N5946));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1708 (.Y(N6201), .A(N6072), .B(N6600));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1709 (.Y(N6557), .A(N6126), .B(N6416), .C(N6470), .D(N6372));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1710 (.Y(N5907), .A(N5938), .B(N5914), .C(N5925), .D(N6138));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1711 (.Y(N6095), .A(N5971), .B(N6281), .C(N5856), .D(N6014));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1712 (.Y(N6285), .A(N6383), .B(N6518), .C(N6050), .D(N6321));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1713 (.Y(N6458), .A(N6676), .B(N6275), .C(N6291), .D(N6487));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1714 (.Y(N6635), .A(N6490), .B(N6411), .C(N6626), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1715 (.Y(N5994), .A(N6201), .B(N6557), .C(N6285), .D(N6095));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1716 (.Y(N6174), .A(N5907));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1717 (.Y(N6357), .A(N6635));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1718 (.Y(N6525), .A(N6458));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1719 (.Y(inst_cellmath__195[25]), .A(N6174), .B(N6357), .C(N6525), .D(N5994));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1720 (.Y(N5959), .A(N6372), .B(N5914), .C(N5943), .D(N6650));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1721 (.Y(N6141), .A(N6120), .B(N6244), .C(N6050), .D(N6321));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1722 (.Y(N6033), .AN(N6487), .B(N6201), .C(N6504), .D(N6517));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1723 (.Y(N6391), .A(N6225), .B(N6208), .C(N6180), .D(N6432));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1724 (.Y(N5927), .A(N6425), .B(N6141), .C(N5959), .D(N6391));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1725 (.Y(inst_cellmath__195[26]), .AN(N6328), .B(N6033), .C(N5927));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1726 (.Y(N6538), .A(N6372), .B(N6563), .C(N5889), .D(N6050));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1727 (.Y(N5890), .A(N6321), .B(N6676), .C(N6275), .D(N6338));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1728 (.Y(N6074), .A(N6487), .B(N5850), .C(N6490), .D(N5897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1729 (.Y(N6440), .A(N6600), .B(N6545), .C(N6411), .D(N6164));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1730 (.Y(N6618), .A(N6643), .B(N6027), .C(N6225), .D(N6180));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1731 (.Y(N6156), .A(N6255), .B(N6538), .C(N6618), .D(N5890));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1732 (.Y(N6509), .A(N6440));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1733 (.Y(inst_cellmath__195[27]), .AN(N6074), .B(N6509), .C(N6156));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1734 (.Y(N6127), .A(N6192), .B(N6386), .C(N6370), .D(N5916));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1735 (.Y(N6483), .A(N6291), .B(N6487), .C(N5897), .D(N6476));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1736 (.Y(N6667), .A(N6545), .B(N6411), .C(N6164), .D(N6643));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1737 (.Y(N6018), .A(N6208), .B(N6180), .C(N6115), .D(N6626));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1738 (.Y(N6197), .A(N6042), .B(N6127), .C(N6018), .D(N6218));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1739 (.Y(N6552), .A(N6667));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1740 (.Y(inst_cellmath__195[28]), .AN(N6483), .B(N6552), .C(N6197));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1741 (.Y(N6633), .A(N5954), .B(N6583));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1742 (.Y(N6171), .A(N6370), .B(N6070), .C(N6050), .D(N6321));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1743 (.Y(N6355), .A(N6676), .B(N6275), .C(N6338), .D(N6487));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1744 (.Y(N6521), .A(N5850), .B(N5897), .C(N6476), .D(N6545));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1745 (.Y(N5869), .A(N6411), .B(N6164), .C(N6225), .D(N6208));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1746 (.Y(N6057), .A(N6115), .B(N6626), .C(N6432), .D(N5969));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1747 (.Y(N6248), .A(N6633), .B(N6171), .C(N5869), .D(N6057));
INVX1 inst_cellmath__198_0_I1750 (.Y(N7958), .A(inst_cellmath__61[1]));
INVXL inst_cellmath__198_0_I1751 (.Y(N7696), .A(inst_cellmath__61[2]));
INVXL inst_cellmath__198_0_I1752 (.Y(N7990), .A(inst_cellmath__61[3]));
INVXL inst_cellmath__198_0_I1753 (.Y(N7726), .A(inst_cellmath__61[4]));
INVXL inst_cellmath__198_0_I1754 (.Y(N7842), .A(inst_cellmath__61[5]));
INVXL inst_cellmath__198_0_I1755 (.Y(N7578), .A(inst_cellmath__61[6]));
INVXL inst_cellmath__198_0_I1756 (.Y(N7704), .A(inst_cellmath__61[7]));
INVXL inst_cellmath__198_0_I1757 (.Y(N7823), .A(inst_cellmath__61[8]));
INVXL inst_cellmath__198_0_I1758 (.Y(N7946), .A(inst_cellmath__61[9]));
INVXL inst_cellmath__198_0_I1759 (.Y(N8074), .A(inst_cellmath__61[10]));
INVXL inst_cellmath__198_0_I1760 (.Y(N7627), .A(inst_cellmath__61[11]));
INVXL inst_cellmath__198_0_I1761 (.Y(N7755), .A(inst_cellmath__61[12]));
INVXL inst_cellmath__198_0_I1762 (.Y(N7875), .A(inst_cellmath__61[13]));
INVXL inst_cellmath__198_0_I1763 (.Y(N8000), .A(inst_cellmath__61[14]));
INVXL inst_cellmath__198_0_I1764 (.Y(N7555), .A(inst_cellmath__61[15]));
INVXL inst_cellmath__198_0_I1765 (.Y(N7683), .A(inst_cellmath__115__W1[0]));
XOR2XL inst_cellmath__198_0_I8425 (.Y(N7975), .A(N733), .B(N5778));
NOR2XL inst_cellmath__198_0_I1770 (.Y(N7587), .A(N7975), .B(N7990));
NOR2XL inst_cellmath__198_0_I1771 (.Y(N7833), .A(N7975), .B(N7726));
NOR2XL inst_cellmath__198_0_I1772 (.Y(N8084), .A(N7975), .B(N7842));
NOR2XL inst_cellmath__198_0_I1773 (.Y(N7766), .A(N7975), .B(N7578));
NOR2XL inst_cellmath__198_0_I1774 (.Y(N8010), .A(N7975), .B(N7704));
NOR2XL inst_cellmath__198_0_I1775 (.Y(N7694), .A(N7975), .B(N7823));
NOR2XL inst_cellmath__198_0_I1776 (.Y(N7935), .A(N7975), .B(N7946));
NOR2XL inst_cellmath__198_0_I1777 (.Y(N7616), .A(N7975), .B(N8074));
NOR2XL inst_cellmath__198_0_I1778 (.Y(N7862), .A(N7975), .B(N7627));
NOR2XL inst_cellmath__198_0_I1779 (.Y(N7542), .A(N7975), .B(N7755));
NOR2XL inst_cellmath__198_0_I1780 (.Y(N7791), .A(N7975), .B(N7875));
NOR2XL inst_cellmath__198_0_I1781 (.Y(N8038), .A(N7975), .B(N8000));
NOR2XL inst_cellmath__198_0_I1782 (.Y(N7724), .A(N7975), .B(N7555));
OR2XL inst_cellmath__198_0_I1783 (.Y(N7764), .A(N7975), .B(N7683));
NOR2XL inst_cellmath__198_0_I1784 (.Y(N7681), .A(N7958), .B(N7696));
NOR2XL inst_cellmath__198_0_I1785 (.Y(N7925), .A(N7958), .B(N7990));
NOR2XL inst_cellmath__198_0_I1786 (.Y(N7604), .A(N7958), .B(N7726));
NOR2XL inst_cellmath__198_0_I1787 (.Y(N7851), .A(N7958), .B(N7842));
NOR2XL inst_cellmath__198_0_I1788 (.Y(N7531), .A(N7958), .B(N7578));
NOR2XL inst_cellmath__198_0_I1789 (.Y(N7780), .A(N7958), .B(N7704));
NOR2XL inst_cellmath__198_0_I1790 (.Y(N8027), .A(N7958), .B(N7823));
NOR2XL inst_cellmath__198_0_I1791 (.Y(N7713), .A(N7958), .B(N7946));
NOR2XL inst_cellmath__198_0_I1792 (.Y(N7954), .A(N7958), .B(N8074));
NOR2XL inst_cellmath__198_0_I1793 (.Y(N7637), .A(N7958), .B(N7627));
NOR2XL inst_cellmath__198_0_I1794 (.Y(N7884), .A(N7958), .B(N7755));
NOR2XL inst_cellmath__198_0_I1795 (.Y(N7564), .A(N7958), .B(N7875));
NOR2XL inst_cellmath__198_0_I1796 (.Y(N7809), .A(N7958), .B(N8000));
NOR2XL inst_cellmath__198_0_I1797 (.Y(N8059), .A(N7958), .B(N7555));
OR2XL inst_cellmath__198_0_I1798 (.Y(N7885), .A(N7958), .B(N7683));
INVXL inst_cellmath__198_0_I1799 (.Y(N7517), .A(N7696));
NOR2XL inst_cellmath__198_0_I1800 (.Y(N8014), .A(N7696), .B(N7990));
NOR2XL inst_cellmath__198_0_I1801 (.Y(N7699), .A(N7696), .B(N7726));
NOR2XL inst_cellmath__198_0_I1802 (.Y(N7941), .A(N7696), .B(N7842));
NOR2XL inst_cellmath__198_0_I1803 (.Y(N7621), .A(N7696), .B(N7578));
NOR2XL inst_cellmath__198_0_I1804 (.Y(N7870), .A(N7696), .B(N7704));
NOR2XL inst_cellmath__198_0_I1805 (.Y(N7549), .A(N7696), .B(N7823));
NOR2XL inst_cellmath__198_0_I1806 (.Y(N7798), .A(N7696), .B(N7946));
NOR2XL inst_cellmath__198_0_I1807 (.Y(N8046), .A(N7696), .B(N8074));
NOR2XL inst_cellmath__198_0_I1808 (.Y(N7730), .A(N7696), .B(N7627));
NOR2XL inst_cellmath__198_0_I1809 (.Y(N7971), .A(N7696), .B(N7755));
NOR2XL inst_cellmath__198_0_I1810 (.Y(N7655), .A(N7696), .B(N7875));
NOR2XL inst_cellmath__198_0_I1811 (.Y(N7900), .A(N7696), .B(N8000));
NOR2XL inst_cellmath__198_0_I1812 (.Y(N7582), .A(N7696), .B(N7555));
OR2XL inst_cellmath__198_0_I1813 (.Y(N8007), .A(N7696), .B(N7683));
INVXL inst_cellmath__198_0_I1814 (.Y(N7608), .A(N7990));
NOR2XL inst_cellmath__198_0_I1815 (.Y(N7536), .A(N7990), .B(N7726));
NOR2XL inst_cellmath__198_0_I1816 (.Y(N7785), .A(N7990), .B(N7842));
NOR2XL inst_cellmath__198_0_I1817 (.Y(N8033), .A(N7990), .B(N7578));
NOR2XL inst_cellmath__198_0_I1818 (.Y(N7718), .A(N7990), .B(N7704));
NOR2XL inst_cellmath__198_0_I1819 (.Y(N7961), .A(N7990), .B(N7823));
NOR2XL inst_cellmath__198_0_I1820 (.Y(N7643), .A(N7990), .B(N7946));
NOR2XL inst_cellmath__198_0_I1821 (.Y(N7890), .A(N7990), .B(N8074));
NOR2XL inst_cellmath__198_0_I1822 (.Y(N7570), .A(N7990), .B(N7627));
NOR2XL inst_cellmath__198_0_I1823 (.Y(N7816), .A(N7990), .B(N7755));
NOR2XL inst_cellmath__198_0_I1824 (.Y(N8065), .A(N7990), .B(N7875));
NOR2XL inst_cellmath__198_0_I1825 (.Y(N7749), .A(N7990), .B(N8000));
NOR2XL inst_cellmath__198_0_I1826 (.Y(N7992), .A(N7990), .B(N7555));
OR2XL inst_cellmath__198_0_I1827 (.Y(N7565), .A(N7990), .B(N7683));
INVXL inst_cellmath__198_0_I1828 (.Y(N8020), .A(N7726));
NOR2XL inst_cellmath__198_0_I1829 (.Y(N7948), .A(N7726), .B(N7842));
NOR2XL inst_cellmath__198_0_I1830 (.Y(N7630), .A(N7726), .B(N7578));
NOR2XL inst_cellmath__198_0_I1831 (.Y(N7877), .A(N7726), .B(N7704));
NOR2XL inst_cellmath__198_0_I1832 (.Y(N7557), .A(N7726), .B(N7823));
NOR2XL inst_cellmath__198_0_I1833 (.Y(N7804), .A(N7726), .B(N7946));
NOR2XL inst_cellmath__198_0_I1834 (.Y(N8053), .A(N7726), .B(N8074));
NOR2XL inst_cellmath__198_0_I1835 (.Y(N7737), .A(N7726), .B(N7627));
NOR2XL inst_cellmath__198_0_I1836 (.Y(N7977), .A(N7726), .B(N7755));
NOR2XL inst_cellmath__198_0_I1837 (.Y(N7664), .A(N7726), .B(N7875));
NOR2XL inst_cellmath__198_0_I1838 (.Y(N7906), .A(N7726), .B(N8000));
NOR2XL inst_cellmath__198_0_I1839 (.Y(N7588), .A(N7726), .B(N7555));
OR2XL inst_cellmath__198_0_I1840 (.Y(N7693), .A(N7726), .B(N7683));
INVXL inst_cellmath__198_0_I1841 (.Y(N7617), .A(N7842));
NOR2XL inst_cellmath__198_0_I1842 (.Y(N7543), .A(N7842), .B(N7578));
NOR2XL inst_cellmath__198_0_I1843 (.Y(N7792), .A(N7842), .B(N7704));
NOR2XL inst_cellmath__198_0_I1844 (.Y(N8040), .A(N7842), .B(N7823));
NOR2XL inst_cellmath__198_0_I1845 (.Y(N7725), .A(N7842), .B(N7946));
NOR2XL inst_cellmath__198_0_I1846 (.Y(N7967), .A(N7842), .B(N8074));
NOR2XL inst_cellmath__198_0_I1847 (.Y(N7649), .A(N7842), .B(N7627));
NOR2XL inst_cellmath__198_0_I1848 (.Y(N7895), .A(N7842), .B(N7755));
NOR2XL inst_cellmath__198_0_I1849 (.Y(N7577), .A(N7842), .B(N7875));
NOR2XL inst_cellmath__198_0_I1850 (.Y(N7822), .A(N7842), .B(N8000));
NOR2XL inst_cellmath__198_0_I1851 (.Y(N8073), .A(N7842), .B(N7555));
OR2XL inst_cellmath__198_0_I1852 (.Y(N7811), .A(N7842), .B(N7683));
INVXL inst_cellmath__198_0_I1853 (.Y(N7532), .A(N7578));
NOR2XL inst_cellmath__198_0_I1854 (.Y(N8029), .A(N7578), .B(N7704));
NOR2XL inst_cellmath__198_0_I1855 (.Y(N7714), .A(N7578), .B(N7823));
NOR2XL inst_cellmath__198_0_I1856 (.Y(N7955), .A(N7578), .B(N7946));
NOR2XL inst_cellmath__198_0_I1857 (.Y(N7639), .A(N7578), .B(N8074));
NOR2XL inst_cellmath__198_0_I1858 (.Y(N7886), .A(N7578), .B(N7627));
NOR2XL inst_cellmath__198_0_I1859 (.Y(N7566), .A(N7578), .B(N7755));
NOR2XL inst_cellmath__198_0_I1860 (.Y(N7813), .A(N7578), .B(N7875));
NOR2XL inst_cellmath__198_0_I1861 (.Y(N8061), .A(N7578), .B(N8000));
NOR2XL inst_cellmath__198_0_I1862 (.Y(N7745), .A(N7578), .B(N7555));
OR2XL inst_cellmath__198_0_I1863 (.Y(N7933), .A(N7578), .B(N7683));
INVXL inst_cellmath__198_0_I1864 (.Y(N7770), .A(N7704));
NOR2XL inst_cellmath__198_0_I1865 (.Y(N7702), .A(N7704), .B(N7823));
NOR2XL inst_cellmath__198_0_I1866 (.Y(N7943), .A(N7704), .B(N7946));
NOR2XL inst_cellmath__198_0_I1867 (.Y(N7624), .A(N7704), .B(N8074));
NOR2XL inst_cellmath__198_0_I1868 (.Y(N7873), .A(N7704), .B(N7627));
NOR2XL inst_cellmath__198_0_I1869 (.Y(N7551), .A(N7704), .B(N7755));
NOR2XL inst_cellmath__198_0_I1870 (.Y(N7801), .A(N7704), .B(N7875));
NOR2XL inst_cellmath__198_0_I1871 (.Y(N8049), .A(N7704), .B(N8000));
NOR2XL inst_cellmath__198_0_I1872 (.Y(N7732), .A(N7704), .B(N7555));
OR2XL inst_cellmath__198_0_I1873 (.Y(N8060), .A(N7704), .B(N7683));
INVXL inst_cellmath__198_0_I1874 (.Y(N7762), .A(N7823));
NOR2XL inst_cellmath__198_0_I1875 (.Y(N7690), .A(N7823), .B(N7946));
NOR2XL inst_cellmath__198_0_I1876 (.Y(N7932), .A(N7823), .B(N8074));
NOR2XL inst_cellmath__198_0_I1877 (.Y(N7611), .A(N7823), .B(N7627));
NOR2XL inst_cellmath__198_0_I1878 (.Y(N7859), .A(N7823), .B(N7755));
NOR2XL inst_cellmath__198_0_I1879 (.Y(N7539), .A(N7823), .B(N7875));
NOR2XL inst_cellmath__198_0_I1880 (.Y(N7788), .A(N7823), .B(N8000));
NOR2XL inst_cellmath__198_0_I1881 (.Y(N8035), .A(N7823), .B(N7555));
OR2XL inst_cellmath__198_0_I1882 (.Y(N7613), .A(N7823), .B(N7683));
INVXL inst_cellmath__198_0_I1883 (.Y(N8068), .A(N7946));
NOR2XL inst_cellmath__198_0_I1884 (.Y(N7994), .A(N7946), .B(N8074));
NOR2XL inst_cellmath__198_0_I1885 (.Y(N7677), .A(N7946), .B(N7627));
NOR2XL inst_cellmath__198_0_I1886 (.Y(N7920), .A(N7946), .B(N7755));
NOR2XL inst_cellmath__198_0_I1887 (.Y(N7599), .A(N7946), .B(N7875));
NOR2XL inst_cellmath__198_0_I1888 (.Y(N7847), .A(N7946), .B(N8000));
NOR2XL inst_cellmath__198_0_I1889 (.Y(N7527), .A(N7946), .B(N7555));
OR2XL inst_cellmath__198_0_I1890 (.Y(N7744), .A(N7946), .B(N7683));
INVXL inst_cellmath__198_0_I1891 (.Y(N7560), .A(N8074));
NOR2XL inst_cellmath__198_0_I1892 (.Y(N8057), .A(N8074), .B(N7627));
NOR2XL inst_cellmath__198_0_I1893 (.Y(N7741), .A(N8074), .B(N7755));
NOR2XL inst_cellmath__198_0_I1894 (.Y(N7981), .A(N8074), .B(N7875));
NOR2XL inst_cellmath__198_0_I1895 (.Y(N7667), .A(N8074), .B(N8000));
NOR2XL inst_cellmath__198_0_I1896 (.Y(N7910), .A(N8074), .B(N7555));
OR2XL inst_cellmath__198_0_I1897 (.Y(N7861), .A(N8074), .B(N7683));
INVXL inst_cellmath__198_0_I1898 (.Y(N7938), .A(N7627));
NOR2XL inst_cellmath__198_0_I1899 (.Y(N7867), .A(N7627), .B(N7755));
NOR2XL inst_cellmath__198_0_I1900 (.Y(N7546), .A(N7627), .B(N7875));
NOR2XL inst_cellmath__198_0_I1901 (.Y(N7794), .A(N7627), .B(N8000));
NOR2XL inst_cellmath__198_0_I1902 (.Y(N8043), .A(N7627), .B(N7555));
OR2XL inst_cellmath__198_0_I1903 (.Y(N7986), .A(N7627), .B(N7683));
INVXL inst_cellmath__198_0_I1904 (.Y(N8077), .A(N7755));
NOR2XL inst_cellmath__198_0_I1905 (.Y(N8002), .A(N7755), .B(N7875));
NOR2XL inst_cellmath__198_0_I1906 (.Y(N7685), .A(N7755), .B(N8000));
NOR2XL inst_cellmath__198_0_I1907 (.Y(N7927), .A(N7755), .B(N7555));
OR2XL inst_cellmath__198_0_I1908 (.Y(N7540), .A(N7755), .B(N7683));
INVXL inst_cellmath__198_0_I1909 (.Y(N7957), .A(N7875));
NOR2XL inst_cellmath__198_0_I1910 (.Y(N7888), .A(N7875), .B(N8000));
NOR2XL inst_cellmath__198_0_I1911 (.Y(N7568), .A(N7875), .B(N7555));
OR2XL inst_cellmath__198_0_I1912 (.Y(N7670), .A(N7875), .B(N7683));
INVXL inst_cellmath__198_0_I1913 (.Y(N7595), .A(N8000));
NOR2XL inst_cellmath__198_0_I1914 (.Y(N7522), .A(N8000), .B(N7555));
OR2XL inst_cellmath__198_0_I1915 (.Y(N7789), .A(N8000), .B(N7683));
INVXL inst_cellmath__198_0_I1916 (.Y(N7554), .A(N7555));
ADDHX1 inst_cellmath__198_0_I1917 (.CO(N8037), .S(N7914), .A(N7587), .B(N7681));
ADDHX1 inst_cellmath__198_0_I1918 (.CO(N7722), .S(N7593), .A(N7925), .B(N7833));
ADDHX1 inst_cellmath__198_0_I1919 (.CO(N7965), .S(N7840), .A(N8084), .B(N7608));
ADDFX1 inst_cellmath__198_0_I1920 (.CO(N7646), .S(N7518), .A(N8014), .B(N7604), .CI(N7840));
ADDHX1 inst_cellmath__198_0_I1921 (.CO(N7892), .S(N7769), .A(N7851), .B(N7766));
ADDFX1 inst_cellmath__198_0_I1922 (.CO(N7574), .S(N8015), .A(N7965), .B(N7699), .CI(N7769));
ADDHX1 inst_cellmath__198_0_I1923 (.CO(N7819), .S(N7700), .A(N8010), .B(N7536));
ADDFX1 inst_cellmath__198_0_I1924 (.CO(N8069), .S(N7942), .A(N8020), .B(N7531), .CI(N7941));
ADDFX1 inst_cellmath__198_0_I1925 (.CO(N7752), .S(N7622), .A(N7700), .B(N7892), .CI(N7942));
ADDHX1 inst_cellmath__198_0_I1926 (.CO(N7996), .S(N7871), .A(N7780), .B(N7785));
ADDFX1 inst_cellmath__198_0_I1927 (.CO(N7678), .S(N7550), .A(N7621), .B(N7694), .CI(N7819));
ADDFX1 inst_cellmath__198_0_I1928 (.CO(N7922), .S(N7799), .A(N8069), .B(N7871), .CI(N7550));
ADDHX1 inst_cellmath__198_0_I1929 (.CO(N7601), .S(N8047), .A(N7935), .B(N7617));
ADDFX1 inst_cellmath__198_0_I1930 (.CO(N7848), .S(N7731), .A(N8027), .B(N8033), .CI(N7948));
ADDFX1 inst_cellmath__198_0_I1931 (.CO(N7528), .S(N7972), .A(N7996), .B(N7870), .CI(N8047));
ADDFX1 inst_cellmath__198_0_I1932 (.CO(N7777), .S(N7656), .A(N7731), .B(N7678), .CI(N7972));
ADDHX1 inst_cellmath__198_0_I1933 (.CO(N8024), .S(N7901), .A(N7713), .B(N7718));
ADDFX1 inst_cellmath__198_0_I1934 (.CO(N7710), .S(N7583), .A(N7630), .B(N7616), .CI(N7549));
ADDFX1 inst_cellmath__198_0_I1935 (.CO(N7951), .S(N7828), .A(N7901), .B(N7601), .CI(N7848));
ADDFX1 inst_cellmath__198_0_I1936 (.CO(N7634), .S(N8081), .A(N7583), .B(N7528), .CI(N7828));
ADDHX1 inst_cellmath__198_0_I1937 (.CO(N7881), .S(N7760), .A(N7862), .B(N7543));
ADDFX1 inst_cellmath__198_0_I1938 (.CO(N7561), .S(N8005), .A(N7954), .B(N7961), .CI(N7798));
ADDFX1 inst_cellmath__198_0_I1939 (.CO(N7806), .S(N7689), .A(N7877), .B(N7532), .CI(N8024));
ADDFX1 inst_cellmath__198_0_I1940 (.CO(N8058), .S(N7930), .A(N7710), .B(N7760), .CI(N8005));
ADDFX1 inst_cellmath__198_0_I1941 (.CO(N7742), .S(N7609), .A(N7951), .B(N7689), .CI(N7930));
ADDHX1 inst_cellmath__198_0_I1942 (.CO(N7983), .S(N7858), .A(N7637), .B(N7643));
ADDFX1 inst_cellmath__198_0_I1943 (.CO(N7668), .S(N7537), .A(N7542), .B(N7792), .CI(N7557));
ADDFX1 inst_cellmath__198_0_I1944 (.CO(N7912), .S(N7786), .A(N7881), .B(N8046), .CI(N7858));
ADDFX1 inst_cellmath__198_0_I1945 (.CO(N7591), .S(N8034), .A(N7806), .B(N7561), .CI(N7537));
ADDFX1 inst_cellmath__198_0_I1946 (.CO(N7838), .S(N7719), .A(N8058), .B(N7786), .CI(N8034));
ADDHX1 inst_cellmath__198_0_I1947 (.CO(N7515), .S(N7962), .A(N7770), .B(N7791));
ADDFX1 inst_cellmath__198_0_I1948 (.CO(N7768), .S(N7644), .A(N7890), .B(N8040), .CI(N7730));
ADDFX1 inst_cellmath__198_0_I1949 (.CO(N8013), .S(N7891), .A(N8029), .B(N7884), .CI(N7804));
ADDFX1 inst_cellmath__198_0_I1950 (.CO(N7698), .S(N7571), .A(N7962), .B(N7983), .CI(N7668));
ADDFX1 inst_cellmath__198_0_I1951 (.CO(N7939), .S(N7817), .A(N7912), .B(N7644), .CI(N7891));
ADDFX1 inst_cellmath__198_0_I1952 (.CO(N7619), .S(N8066), .A(N7591), .B(N7571), .CI(N7817));
ADDHX1 inst_cellmath__198_0_I1953 (.CO(N7868), .S(N7750), .A(N7564), .B(N7570));
ADDFX1 inst_cellmath__198_0_I1954 (.CO(N7548), .S(N7993), .A(N8038), .B(N7725), .CI(N7971));
ADDFX1 inst_cellmath__198_0_I1955 (.CO(N7796), .S(N7675), .A(N8053), .B(N7714), .CI(N7515));
ADDFX1 inst_cellmath__198_0_I1956 (.CO(N8044), .S(N7918), .A(N7768), .B(N7750), .CI(N8013));
ADDFX1 inst_cellmath__198_0_I1957 (.CO(N7729), .S(N7598), .A(N7675), .B(N7993), .CI(N7698));
ADDFX1 inst_cellmath__198_0_I1958 (.CO(N7970), .S(N7844), .A(N7939), .B(N7918), .CI(N7598));
ADDHX1 inst_cellmath__198_0_I1959 (.CO(N7652), .S(N7524), .A(N7724), .B(N7702));
ADDFX1 inst_cellmath__198_0_I1960 (.CO(N7898), .S(N7774), .A(N7809), .B(N7762), .CI(N7655));
ADDFX1 inst_cellmath__198_0_I1961 (.CO(N7580), .S(N8021), .A(N7816), .B(N7967), .CI(N7737));
ADDFX1 inst_cellmath__198_0_I1962 (.CO(N7826), .S(N7706), .A(N7868), .B(N7955), .CI(N7524));
ADDFX1 inst_cellmath__198_0_I1963 (.CO(N8078), .S(N7949), .A(N7796), .B(N7548), .CI(N8021));
ADDFX1 inst_cellmath__198_0_I1964 (.CO(N7757), .S(N7631), .A(N8044), .B(N7774), .CI(N7706));
ADDFX1 inst_cellmath__198_0_I1965 (.CO(N8003), .S(N7878), .A(N7949), .B(N7729), .CI(N7631));
XNOR2X1 inst_cellmath__198_0_I1966 (.Y(N7558), .A(N8059), .B(N8065));
OR2XL inst_cellmath__198_0_I1967 (.Y(N7687), .A(N8059), .B(N8065));
ADDFX1 inst_cellmath__198_0_I1968 (.CO(N7606), .S(N8054), .A(N7649), .B(N7943), .CI(N7639));
ADDFX1 inst_cellmath__198_0_I1969 (.CO(N7855), .S(N7738), .A(N7764), .B(N7977), .CI(N7900));
ADDFX1 inst_cellmath__198_0_I1970 (.CO(N7534), .S(N7978), .A(N7558), .B(N7652), .CI(N7580));
ADDFX1 inst_cellmath__198_0_I1971 (.CO(N7783), .S(N7665), .A(N8054), .B(N7898), .CI(N7738));
ADDFX1 inst_cellmath__198_0_I1972 (.CO(N8031), .S(N7907), .A(N7978), .B(N7826), .CI(N8078));
ADDFX1 inst_cellmath__198_0_I1973 (.CO(N7716), .S(N7589), .A(N7757), .B(N7665), .CI(N7907));
ADDFX1 inst_cellmath__198_0_I1974 (.CO(N7959), .S(N7834), .A(N7624), .B(N8068), .CI(N7885));
ADDFX1 inst_cellmath__198_0_I1975 (.CO(N7642), .S(N8088), .A(N7749), .B(N7895), .CI(N7582));
ADDFX1 inst_cellmath__198_0_I1976 (.CO(N7889), .S(N7767), .A(N7886), .B(N7690), .CI(N7664));
ADDFX1 inst_cellmath__198_0_I1977 (.CO(N7569), .S(N8011), .A(N7606), .B(N7687), .CI(N7855));
ADDFX1 inst_cellmath__198_0_I1978 (.CO(N7815), .S(N7697), .A(N8088), .B(N7834), .CI(N7767));
ADDFX1 inst_cellmath__198_0_I1979 (.CO(N8064), .S(N7936), .A(N8011), .B(N7534), .CI(N7783));
ADDFX1 inst_cellmath__198_0_I1980 (.CO(N7748), .S(N7618), .A(N8031), .B(N7697), .CI(N7936));
ADDFX1 inst_cellmath__198_0_I1981 (.CO(N7989), .S(N7865), .A(N7577), .B(N7873), .CI(N7992));
ADDFX1 inst_cellmath__198_0_I1982 (.CO(N7674), .S(N7544), .A(N7566), .B(N7932), .CI(N7906));
ADDFX1 inst_cellmath__198_0_I1983 (.CO(N7916), .S(N7793), .A(N7959), .B(N8007), .CI(N7889));
ADDFX1 inst_cellmath__198_0_I1984 (.CO(N7596), .S(N8041), .A(N7865), .B(N7642), .CI(N7544));
ADDFX1 inst_cellmath__198_0_I1985 (.CO(N7843), .S(N7727), .A(N7815), .B(N7569), .CI(N7793));
ADDFX1 inst_cellmath__198_0_I1986 (.CO(N7523), .S(N7968), .A(N8064), .B(N8041), .CI(N7727));
ADDFX1 inst_cellmath__198_0_I1987 (.CO(N7772), .S(N7650), .A(N7994), .B(N7560), .CI(N7565));
ADDFX1 inst_cellmath__198_0_I1988 (.CO(N8019), .S(N7896), .A(N7822), .B(N7551), .CI(N7588));
ADDFX1 inst_cellmath__198_0_I1989 (.CO(N7705), .S(N7579), .A(N7813), .B(N7611), .CI(N7989));
ADDFX1 inst_cellmath__198_0_I1990 (.CO(N7947), .S(N7824), .A(N7650), .B(N7674), .CI(N7896));
ADDFX1 inst_cellmath__198_0_I1991 (.CO(N7628), .S(N8075), .A(N7579), .B(N7916), .CI(N7596));
ADDFX1 inst_cellmath__198_0_I1992 (.CO(N7876), .S(N7756), .A(N7843), .B(N7824), .CI(N8075));
ADDFX1 inst_cellmath__198_0_I1993 (.CO(N7556), .S(N8001), .A(N7801), .B(N7677), .CI(N8073));
ADDFX1 inst_cellmath__198_0_I1994 (.CO(N7803), .S(N7684), .A(N8061), .B(N7859), .CI(N7693));
ADDFX1 inst_cellmath__198_0_I1995 (.CO(N8052), .S(N7926), .A(N8019), .B(N7772), .CI(N8001));
ADDFX1 inst_cellmath__198_0_I1996 (.CO(N7736), .S(N7605), .A(N7705), .B(N7684), .CI(N7947));
ADDFX1 inst_cellmath__198_0_I1997 (.CO(N7976), .S(N7853), .A(N7628), .B(N7926), .CI(N7605));
ADDFX1 inst_cellmath__198_0_I1998 (.CO(N7662), .S(N7533), .A(N7920), .B(N7938), .CI(N7811));
ADDFX1 inst_cellmath__198_0_I1999 (.CO(N7905), .S(N7782), .A(N7745), .B(N8049), .CI(N7539));
ADDFX1 inst_cellmath__198_0_I2000 (.CO(N7586), .S(N8030), .A(N7556), .B(N8057), .CI(N7803));
ADDFX1 inst_cellmath__198_0_I2001 (.CO(N7832), .S(N7715), .A(N7782), .B(N7533), .CI(N8052));
ADDFX1 inst_cellmath__198_0_I2002 (.CO(N8086), .S(N7956), .A(N7736), .B(N8030), .CI(N7715));
ADDFX1 inst_cellmath__198_0_I2003 (.CO(N7765), .S(N7641), .A(N7732), .B(N7599), .CI(N7741));
ADDFX1 inst_cellmath__198_0_I2004 (.CO(N8009), .S(N7887), .A(N7933), .B(N7788), .CI(N7662));
ADDFX1 inst_cellmath__198_0_I2005 (.CO(N7695), .S(N7567), .A(N7641), .B(N7905), .CI(N7586));
ADDFX1 inst_cellmath__198_0_I2006 (.CO(N7934), .S(N7814), .A(N7832), .B(N7887), .CI(N7567));
ADDFX1 inst_cellmath__198_0_I2007 (.CO(N7615), .S(N8062), .A(N7867), .B(N8077), .CI(N8060));
ADDFX1 inst_cellmath__198_0_I2008 (.CO(N7864), .S(N7747), .A(N8035), .B(N7847), .CI(N7981));
ADDFX1 inst_cellmath__198_0_I2009 (.CO(N7541), .S(N7987), .A(N8062), .B(N7765), .CI(N7747));
ADDFX1 inst_cellmath__198_0_I2010 (.CO(N7790), .S(N7672), .A(N7695), .B(N8009), .CI(N7987));
ADDFX1 inst_cellmath__198_0_I2011 (.CO(N8039), .S(N7915), .A(N7527), .B(N7546), .CI(N7667));
ADDFX1 inst_cellmath__198_0_I2012 (.CO(N7723), .S(N7594), .A(N7615), .B(N7613), .CI(N7864));
ADDFX1 inst_cellmath__198_0_I2013 (.CO(N7966), .S(N7841), .A(N7541), .B(N7915), .CI(N7594));
ADDFX1 inst_cellmath__198_0_I2014 (.CO(N7648), .S(N7521), .A(N8002), .B(N7957), .CI(N7744));
ADDFX1 inst_cellmath__198_0_I2015 (.CO(N7894), .S(N7771), .A(N7910), .B(N7794), .CI(N8039));
ADDFX1 inst_cellmath__198_0_I2016 (.CO(N7576), .S(N8017), .A(N7723), .B(N7521), .CI(N7771));
ADDFX1 inst_cellmath__198_0_I2017 (.CO(N7821), .S(N7703), .A(N7685), .B(N8043), .CI(N7861));
ADDFX1 inst_cellmath__198_0_I2018 (.CO(N8072), .S(N7945), .A(N7703), .B(N7648), .CI(N7894));
ADDFX1 inst_cellmath__198_0_I2019 (.CO(N7754), .S(N7626), .A(N7927), .B(N7595), .CI(N7986));
ADDFX1 inst_cellmath__198_0_I2020 (.CO(N7998), .S(N7874), .A(N7821), .B(N7888), .CI(N7626));
ADDFX1 inst_cellmath__198_0_I2021 (.CO(N7680), .S(N7553), .A(N7540), .B(N7568), .CI(N7754));
ADDFX1 inst_cellmath__198_0_I2022 (.CO(N7924), .S(N7802), .A(N7522), .B(N7554), .CI(N7670));
AND2XL inst_cellmath__198_0_I2025 (.Y(N7850), .A(N7517), .B(N7914));
NOR2XL inst_cellmath__198_0_I2026 (.Y(N7974), .A(N8037), .B(N7593));
NAND2XL inst_cellmath__198_0_I2027 (.Y(N7530), .A(N8037), .B(N7593));
AND2XL inst_cellmath__198_0_I2029 (.Y(N7779), .A(N7722), .B(N7518));
NOR2XL inst_cellmath__198_0_I2030 (.Y(N7903), .A(N7646), .B(N8015));
NAND2XL inst_cellmath__198_0_I2031 (.Y(N8026), .A(N7646), .B(N8015));
AND2XL inst_cellmath__198_0_I2033 (.Y(N7712), .A(N7574), .B(N7622));
NOR2XL inst_cellmath__198_0_I2034 (.Y(N7830), .A(N7752), .B(N7799));
NAND2XL inst_cellmath__198_0_I2035 (.Y(N7953), .A(N7752), .B(N7799));
NOR2XL inst_cellmath__198_0_I2036 (.Y(N8083), .A(N7922), .B(N7656));
NAND2XL inst_cellmath__198_0_I2037 (.Y(N7636), .A(N7922), .B(N7656));
AND2XL inst_cellmath__198_0_I2039 (.Y(N7883), .A(N7777), .B(N8081));
NOR2XL inst_cellmath__198_0_I2040 (.Y(N8006), .A(N7634), .B(N7609));
NAND2XL inst_cellmath__198_0_I2041 (.Y(N7563), .A(N7634), .B(N7609));
NOR2XL inst_cellmath__198_0_I2042 (.Y(N7692), .A(N7742), .B(N7719));
NAND2XL inst_cellmath__198_0_I2043 (.Y(N7808), .A(N7742), .B(N7719));
NOR3XL inst_cellmath__198_0_I8489 (.Y(N7612), .A(N7975), .B(N7958), .C(N7696));
OAI22XL inst_cellmath__198_0_I8428 (.Y(N7721), .A0(N7850), .A1(N7612), .B0(N7517), .B1(N7914));
AOI21XL inst_cellmath__198_0_I2048 (.Y(N7573), .A0(N7530), .A1(N7721), .B0(N7974));
OAI22XL inst_cellmath__198_0_I8429 (.Y(N7921), .A0(N7779), .A1(N7573), .B0(N7722), .B1(N7518));
AOI21XL inst_cellmath__198_0_I2052 (.Y(N7709), .A0(N8026), .A1(N7921), .B0(N7903));
OAI22XL inst_cellmath__198_0_I8430 (.Y(N7982), .A0(N7712), .A1(N7709), .B0(N7574), .B1(N7622));
AOI21XL inst_cellmath__198_0_I2056 (.Y(N7911), .A0(N7636), .A1(N7830), .B0(N8083));
INVXL inst_cellmath__198_0_I2057 (.Y(N7520), .A(N7911));
AOI31X1 inst_cellmath__198_0_I2059 (.Y(N7795), .A0(N7636), .A1(N7953), .A2(N7982), .B0(N7520));
OAI22XL inst_cellmath__198_0_I8431 (.Y(N7686), .A0(N7883), .A1(N7795), .B0(N7777), .B1(N8081));
AO21XL inst_cellmath__198_0_I2063 (.Y(N7660), .A0(N7808), .A1(N8006), .B0(N7692));
AOI31X1 inst_cellmath__198_0_I2065 (.Y(N7673), .A0(N7808), .A1(N7563), .A2(N7686), .B0(N7660));
NOR2XL inst_cellmath__198_0_I2090 (.Y(N8016), .A(N7619), .B(N7844));
XOR2XL inst_cellmath__198_0_I2091 (.Y(N7575), .A(N7619), .B(N7844));
NOR2XL inst_cellmath__198_0_I2092 (.Y(N7701), .A(N7970), .B(N7878));
XOR2XL inst_cellmath__198_0_I2093 (.Y(N7820), .A(N7970), .B(N7878));
NOR2XL inst_cellmath__198_0_I2094 (.Y(N7944), .A(N8003), .B(N7589));
XOR2XL inst_cellmath__198_0_I2095 (.Y(N8070), .A(N8003), .B(N7589));
NOR2XL inst_cellmath__198_0_I2096 (.Y(N7623), .A(N7716), .B(N7618));
XOR2XL inst_cellmath__198_0_I2097 (.Y(N7753), .A(N7716), .B(N7618));
NOR2XL inst_cellmath__198_0_I2098 (.Y(N7872), .A(N7748), .B(N7968));
XOR2XL inst_cellmath__198_0_I2099 (.Y(N7997), .A(N7748), .B(N7968));
NOR2XL inst_cellmath__198_0_I2100 (.Y(N7552), .A(N7523), .B(N7756));
XOR2XL inst_cellmath__198_0_I2101 (.Y(N7679), .A(N7523), .B(N7756));
NOR2XL inst_cellmath__198_0_I2102 (.Y(N7800), .A(N7876), .B(N7853));
XOR2XL inst_cellmath__198_0_I2103 (.Y(N7923), .A(N7876), .B(N7853));
NOR2XL inst_cellmath__198_0_I2104 (.Y(N8048), .A(N7976), .B(N7956));
XOR2XL inst_cellmath__198_0_I2105 (.Y(N7602), .A(N7976), .B(N7956));
NOR2XL inst_cellmath__198_0_I2106 (.Y(N7733), .A(N8086), .B(N7814));
XOR2XL inst_cellmath__198_0_I2107 (.Y(N7849), .A(N8086), .B(N7814));
NOR2XL inst_cellmath__198_0_I2108 (.Y(N7973), .A(N7934), .B(N7672));
XOR2XL inst_cellmath__198_0_I2109 (.Y(N7529), .A(N7934), .B(N7672));
NOR2XL inst_cellmath__198_0_I2110 (.Y(N7657), .A(N7790), .B(N7841));
XOR2XL inst_cellmath__198_0_I2111 (.Y(N7778), .A(N7790), .B(N7841));
NOR2XL inst_cellmath__198_0_I2112 (.Y(N7902), .A(N7966), .B(N8017));
XOR2XL inst_cellmath__198_0_I2113 (.Y(N8025), .A(N7966), .B(N8017));
NOR2XL inst_cellmath__198_0_I2114 (.Y(N7584), .A(N7945), .B(N7576));
XOR2XL inst_cellmath__198_0_I2115 (.Y(N7711), .A(N7945), .B(N7576));
NOR2XL inst_cellmath__198_0_I2116 (.Y(N7829), .A(N8072), .B(N7874));
XOR2XL inst_cellmath__198_0_I2117 (.Y(N7952), .A(N8072), .B(N7874));
NOR2XL inst_cellmath__198_0_I2118 (.Y(N8082), .A(N7553), .B(N7998));
XOR2XL inst_cellmath__198_0_I2119 (.Y(N7635), .A(N7553), .B(N7998));
NOR2XL inst_cellmath__198_0_I2120 (.Y(N7761), .A(N7802), .B(N7680));
XOR2XL inst_cellmath__198_0_I2121 (.Y(N7882), .A(N7802), .B(N7680));
XNOR2X1 inst_cellmath__198_0_I2122 (.Y(N7825), .A(N7789), .B(N7924));
NAND2BXL inst_cellmath__198_0_I2123 (.Y(N7807), .AN(N7683), .B(N7555));
OR2XL cmp_A_I8515 (.Y(N19018), .A(N7838), .B(N8066));
AO22XL cmp_A_I8516 (.Y(N7931), .A0(N19018), .A1(N7673), .B0(N7838), .B1(N8066));
AOI21XL inst_cellmath__198_0_I2125 (.Y(N7610), .A0(N7820), .A1(N8016), .B0(N7701));
NAND2XL inst_cellmath__198_0_I2126 (.Y(N7743), .A(N7820), .B(N7575));
AOI21XL inst_cellmath__198_0_I2127 (.Y(N7860), .A0(N7753), .A1(N7944), .B0(N7623));
NAND2XL inst_cellmath__198_0_I2128 (.Y(N7984), .A(N7753), .B(N8070));
AOI21XL inst_cellmath__198_0_I2129 (.Y(N7538), .A0(N7679), .A1(N7872), .B0(N7552));
NAND2XL inst_cellmath__198_0_I2130 (.Y(N7669), .A(N7679), .B(N7997));
AOI21XL inst_cellmath__198_0_I2131 (.Y(N7787), .A0(N7602), .A1(N7800), .B0(N8048));
NAND2XL inst_cellmath__198_0_I2132 (.Y(N7913), .A(N7602), .B(N7923));
AOI21XL inst_cellmath__198_0_I2133 (.Y(N8036), .A0(N7529), .A1(N7733), .B0(N7973));
NAND2XL inst_cellmath__198_0_I2134 (.Y(N7592), .A(N7529), .B(N7849));
AOI21XL inst_cellmath__198_0_I2135 (.Y(N7720), .A0(N8025), .A1(N7657), .B0(N7902));
NAND2XL inst_cellmath__198_0_I2136 (.Y(N7839), .A(N8025), .B(N7778));
AOI21XL inst_cellmath__198_0_I2137 (.Y(N7963), .A0(N7952), .A1(N7584), .B0(N7829));
NAND2XL inst_cellmath__198_0_I2138 (.Y(N7516), .A(N7952), .B(N7711));
AOI21XL inst_cellmath__198_0_I2139 (.Y(N7645), .A0(N7882), .A1(N8082), .B0(N7761));
OAI21XL inst_cellmath__198_0_I2140 (.Y(N7572), .A0(N7743), .A1(N7931), .B0(N7610));
OAI21XL inst_cellmath__198_0_I2141 (.Y(N7818), .A0(N7669), .A1(N7860), .B0(N7538));
NOR2XL inst_cellmath__198_0_I2142 (.Y(N7940), .A(N7669), .B(N7984));
OAI21XL inst_cellmath__198_0_I2143 (.Y(N8067), .A0(N7592), .A1(N7787), .B0(N8036));
NOR2XL inst_cellmath__198_0_I2144 (.Y(N7620), .A(N7592), .B(N7913));
OAI21XL inst_cellmath__198_0_I2145 (.Y(N7751), .A0(N7516), .A1(N7720), .B0(N7963));
NOR2XL inst_cellmath__198_0_I2146 (.Y(N7869), .A(N7516), .B(N7839));
AOI21XL inst_cellmath__198_0_I2147 (.Y(N7995), .A0(N7940), .A1(N7572), .B0(N7818));
AOI21XL inst_cellmath__198_0_I2148 (.Y(N7676), .A0(N7869), .A1(N8067), .B0(N7751));
NAND2XL inst_cellmath__198_0_I2149 (.Y(N7797), .A(N7869), .B(N7620));
INVXL inst_cellmath__198_0_I2150 (.Y(N7919), .A(N7620));
INVXL inst_cellmath__198_0_I2151 (.Y(N8045), .A(N8067));
OAI21XL inst_cellmath__198_0_I2152 (.Y(N7600), .A0(N7919), .A1(N7995), .B0(N8045));
OAI21XL inst_cellmath__198_0_I2153 (.Y(N7846), .A0(N7797), .A1(N7995), .B0(N7676));
INVXL inst_cellmath__198_0_I2154 (.Y(N7526), .A(N7984));
INVXL inst_cellmath__198_0_I2155 (.Y(N7654), .A(N7860));
AOI21XL inst_cellmath__198_0_I2156 (.Y(N7776), .A0(N7526), .A1(N7572), .B0(N7654));
INVXL inst_cellmath__198_0_I2157 (.Y(N7562), .A(N7995));
OAI21XL inst_cellmath__198_0_I2158 (.Y(N7708), .A0(N7913), .A1(N7995), .B0(N7787));
INVXL inst_cellmath__198_0_I2159 (.Y(N7691), .A(N7600));
INVXL inst_cellmath__198_0_I2160 (.Y(N7633), .A(N7839));
INVXL inst_cellmath__198_0_I2161 (.Y(N7759), .A(N7720));
AOI21XL inst_cellmath__198_0_I2162 (.Y(N7880), .A0(N7633), .A1(N7600), .B0(N7759));
INVXL inst_cellmath__198_0_I2163 (.Y(N7810), .A(N7846));
INVXL inst_cellmath__198_0_I2164 (.Y(N7929), .A(N7645));
AOI31X1 inst_cellmath__198_0_I2165 (.Y(N8056), .A0(N7882), .A1(N7635), .A2(N7846), .B0(N7929));
AOI21XL inst_cellmath__198_0_I2169 (.Y(N7909), .A0(N8070), .A1(N7572), .B0(N7944));
INVXL inst_cellmath__198_0_I2170 (.Y(N7836), .A(N7997));
INVXL inst_cellmath__198_0_I2171 (.Y(N7960), .A(N7872));
OAI21XL inst_cellmath__198_0_I2172 (.Y(N8089), .A0(N7836), .A1(N7776), .B0(N7960));
AOI21XL inst_cellmath__198_0_I2173 (.Y(N8012), .A0(N7923), .A1(N7562), .B0(N7800));
AOI21XL inst_cellmath__198_0_I2174 (.Y(N7937), .A0(N7849), .A1(N7708), .B0(N7733));
INVXL inst_cellmath__198_0_I2175 (.Y(N7866), .A(N7778));
INVXL inst_cellmath__198_0_I2176 (.Y(N7991), .A(N7657));
OAI21XL inst_cellmath__198_0_I2177 (.Y(N7545), .A0(N7866), .A1(N7691), .B0(N7991));
INVXL inst_cellmath__198_0_I2178 (.Y(N8042), .A(N7711));
INVXL inst_cellmath__198_0_I2179 (.Y(N7597), .A(N7584));
OAI21XL inst_cellmath__198_0_I2180 (.Y(N7728), .A0(N8042), .A1(N7880), .B0(N7597));
INVXL inst_cellmath__198_0_I2181 (.Y(N7651), .A(N7635));
INVXL inst_cellmath__198_0_I2182 (.Y(N7773), .A(N8082));
OAI21XL inst_cellmath__198_0_I2183 (.Y(N7897), .A0(N7651), .A1(N7810), .B0(N7773));
OAI22XL inst_cellmath__198_0_I2184 (.Y(N8076), .A0(N7825), .A1(N8056), .B0(N7789), .B1(N7924));
XOR2XL inst_cellmath__198_0_I2189 (.Y(inst_cellmath__198[18]), .A(N7909), .B(N7753));
XOR2XL inst_cellmath__198_0_I2190 (.Y(inst_cellmath__198[19]), .A(N7776), .B(N7997));
XNOR2X1 inst_cellmath__198_0_I2191 (.Y(inst_cellmath__198[20]), .A(N8089), .B(N7679));
XNOR2X1 inst_cellmath__198_0_I2192 (.Y(inst_cellmath__198[21]), .A(N7562), .B(N7923));
XOR2XL inst_cellmath__198_0_I2193 (.Y(inst_cellmath__198[22]), .A(N8012), .B(N7602));
XNOR2X1 inst_cellmath__198_0_I2194 (.Y(inst_cellmath__198[23]), .A(N7708), .B(N7849));
XOR2XL inst_cellmath__198_0_I2195 (.Y(inst_cellmath__198[24]), .A(N7937), .B(N7529));
XOR2XL inst_cellmath__198_0_I2196 (.Y(inst_cellmath__198[25]), .A(N7691), .B(N7778));
XNOR2X1 inst_cellmath__198_0_I2197 (.Y(inst_cellmath__198[26]), .A(N7545), .B(N8025));
XOR2XL inst_cellmath__198_0_I2198 (.Y(inst_cellmath__198[27]), .A(N7880), .B(N7711));
XNOR2X1 inst_cellmath__198_0_I2199 (.Y(inst_cellmath__198[28]), .A(N7728), .B(N7952));
XOR2XL inst_cellmath__198_0_I2200 (.Y(inst_cellmath__198[29]), .A(N7810), .B(N7635));
XNOR2X1 inst_cellmath__198_0_I2201 (.Y(inst_cellmath__198[30]), .A(N7897), .B(N7882));
XNOR2X1 inst_cellmath__198_0_I2202 (.Y(inst_cellmath__198[31]), .A(N8056), .B(N7825));
XNOR2X1 inst_cellmath__198_0_I2203 (.Y(inst_cellmath__198[32]), .A(N8076), .B(N7807));
NOR3XL inst_cellmath__203_0_I8433 (.Y(N10310), .A(N6061), .B(N5958), .C(N6252));
NOR3BX1 inst_cellmath__203_0_I8491 (.Y(N8975), .AN(N6186), .B(N6296), .C(N6651));
NOR2BX1 inst_cellmath__203_0_I8435 (.Y(N9352), .AN(N6234), .B(N6045));
NOR3BX1 inst_cellmath__203_0_I8492 (.Y(N9745), .AN(N6282), .B(N6196), .C(N5903));
NOR4X1 inst_cellmath__203_0_I8437 (.Y(N10108), .A(N5955), .B(N6030), .C(N6139), .D(N6328));
NAND2XL hyperpropagate_3_1_A_I8517 (.Y(N19025), .A(N6535), .B(N6435));
NOR2XL hyperpropagate_3_1_A_I8518 (.Y(N8774), .A(N5884), .B(N19025));
NOR3BX1 inst_cellmath__203_0_I8493 (.Y(N9125), .AN(N6661), .B(N6121), .C(N6309));
NOR3BX1 inst_cellmath__203_0_I8494 (.Y(N9517), .AN(N5867), .B(N6519), .C(N6351));
NOR3BX1 inst_cellmath__203_0_I8495 (.Y(N9894), .AN(N6565), .B(N6026), .C(N6385));
NOR3BX1 inst_cellmath__203_0_I8496 (.Y(N10255), .AN(N6433), .B(N6532), .C(N6260));
NOR3BX1 inst_cellmath__203_0_I8497 (.Y(N8914), .AN(N6304), .B(N6114), .C(N5935));
NOR3BX1 inst_cellmath__203_0_I8498 (.Y(N9677), .AN(N6638), .B(N6098), .C(N6287));
AND2XL inst_cellmath__203_0_I8445 (.Y(N9064), .A(N6556), .B(N6457));
NOR4X1 inst_cellmath__203_0_I8446 (.Y(N9447), .A(N5872), .B(N6423), .C(N6060), .D(N6251));
NOR3BX1 inst_cellmath__203_0_I8499 (.Y(N9832), .AN(N6109), .B(N5924), .C(N6390));
NOR3BX1 inst_cellmath__203_0_I8500 (.Y(N10191), .AN(N6155), .B(N6617), .C(N5975));
NOR2BX1 inst_cellmath__203_0_I8449 (.Y(N8851), .AN(N6017), .B(N6482));
XOR2XL inst_cellmath__203_0_I8450 (.Y(N9219), .A(N7572), .B(N8070));
NOR2XL inst_cellmath__203_0_I2226 (.Y(N10277), .A(N9219), .B(N8975));
NOR2XL inst_cellmath__203_0_I2227 (.Y(N9311), .A(N9219), .B(N9352));
NOR2XL inst_cellmath__203_0_I2228 (.Y(N10069), .A(N9219), .B(N9745));
NOR2XL inst_cellmath__203_0_I2229 (.Y(N9084), .A(N9219), .B(N10108));
NOR2XL inst_cellmath__203_0_I2230 (.Y(N9859), .A(N9219), .B(N8774));
NOR2XL inst_cellmath__203_0_I2231 (.Y(N8874), .A(N9219), .B(N9125));
NOR2XL inst_cellmath__203_0_I2232 (.Y(N9635), .A(N9219), .B(N9517));
NOR2XL inst_cellmath__203_0_I2233 (.Y(N8691), .A(N9219), .B(N9894));
NOR2XL inst_cellmath__203_0_I2234 (.Y(N9405), .A(N9219), .B(N10255));
NOR2XL inst_cellmath__203_0_I2235 (.Y(N10152), .A(N9219), .B(N8914));
NOR2XL inst_cellmath__203_0_I2236 (.Y(N9177), .A(N9219), .B(N9284));
NOR2XL inst_cellmath__203_0_I2237 (.Y(N9949), .A(N9219), .B(N9677));
NOR2XL inst_cellmath__203_0_I2238 (.Y(N8960), .A(N9219), .B(N10044));
NOR2XL inst_cellmath__203_0_I2239 (.Y(N9734), .A(N9219), .B(N6236));
NOR2XL inst_cellmath__203_0_I2240 (.Y(N8763), .A(N9219), .B(N9064));
NOR2XL inst_cellmath__203_0_I2241 (.Y(N9501), .A(N9219), .B(N9447));
NOR2XL inst_cellmath__203_0_I2242 (.Y(N10245), .A(N9219), .B(N9832));
NOR2XL inst_cellmath__203_0_I2243 (.Y(N9272), .A(N9219), .B(N10191));
NOR2XL inst_cellmath__203_0_I2244 (.Y(N10034), .A(N9219), .B(N8851));
INVXL inst_cellmath__203_0_I2245 (.Y(N8669), .A(inst_cellmath__198[18]));
NAND2BX1 inst_cellmath__203_0_I2246 (.Y(N9001), .AN(inst_cellmath__198[19]), .B(inst_cellmath__198[18]));
INVXL inst_cellmath__203_0_I2247 (.Y(N9381), .A(inst_cellmath__198[19]));
NOR2XL inst_cellmath__203_0_I2248 (.Y(N9704), .A(N10310), .B(N8669));
MXI2XL inst_cellmath__203_0_I2249 (.Y(inst_cellmath__203__W0[1]), .A(N9381), .B(N9001), .S0(N9704));
MXI2XL inst_cellmath__203_0_I2250 (.Y(N9637), .A(N8975), .B(N10310), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2251 (.Y(N9366), .A(N9381), .B(N9001), .S0(N9637));
MXI2XL inst_cellmath__203_0_I2252 (.Y(N9570), .A(N9352), .B(N8975), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2253 (.Y(N9759), .A(N9381), .B(N9001), .S0(N9570));
MXI2XL inst_cellmath__203_0_I2254 (.Y(N9504), .A(N9745), .B(N9352), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2255 (.Y(N10122), .A(N9381), .B(N9001), .S0(N9504));
MXI2XL inst_cellmath__203_0_I2256 (.Y(N9436), .A(N10108), .B(N9745), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2257 (.Y(N8786), .A(N9381), .B(N9001), .S0(N9436));
MXI2XL inst_cellmath__203_0_I2258 (.Y(N9369), .A(N8774), .B(N10108), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2259 (.Y(N9139), .A(N9381), .B(N9001), .S0(N9369));
MXI2XL inst_cellmath__203_0_I2260 (.Y(N9304), .A(N9125), .B(N8774), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2261 (.Y(N9532), .A(N9381), .B(N9001), .S0(N9304));
MXI2XL inst_cellmath__203_0_I2262 (.Y(N9240), .A(N9517), .B(N9125), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2263 (.Y(N9912), .A(N9381), .B(N9001), .S0(N9240));
MXI2XL inst_cellmath__203_0_I2264 (.Y(N9170), .A(N9894), .B(N9517), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2265 (.Y(N10268), .A(N9381), .B(N9001), .S0(N9170));
MXI2XL inst_cellmath__203_0_I2266 (.Y(N9104), .A(N10255), .B(N9894), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2267 (.Y(N8928), .A(N9381), .B(N9001), .S0(N9104));
MXI2XL inst_cellmath__203_0_I2268 (.Y(N9046), .A(N8914), .B(N10255), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2269 (.Y(N9300), .A(N9381), .B(N9001), .S0(N9046));
MXI2XL inst_cellmath__203_0_I2270 (.Y(N8983), .A(N9284), .B(N8914), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2271 (.Y(N9694), .A(N9381), .B(N9001), .S0(N8983));
MXI2XL inst_cellmath__203_0_I2272 (.Y(N8923), .A(N9677), .B(N9284), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2273 (.Y(N10060), .A(N9381), .B(N9001), .S0(N8923));
MXI2XL inst_cellmath__203_0_I2274 (.Y(N8862), .A(N10044), .B(N9677), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2275 (.Y(N8736), .A(N9381), .B(N9001), .S0(N8862));
MXI2XL inst_cellmath__203_0_I2276 (.Y(N8805), .A(N6236), .B(N10044), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2277 (.Y(N9076), .A(N9381), .B(N9001), .S0(N8805));
MXI2XL inst_cellmath__203_0_I2278 (.Y(N8751), .A(N9064), .B(N6236), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2279 (.Y(N9464), .A(N9381), .B(N9001), .S0(N8751));
MXI2XL inst_cellmath__203_0_I2280 (.Y(N8704), .A(N9447), .B(N9064), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2281 (.Y(N9851), .A(N9381), .B(N9001), .S0(N8704));
MXI2XL inst_cellmath__203_0_I2282 (.Y(N8651), .A(N9832), .B(N9447), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2283 (.Y(N10207), .A(N9381), .B(N9001), .S0(N8651));
MXI2XL inst_cellmath__203_0_I2284 (.Y(N10259), .A(N10191), .B(N9832), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2285 (.Y(N8868), .A(N9381), .B(N9001), .S0(N10259));
MXI2XL inst_cellmath__203_0_I2286 (.Y(N10196), .A(N8851), .B(N10191), .S0(N8669));
MXI2XL inst_cellmath__203_0_I2287 (.Y(N9236), .A(N9381), .B(N9001), .S0(N10196));
NAND2XL inst_cellmath__203_0_I2288 (.Y(N10133), .A(N8851), .B(N8669));
MXI2XL inst_cellmath__203_0_I2289 (.Y(N9628), .A(N9381), .B(N9001), .S0(N10133));
XNOR2X1 inst_cellmath__203_0_I2290 (.Y(N9402), .A(inst_cellmath__198[20]), .B(inst_cellmath__198[19]));
NOR2XL inst_cellmath__203_0_I2291 (.Y(N9092), .A(inst_cellmath__198[20]), .B(inst_cellmath__198[19]));
OAI2BB1X1 inst_cellmath__203_0_I2292 (.Y(N9017), .A0N(inst_cellmath__198[20]), .A1N(inst_cellmath__198[19]), .B0(inst_cellmath__198[21]));
INVXL inst_cellmath__203_0_I2293 (.Y(N9768), .A(N9017));
OR2XL inst_cellmath__203_0_I2294 (.Y(N9153), .A(N9092), .B(inst_cellmath__198[21]));
INVXL inst_cellmath__203_0_I2295 (.Y(N9545), .A(N9768));
NOR2XL inst_cellmath__203_0_I2296 (.Y(N9801), .A(N10310), .B(N9402));
MXI2XL inst_cellmath__203_0_I2297 (.Y(N9942), .A(N9545), .B(N9153), .S0(N9801));
MXI2XL inst_cellmath__203_0_I2298 (.Y(N9741), .A(N8975), .B(N10310), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2299 (.Y(N10292), .A(N9545), .B(N9153), .S0(N9741));
MXI2XL inst_cellmath__203_0_I2300 (.Y(N9673), .A(N9352), .B(N8975), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2301 (.Y(N8952), .A(N9545), .B(N9153), .S0(N9673));
MXI2XL inst_cellmath__203_0_I2302 (.Y(N9606), .A(N9745), .B(N9352), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2303 (.Y(N9334), .A(N9545), .B(N9153), .S0(N9606));
MXI2XL inst_cellmath__203_0_I2304 (.Y(N9542), .A(N10108), .B(N9745), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2305 (.Y(N9725), .A(N9545), .B(N9153), .S0(N9542));
MXI2XL inst_cellmath__203_0_I2306 (.Y(N9471), .A(N8774), .B(N10108), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2307 (.Y(N10088), .A(N9545), .B(N9153), .S0(N9471));
MXI2XL inst_cellmath__203_0_I2308 (.Y(N9406), .A(N9125), .B(N8774), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2309 (.Y(N8757), .A(N9545), .B(N9153), .S0(N9406));
MXI2XL inst_cellmath__203_0_I2310 (.Y(N9339), .A(N9517), .B(N9125), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2311 (.Y(N9103), .A(N9545), .B(N9153), .S0(N9339));
MXI2XL inst_cellmath__203_0_I2312 (.Y(N9273), .A(N9894), .B(N9517), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2313 (.Y(N9494), .A(N9545), .B(N9153), .S0(N9273));
MXI2XL inst_cellmath__203_0_I2314 (.Y(N9204), .A(N10255), .B(N9894), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2315 (.Y(N9879), .A(N9545), .B(N9153), .S0(N9204));
MXI2XL inst_cellmath__203_0_I2316 (.Y(N9140), .A(N8914), .B(N10255), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2317 (.Y(N10236), .A(N9545), .B(N9153), .S0(N9140));
MXI2XL inst_cellmath__203_0_I2318 (.Y(N9077), .A(N9284), .B(N8914), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2319 (.Y(N8893), .A(N9545), .B(N9153), .S0(N9077));
MXI2XL inst_cellmath__203_0_I2320 (.Y(N9018), .A(N9677), .B(N9284), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2321 (.Y(N9267), .A(N9545), .B(N9153), .S0(N9018));
MXI2XL inst_cellmath__203_0_I2322 (.Y(N8953), .A(N10044), .B(N9677), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2323 (.Y(N9661), .A(N9545), .B(N9153), .S0(N8953));
MXI2XL inst_cellmath__203_0_I2324 (.Y(N8894), .A(N6236), .B(N10044), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2325 (.Y(N10025), .A(N9545), .B(N9153), .S0(N8894));
MXI2XL inst_cellmath__203_0_I2326 (.Y(N8834), .A(N9064), .B(N6236), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2327 (.Y(N8709), .A(N9545), .B(N9153), .S0(N8834));
MXI2XL inst_cellmath__203_0_I2328 (.Y(N8781), .A(N9447), .B(N9064), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2329 (.Y(N9045), .A(N9545), .B(N9153), .S0(N8781));
MXI2XL inst_cellmath__203_0_I2330 (.Y(N8730), .A(N9832), .B(N9447), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2331 (.Y(N9427), .A(N9545), .B(N9153), .S0(N8730));
MXI2XL inst_cellmath__203_0_I2332 (.Y(N8677), .A(N10191), .B(N9832), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2333 (.Y(N9815), .A(N9545), .B(N9153), .S0(N8677));
MXI2XL inst_cellmath__203_0_I2334 (.Y(N10285), .A(N8851), .B(N10191), .S0(N9402));
MXI2XL inst_cellmath__203_0_I2335 (.Y(N10172), .A(N9545), .B(N9153), .S0(N10285));
NAND2XL inst_cellmath__203_0_I2336 (.Y(N10228), .A(N8851), .B(N9402));
MXI2XL inst_cellmath__203_0_I2337 (.Y(N8833), .A(N9545), .B(N9153), .S0(N10228));
XNOR2X1 inst_cellmath__203_0_I2338 (.Y(N8655), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
NOR2XL inst_cellmath__203_0_I2339 (.Y(N9193), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
OAI2BB1X1 inst_cellmath__203_0_I2340 (.Y(N9966), .A0N(inst_cellmath__198[22]), .A1N(inst_cellmath__198[21]), .B0(inst_cellmath__198[23]));
INVXL inst_cellmath__203_0_I2341 (.Y(N9925), .A(N9966));
OR2XL inst_cellmath__203_0_I2342 (.Y(N9317), .A(N9193), .B(inst_cellmath__198[23]));
INVXL inst_cellmath__203_0_I2343 (.Y(N9706), .A(N9925));
NOR2XL inst_cellmath__203_0_I2344 (.Y(N9895), .A(N10310), .B(N8655));
MXI2XL inst_cellmath__203_0_I2345 (.Y(N9133), .A(N9706), .B(N9317), .S0(N9895));
MXI2XL inst_cellmath__203_0_I2346 (.Y(N9834), .A(N8975), .B(N10310), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2347 (.Y(N9527), .A(N9706), .B(N9317), .S0(N9834));
MXI2XL inst_cellmath__203_0_I2348 (.Y(N9770), .A(N9352), .B(N8975), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2349 (.Y(N9903), .A(N9706), .B(N9317), .S0(N9770));
MXI2XL inst_cellmath__203_0_I2350 (.Y(N9708), .A(N9745), .B(N9352), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2351 (.Y(N10262), .A(N9706), .B(N9317), .S0(N9708));
MXI2XL inst_cellmath__203_0_I2352 (.Y(N9641), .A(N10108), .B(N9745), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2353 (.Y(N8921), .A(N9706), .B(N9317), .S0(N9641));
MXI2XL inst_cellmath__203_0_I2354 (.Y(N9573), .A(N8774), .B(N10108), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2355 (.Y(N9293), .A(N9706), .B(N9317), .S0(N9573));
MXI2XL inst_cellmath__203_0_I2356 (.Y(N9508), .A(N9125), .B(N8774), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2357 (.Y(N9686), .A(N9706), .B(N9317), .S0(N9508));
MXI2XL inst_cellmath__203_0_I2358 (.Y(N9439), .A(N9517), .B(N9125), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2359 (.Y(N10052), .A(N9706), .B(N9317), .S0(N9439));
MXI2XL inst_cellmath__203_0_I2360 (.Y(N9372), .A(N9894), .B(N9517), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2361 (.Y(N8729), .A(N9706), .B(N9317), .S0(N9372));
MXI2XL inst_cellmath__203_0_I2362 (.Y(N9310), .A(N10255), .B(N9894), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2363 (.Y(N9071), .A(N9706), .B(N9317), .S0(N9310));
MXI2XL inst_cellmath__203_0_I2364 (.Y(N9244), .A(N8914), .B(N10255), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2365 (.Y(N9458), .A(N9706), .B(N9317), .S0(N9244));
MXI2XL inst_cellmath__203_0_I2366 (.Y(N9174), .A(N9284), .B(N8914), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2367 (.Y(N9842), .A(N9706), .B(N9317), .S0(N9174));
MXI2XL inst_cellmath__203_0_I2368 (.Y(N9109), .A(N9677), .B(N9284), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2369 (.Y(N10200), .A(N9706), .B(N9317), .S0(N9109));
MXI2XL inst_cellmath__203_0_I2370 (.Y(N9050), .A(N10044), .B(N9677), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2371 (.Y(N8860), .A(N9706), .B(N9317), .S0(N9050));
MXI2XL inst_cellmath__203_0_I2372 (.Y(N8987), .A(N6236), .B(N10044), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2373 (.Y(N9228), .A(N9706), .B(N9317), .S0(N8987));
MXI2XL inst_cellmath__203_0_I2374 (.Y(N8926), .A(N9064), .B(N6236), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2375 (.Y(N9619), .A(N9706), .B(N9317), .S0(N8926));
MXI2XL inst_cellmath__203_0_I2376 (.Y(N8865), .A(N9447), .B(N9064), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2377 (.Y(N9992), .A(N9706), .B(N9317), .S0(N8865));
MXI2XL inst_cellmath__203_0_I2378 (.Y(N8809), .A(N9832), .B(N9447), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2379 (.Y(N8676), .A(N9706), .B(N9317), .S0(N8809));
MXI2XL inst_cellmath__203_0_I2380 (.Y(N8755), .A(N10191), .B(N9832), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2381 (.Y(N9011), .A(N9706), .B(N9317), .S0(N8755));
MXI2XL inst_cellmath__203_0_I2382 (.Y(N8707), .A(N8851), .B(N10191), .S0(N8655));
MXI2XL inst_cellmath__203_0_I2383 (.Y(N9393), .A(N9706), .B(N9317), .S0(N8707));
NAND2XL inst_cellmath__203_0_I2384 (.Y(N8654), .A(N8851), .B(N8655));
MXI2XL inst_cellmath__203_0_I2385 (.Y(N9778), .A(N9706), .B(N9317), .S0(N8654));
XNOR2X1 inst_cellmath__203_0_I2386 (.Y(N9555), .A(inst_cellmath__198[24]), .B(inst_cellmath__198[23]));
NOR2XL inst_cellmath__203_0_I2387 (.Y(N9291), .A(inst_cellmath__198[24]), .B(inst_cellmath__198[23]));
OAI2BB1X1 inst_cellmath__203_0_I2388 (.Y(N9161), .A0N(inst_cellmath__198[24]), .A1N(inst_cellmath__198[23]), .B0(inst_cellmath__198[25]));
INVXL inst_cellmath__203_0_I2389 (.Y(N10071), .A(N9161));
OR2XL inst_cellmath__203_0_I2390 (.Y(N9475), .A(N9291), .B(inst_cellmath__198[25]));
INVXL inst_cellmath__203_0_I2391 (.Y(N9861), .A(N10071));
NOR2XL inst_cellmath__203_0_I2392 (.Y(N9989), .A(N10310), .B(N9555));
MXI2XL inst_cellmath__203_0_I2393 (.Y(N10078), .A(N9861), .B(N9475), .S0(N9989));
MXI2XL inst_cellmath__203_0_I2394 (.Y(N9931), .A(N8975), .B(N10310), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2395 (.Y(N8749), .A(N9861), .B(N9475), .S0(N9931));
MXI2XL inst_cellmath__203_0_I2396 (.Y(N9868), .A(N9352), .B(N8975), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2397 (.Y(N9097), .A(N9861), .B(N9475), .S0(N9868));
MXI2XL inst_cellmath__203_0_I2398 (.Y(N9804), .A(N9745), .B(N9352), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2399 (.Y(N9485), .A(N9861), .B(N9475), .S0(N9804));
MXI2XL inst_cellmath__203_0_I2400 (.Y(N9744), .A(N10108), .B(N9745), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2401 (.Y(N9870), .A(N9861), .B(N9475), .S0(N9744));
MXI2XL inst_cellmath__203_0_I2402 (.Y(N9676), .A(N8774), .B(N10108), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2403 (.Y(N10227), .A(N9861), .B(N9475), .S0(N9676));
MXI2XL inst_cellmath__203_0_I2404 (.Y(N9608), .A(N9125), .B(N8774), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2405 (.Y(N8886), .A(N9861), .B(N9475), .S0(N9608));
MXI2XL inst_cellmath__203_0_I2406 (.Y(N9544), .A(N9517), .B(N9125), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2407 (.Y(N9258), .A(N9861), .B(N9475), .S0(N9544));
MXI2XL inst_cellmath__203_0_I2408 (.Y(N9474), .A(N9894), .B(N9517), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2409 (.Y(N9649), .A(N9861), .B(N9475), .S0(N9474));
MXI2XL inst_cellmath__203_0_I2410 (.Y(N9409), .A(N10255), .B(N9894), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2411 (.Y(N10016), .A(N9861), .B(N9475), .S0(N9409));
MXI2XL inst_cellmath__203_0_I2412 (.Y(N9342), .A(N8914), .B(N10255), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2413 (.Y(N8700), .A(N9861), .B(N9475), .S0(N9342));
MXI2XL inst_cellmath__203_0_I2414 (.Y(N9275), .A(N9284), .B(N8914), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2415 (.Y(N9036), .A(N9861), .B(N9475), .S0(N9275));
MXI2XL inst_cellmath__203_0_I2416 (.Y(N9206), .A(N9677), .B(N9284), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2417 (.Y(N9419), .A(N9861), .B(N9475), .S0(N9206));
MXI2XL inst_cellmath__203_0_I2418 (.Y(N9142), .A(N10044), .B(N9677), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2419 (.Y(N9805), .A(N9861), .B(N9475), .S0(N9142));
MXI2XL inst_cellmath__203_0_I2420 (.Y(N9080), .A(N6236), .B(N10044), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2421 (.Y(N10164), .A(N9861), .B(N9475), .S0(N9080));
MXI2XL inst_cellmath__203_0_I2422 (.Y(N9021), .A(N9064), .B(N6236), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2423 (.Y(N8827), .A(N9861), .B(N9475), .S0(N9021));
MXI2XL inst_cellmath__203_0_I2424 (.Y(N8954), .A(N9447), .B(N9064), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2425 (.Y(N9192), .A(N9861), .B(N9475), .S0(N8954));
MXI2XL inst_cellmath__203_0_I2426 (.Y(N8898), .A(N9832), .B(N9447), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2427 (.Y(N9581), .A(N9861), .B(N9475), .S0(N8898));
MXI2XL inst_cellmath__203_0_I2428 (.Y(N8837), .A(N10191), .B(N9832), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2429 (.Y(N9959), .A(N9861), .B(N9475), .S0(N8837));
MXI2XL inst_cellmath__203_0_I2430 (.Y(N8782), .A(N8851), .B(N10191), .S0(N9555));
MXI2XL inst_cellmath__203_0_I2431 (.Y(N8649), .A(N9861), .B(N9475), .S0(N8782));
NAND2XL inst_cellmath__203_0_I2432 (.Y(N8734), .A(N8851), .B(N9555));
MXI2XL inst_cellmath__203_0_I2433 (.Y(N8976), .A(N9861), .B(N9475), .S0(N8734));
XNOR2X1 inst_cellmath__203_0_I2434 (.Y(N8775), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
NOR2XL inst_cellmath__203_0_I2435 (.Y(N9396), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
OAI2BB1X1 inst_cellmath__203_0_I2436 (.Y(N10110), .A0N(inst_cellmath__198[26]), .A1N(inst_cellmath__198[25]), .B0(inst_cellmath__198[27]));
INVXL inst_cellmath__203_0_I2437 (.Y(N10219), .A(N10110));
OR2XL inst_cellmath__203_0_I2438 (.Y(N9639), .A(N9396), .B(inst_cellmath__198[27]));
INVXL inst_cellmath__203_0_I2439 (.Y(N10009), .A(N10219));
NOR2XL inst_cellmath__203_0_I2440 (.Y(N10081), .A(N10310), .B(N8775));
MXI2XL inst_cellmath__203_0_I2441 (.Y(N9285), .A(N10009), .B(N9639), .S0(N10081));
MXI2XL inst_cellmath__203_0_I2442 (.Y(N10020), .A(N8975), .B(N10310), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2443 (.Y(N9678), .A(N10009), .B(N9639), .S0(N10020));
MXI2XL inst_cellmath__203_0_I2444 (.Y(N9961), .A(N9352), .B(N8975), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2445 (.Y(N10046), .A(N10009), .B(N9639), .S0(N9961));
MXI2XL inst_cellmath__203_0_I2446 (.Y(N9898), .A(N9745), .B(N9352), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2447 (.Y(N8725), .A(N10009), .B(N9639), .S0(N9898));
MXI2XL inst_cellmath__203_0_I2448 (.Y(N9837), .A(N10108), .B(N9745), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2449 (.Y(N9066), .A(N10009), .B(N9639), .S0(N9837));
MXI2XL inst_cellmath__203_0_I2450 (.Y(N9772), .A(N8774), .B(N10108), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2451 (.Y(N9448), .A(N10009), .B(N9639), .S0(N9772));
MXI2XL inst_cellmath__203_0_I2452 (.Y(N9712), .A(N9125), .B(N8774), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2453 (.Y(N9833), .A(N10009), .B(N9639), .S0(N9712));
MXI2XL inst_cellmath__203_0_I2454 (.Y(N9645), .A(N9517), .B(N9125), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2455 (.Y(N10193), .A(N10009), .B(N9639), .S0(N9645));
MXI2XL inst_cellmath__203_0_I2456 (.Y(N9577), .A(N9894), .B(N9517), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2457 (.Y(N8853), .A(N10009), .B(N9639), .S0(N9577));
MXI2XL inst_cellmath__203_0_I2458 (.Y(N9513), .A(N10255), .B(N9894), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2459 (.Y(N9220), .A(N10009), .B(N9639), .S0(N9513));
MXI2XL inst_cellmath__203_0_I2460 (.Y(N9443), .A(N8914), .B(N10255), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2461 (.Y(N9609), .A(N10009), .B(N9639), .S0(N9443));
MXI2XL inst_cellmath__203_0_I2462 (.Y(N9378), .A(N9284), .B(N8914), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2463 (.Y(N9984), .A(N10009), .B(N9639), .S0(N9378));
MXI2XL inst_cellmath__203_0_I2464 (.Y(N9314), .A(N9677), .B(N9284), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2465 (.Y(N8670), .A(N10009), .B(N9639), .S0(N9314));
MXI2XL inst_cellmath__203_0_I2466 (.Y(N9246), .A(N10044), .B(N9677), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2467 (.Y(N9003), .A(N10009), .B(N9639), .S0(N9246));
MXI2XL inst_cellmath__203_0_I2468 (.Y(N9178), .A(N6236), .B(N10044), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2469 (.Y(N9383), .A(N10009), .B(N9639), .S0(N9178));
MXI2XL inst_cellmath__203_0_I2470 (.Y(N9112), .A(N9064), .B(N6236), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2471 (.Y(N9769), .A(N10009), .B(N9639), .S0(N9112));
MXI2XL inst_cellmath__203_0_I2472 (.Y(N9053), .A(N9447), .B(N9064), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2473 (.Y(N10131), .A(N10009), .B(N9639), .S0(N9053));
MXI2XL inst_cellmath__203_0_I2474 (.Y(N8990), .A(N9832), .B(N9447), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2475 (.Y(N8797), .A(N10009), .B(N9639), .S0(N8990));
MXI2XL inst_cellmath__203_0_I2476 (.Y(N8929), .A(N10191), .B(N9832), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2477 (.Y(N9154), .A(N10009), .B(N9639), .S0(N8929));
MXI2XL inst_cellmath__203_0_I2478 (.Y(N8869), .A(N8851), .B(N10191), .S0(N8775));
MXI2XL inst_cellmath__203_0_I2479 (.Y(N9547), .A(N10009), .B(N9639), .S0(N8869));
NAND2XL inst_cellmath__203_0_I2480 (.Y(N8811), .A(N8851), .B(N8775));
MXI2XL inst_cellmath__203_0_I2481 (.Y(N9927), .A(N10009), .B(N9639), .S0(N8811));
XNOR2X1 inst_cellmath__203_0_I2482 (.Y(N9707), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
NOR2XL inst_cellmath__203_0_I2483 (.Y(N9495), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
OAI2BB1X1 inst_cellmath__203_0_I2484 (.Y(N9319), .A0N(inst_cellmath__198[28]), .A1N(inst_cellmath__198[27]), .B0(inst_cellmath__198[29]));
INVXL inst_cellmath__203_0_I2485 (.Y(N8693), .A(N9319));
OR2XL inst_cellmath__203_0_I2486 (.Y(N9795), .A(N9495), .B(inst_cellmath__198[29]));
INVXL inst_cellmath__203_0_I2487 (.Y(N10157), .A(N8693));
NOR2XL inst_cellmath__203_0_I2488 (.Y(N10173), .A(N10310), .B(N9707));
MXI2XL inst_cellmath__203_0_I2489 (.Y(N10220), .A(N10157), .B(N9795), .S0(N10173));
MXI2XL inst_cellmath__203_0_I2490 (.Y(N10115), .A(N8975), .B(N10310), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2491 (.Y(N8879), .A(N10157), .B(N9795), .S0(N10115));
MXI2XL inst_cellmath__203_0_I2492 (.Y(N10053), .A(N9352), .B(N8975), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2493 (.Y(N9249), .A(N10157), .B(N9795), .S0(N10053));
MXI2XL inst_cellmath__203_0_I2494 (.Y(N9993), .A(N9745), .B(N9352), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2495 (.Y(N9640), .A(N10157), .B(N9795), .S0(N9993));
MXI2XL inst_cellmath__203_0_I2496 (.Y(N9932), .A(N10108), .B(N9745), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2497 (.Y(N10010), .A(N10157), .B(N9795), .S0(N9932));
MXI2XL inst_cellmath__203_0_I2498 (.Y(N9871), .A(N8774), .B(N10108), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2499 (.Y(N8695), .A(N10157), .B(N9795), .S0(N9871));
MXI2XL inst_cellmath__203_0_I2500 (.Y(N9806), .A(N9125), .B(N8774), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2501 (.Y(N9029), .A(N10157), .B(N9795), .S0(N9806));
MXI2XL inst_cellmath__203_0_I2502 (.Y(N9747), .A(N9517), .B(N9125), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2503 (.Y(N9411), .A(N10157), .B(N9795), .S0(N9747));
MXI2XL inst_cellmath__203_0_I2504 (.Y(N9679), .A(N9894), .B(N9517), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2505 (.Y(N9798), .A(N10157), .B(N9795), .S0(N9679));
MXI2XL inst_cellmath__203_0_I2506 (.Y(N9610), .A(N10255), .B(N9894), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2507 (.Y(N10158), .A(N10157), .B(N9795), .S0(N9610));
MXI2XL inst_cellmath__203_0_I2508 (.Y(N9548), .A(N8914), .B(N10255), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2509 (.Y(N8820), .A(N10157), .B(N9795), .S0(N9548));
MXI2XL inst_cellmath__203_0_I2510 (.Y(N9477), .A(N9284), .B(N8914), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2511 (.Y(N9183), .A(N10157), .B(N9795), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2512 (.Y(N9412), .A(N9677), .B(N9284), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2513 (.Y(N9572), .A(N10157), .B(N9795), .S0(N9412));
MXI2XL inst_cellmath__203_0_I2514 (.Y(N9346), .A(N10044), .B(N9677), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2515 (.Y(N9953), .A(N10157), .B(N9795), .S0(N9346));
MXI2XL inst_cellmath__203_0_I2516 (.Y(N9278), .A(N6236), .B(N10044), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2517 (.Y(N10305), .A(N10157), .B(N9795), .S0(N9278));
MXI2XL inst_cellmath__203_0_I2518 (.Y(N9211), .A(N9064), .B(N6236), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2519 (.Y(N8966), .A(N10157), .B(N9795), .S0(N9211));
MXI2XL inst_cellmath__203_0_I2520 (.Y(N9146), .A(N9447), .B(N9064), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2521 (.Y(N9345), .A(N10157), .B(N9795), .S0(N9146));
MXI2XL inst_cellmath__203_0_I2522 (.Y(N9082), .A(N9832), .B(N9447), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2523 (.Y(N9738), .A(N10157), .B(N9795), .S0(N9082));
MXI2XL inst_cellmath__203_0_I2524 (.Y(N9023), .A(N10191), .B(N9832), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2525 (.Y(N10102), .A(N10157), .B(N9795), .S0(N9023));
MXI2XL inst_cellmath__203_0_I2526 (.Y(N8959), .A(N8851), .B(N10191), .S0(N9707));
MXI2XL inst_cellmath__203_0_I2527 (.Y(N8768), .A(N10157), .B(N9795), .S0(N8959));
NAND2XL inst_cellmath__203_0_I2528 (.Y(N8902), .A(N8851), .B(N9707));
MXI2XL inst_cellmath__203_0_I2529 (.Y(N9118), .A(N10157), .B(N9795), .S0(N8902));
XNOR2X1 inst_cellmath__203_0_I2530 (.Y(N8908), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
NOR2XL inst_cellmath__203_0_I2531 (.Y(N9596), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
OAI2BB1X1 inst_cellmath__203_0_I2532 (.Y(N10251), .A0N(inst_cellmath__198[30]), .A1N(inst_cellmath__198[29]), .B0(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I2533 (.Y(N8817), .A(N10251));
OR2XL inst_cellmath__203_0_I2534 (.Y(N9952), .A(N9596), .B(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I2535 (.Y(N10302), .A(N8817));
NOR2XL inst_cellmath__203_0_I2536 (.Y(N10266), .A(N10310), .B(N8908));
MXI2XL inst_cellmath__203_0_I2537 (.Y(N9438), .A(N10302), .B(N9952), .S0(N10266));
MXI2XL inst_cellmath__203_0_I2538 (.Y(N10205), .A(N8975), .B(N10310), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2539 (.Y(N9827), .A(N10302), .B(N9952), .S0(N10205));
MXI2XL inst_cellmath__203_0_I2540 (.Y(N10142), .A(N9352), .B(N8975), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2541 (.Y(N10187), .A(N10302), .B(N9952), .S0(N10142));
MXI2XL inst_cellmath__203_0_I2542 (.Y(N10086), .A(N9745), .B(N9352), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2543 (.Y(N8843), .A(N10302), .B(N9952), .S0(N10086));
MXI2XL inst_cellmath__203_0_I2544 (.Y(N10024), .A(N10108), .B(N9745), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2545 (.Y(N9210), .A(N10302), .B(N9952), .S0(N10024));
MXI2XL inst_cellmath__203_0_I2546 (.Y(N9965), .A(N8774), .B(N10108), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2547 (.Y(N9603), .A(N10302), .B(N9952), .S0(N9965));
MXI2XL inst_cellmath__203_0_I2548 (.Y(N9902), .A(N9125), .B(N8774), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2549 (.Y(N9979), .A(N10302), .B(N9952), .S0(N9902));
MXI2XL inst_cellmath__203_0_I2550 (.Y(N9841), .A(N9517), .B(N9125), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2551 (.Y(N8665), .A(N10302), .B(N9952), .S0(N9841));
MXI2XL inst_cellmath__203_0_I2552 (.Y(N9777), .A(N9894), .B(N9517), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2553 (.Y(N8996), .A(N10302), .B(N9952), .S0(N9777));
MXI2XL inst_cellmath__203_0_I2554 (.Y(N9715), .A(N10255), .B(N9894), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2555 (.Y(N9375), .A(N10302), .B(N9952), .S0(N9715));
MXI2XL inst_cellmath__203_0_I2556 (.Y(N9648), .A(N8914), .B(N10255), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2557 (.Y(N9762), .A(N10302), .B(N9952), .S0(N9648));
MXI2XL inst_cellmath__203_0_I2558 (.Y(N9580), .A(N9284), .B(N8914), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2559 (.Y(N10128), .A(N10302), .B(N9952), .S0(N9580));
MXI2XL inst_cellmath__203_0_I2560 (.Y(N9516), .A(N9677), .B(N9284), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2561 (.Y(N8792), .A(N10302), .B(N9952), .S0(N9516));
MXI2XL inst_cellmath__203_0_I2562 (.Y(N9446), .A(N10044), .B(N9677), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2563 (.Y(N9145), .A(N10302), .B(N9952), .S0(N9446));
MXI2XL inst_cellmath__203_0_I2564 (.Y(N9380), .A(N6236), .B(N10044), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2565 (.Y(N9537), .A(N10302), .B(N9952), .S0(N9380));
MXI2XL inst_cellmath__203_0_I2566 (.Y(N9316), .A(N9064), .B(N6236), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2567 (.Y(N9921), .A(N10302), .B(N9952), .S0(N9316));
MXI2XL inst_cellmath__203_0_I2568 (.Y(N9248), .A(N9447), .B(N9064), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2569 (.Y(N10273), .A(N10302), .B(N9952), .S0(N9248));
MXI2XL inst_cellmath__203_0_I2570 (.Y(N9180), .A(N9832), .B(N9447), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2571 (.Y(N8933), .A(N10302), .B(N9952), .S0(N9180));
MXI2XL inst_cellmath__203_0_I2572 (.Y(N9114), .A(N10191), .B(N9832), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2573 (.Y(N9309), .A(N10302), .B(N9952), .S0(N9114));
MXI2XL inst_cellmath__203_0_I2574 (.Y(N9054), .A(N8851), .B(N10191), .S0(N8908));
MXI2XL inst_cellmath__203_0_I2575 (.Y(N9699), .A(N10302), .B(N9952), .S0(N9054));
NAND2XL inst_cellmath__203_0_I2576 (.Y(N8992), .A(N8851), .B(N8908));
MXI2XL inst_cellmath__203_0_I2577 (.Y(N10067), .A(N10302), .B(N9952), .S0(N8992));
ADDHX1 inst_cellmath__203_0_I2578 (.CO(N10214), .S(N9468), .A(inst_cellmath__198[32]), .B(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I2579 (.Y(N8965), .A(N9468));
INVXL inst_cellmath__203_0_I2580 (.Y(N9343), .A(N10214));
NOR2XL inst_cellmath__203_0_I2581 (.Y(N10149), .A(N8965), .B(N10310));
OAI22XL inst_cellmath__203_0_I2582 (.Y(N9173), .A0(N10310), .A1(N9343), .B0(N8965), .B1(N8975));
OAI22XL inst_cellmath__203_0_I2583 (.Y(N9947), .A0(N8975), .A1(N9343), .B0(N8965), .B1(N9352));
OAI22XL inst_cellmath__203_0_I2584 (.Y(N8957), .A0(N9352), .A1(N9343), .B0(N8965), .B1(N9745));
OAI22XL inst_cellmath__203_0_I2585 (.Y(N9731), .A0(N9745), .A1(N9343), .B0(N8965), .B1(N10108));
OAI22XL inst_cellmath__203_0_I2586 (.Y(N8761), .A0(N10108), .A1(N9343), .B0(N8965), .B1(N8774));
OAI22XL inst_cellmath__203_0_I2587 (.Y(N9498), .A0(N8774), .A1(N9343), .B0(N8965), .B1(N9125));
OAI22XL inst_cellmath__203_0_I2588 (.Y(N10241), .A0(N9125), .A1(N9343), .B0(N8965), .B1(N9517));
OAI22XL inst_cellmath__203_0_I2589 (.Y(N9270), .A0(N9517), .A1(N9343), .B0(N8965), .B1(N9894));
OAI22XL inst_cellmath__203_0_I2590 (.Y(N10031), .A0(N9894), .A1(N9343), .B0(N8965), .B1(N10255));
OAI22XL inst_cellmath__203_0_I2591 (.Y(N9049), .A0(N10255), .A1(N9343), .B0(N8965), .B1(N8914));
OAI22XL inst_cellmath__203_0_I2592 (.Y(N9821), .A0(N8914), .A1(N9343), .B0(N8965), .B1(N9284));
OAI22XL inst_cellmath__203_0_I2593 (.Y(N8839), .A0(N9284), .A1(N9343), .B0(N8965), .B1(N9677));
OAI22XL inst_cellmath__203_0_I2594 (.Y(N9595), .A0(N9677), .A1(N9343), .B0(N8965), .B1(N10044));
OAI22XL inst_cellmath__203_0_I2595 (.Y(N8659), .A0(N10044), .A1(N9343), .B0(N8965), .B1(N6236));
OAI22XL inst_cellmath__203_0_I2596 (.Y(N9363), .A0(N6236), .A1(N9343), .B0(N8965), .B1(N9064));
OAI22XL inst_cellmath__203_0_I2597 (.Y(N10118), .A0(N9064), .A1(N9343), .B0(N8965), .B1(N9447));
OAI22XL inst_cellmath__203_0_I2598 (.Y(N9137), .A0(N9447), .A1(N9343), .B0(N8965), .B1(N9832));
OAI22XL inst_cellmath__203_0_I2599 (.Y(N9909), .A0(N9832), .A1(N9343), .B0(N8965), .B1(N10191));
OAI22XL inst_cellmath__203_0_I2600 (.Y(N8925), .A0(N10191), .A1(N9343), .B0(N8965), .B1(N8851));
OAI21XL inst_cellmath__203_0_I2601 (.Y(N9692), .A0(N9343), .A1(N8851), .B0(N8965));
AND2XL inst_cellmath__203_0_I2602 (.Y(N10192), .A(N9343), .B(N8965));
NOR3BX1 inst_cellmath__203_0_I8501 (.Y(N9736), .AN(N6479), .B(N6585), .C(N6119));
NAND2XL hyperpropagate_3_1_A_I8519 (.Y(N19032), .A(N6053), .B(N5952));
NOR2XL hyperpropagate_3_1_A_I8520 (.Y(N10101), .A(N6167), .B(N19032));
NOR3BX1 inst_cellmath__203_0_I8502 (.Y(N8766), .AN(N6178), .B(N6289), .C(N6640));
NOR3BX1 inst_cellmath__203_0_I8503 (.Y(N9115), .AN(N6222), .B(N6146), .C(N6038));
NOR4X1 inst_cellmath__203_0_I8455 (.Y(N9507), .A(N6544), .B(N5893), .C(N6606), .D(N6272));
AND2XL inst_cellmath__203_0_I8456 (.Y(N9888), .A(N6672), .B(N6486));
NOR4X1 inst_cellmath__203_0_I8457 (.Y(N10248), .A(N6175), .B(N6359), .C(N6527), .D(N6254));
NOR3BX1 inst_cellmath__203_0_I8504 (.Y(N8907), .AN(N6298), .B(N6392), .C(N6573));
AND2XL inst_cellmath__203_0_I8459 (.Y(N8716), .A(N6536), .B(N5887));
NOR3BX1 inst_cellmath__203_0_I8505 (.Y(N9055), .AN(N6587), .B(N6043), .C(N6232));
NOR4X1 inst_cellmath__203_0_I8461 (.Y(N9437), .A(N6247), .B(N5990), .C(N6353), .D(N6418));
NOR3X1 inst_cellmath__203_0_I8462 (.Y(N9825), .A(N6566), .B(N6102), .C(N6000));
NOR2BX1 inst_cellmath__203_0_I8463 (.Y(N10183), .AN(N6227), .B(N5851));
NOR3BX1 inst_cellmath__203_0_I8506 (.Y(N9208), .AN(N6678), .B(N5951), .C(N6135));
NOR2BX1 inst_cellmath__203_0_I8465 (.Y(N9599), .AN(N5964), .B(N6257));
NOR4X1 inst_cellmath__203_0_I8466 (.Y(N9978), .A(N6396), .B(N5931), .C(N6640), .D(N6576));
NOR4X1 inst_cellmath__203_0_I8467 (.Y(N8664), .A(N6542), .B(N6443), .C(N6078), .D(N6270));
NOR2BX1 inst_cellmath__203_0_I8468 (.Y(N8993), .AN(N6131), .B(N6591));
NOR2XL inst_cellmath__203_0_I2626 (.Y(N9564), .A(N7975), .B(N9736));
NOR2XL inst_cellmath__203_0_I2627 (.Y(N10296), .A(N7975), .B(N10101));
NOR2XL inst_cellmath__203_0_I2628 (.Y(N9336), .A(N7975), .B(N8766));
NOR2XL inst_cellmath__203_0_I2629 (.Y(N10091), .A(N7975), .B(N9115));
NOR2XL inst_cellmath__203_0_I2630 (.Y(N9106), .A(N7975), .B(N9507));
NOR2XL inst_cellmath__203_0_I2631 (.Y(N9882), .A(N7975), .B(N9888));
NOR2XL inst_cellmath__203_0_I2632 (.Y(N8897), .A(N7975), .B(N10248));
NOR2XL inst_cellmath__203_0_I2633 (.Y(N9664), .A(N7975), .B(N8907));
NOR2XL inst_cellmath__203_0_I2634 (.Y(N8712), .A(N7975), .B(N9277));
NOR2XL inst_cellmath__203_0_I2635 (.Y(N9430), .A(N7975), .B(N9670));
NOR2XL inst_cellmath__203_0_I2636 (.Y(N10175), .A(N7975), .B(N10038));
NOR2XL inst_cellmath__203_0_I2637 (.Y(N9203), .A(N7975), .B(N8716));
NOR2XL inst_cellmath__203_0_I2638 (.Y(N9969), .A(N7975), .B(N9055));
NOR2XL inst_cellmath__203_0_I2639 (.Y(N8985), .A(N7975), .B(N9437));
NOR2XL inst_cellmath__203_0_I2640 (.Y(N9755), .A(N7975), .B(N9825));
NOR2XL inst_cellmath__203_0_I2641 (.Y(N8784), .A(N7975), .B(N10183));
NOR2XL inst_cellmath__203_0_I2642 (.Y(N9171), .A(N7975), .B(N8842));
NOR2XL inst_cellmath__203_0_I2643 (.Y(N9907), .A(N7975), .B(N9208));
NOR2XL inst_cellmath__203_0_I2644 (.Y(N9297), .A(N7975), .B(N9599));
NOR2XL inst_cellmath__203_0_I2645 (.Y(N8854), .A(N7975), .B(N9978));
NOR2XL inst_cellmath__203_0_I2646 (.Y(N8824), .A(N7975), .B(N8664));
NOR2XL inst_cellmath__203_0_I2647 (.Y(N9847), .A(N7975), .B(N8993));
NAND2BX1 inst_cellmath__203_0_I2649 (.Y(N9144), .AN(inst_cellmath__61[2]), .B(inst_cellmath__61[1]));
NOR2XL inst_cellmath__203_0_I2651 (.Y(N8686), .A(N9736), .B(N7958));
MXI2XL inst_cellmath__203_0_I2652 (.Y(N10138), .A(N7696), .B(N9144), .S0(N8686));
MXI2XL inst_cellmath__203_0_I2653 (.Y(N10297), .A(N10101), .B(N9736), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2654 (.Y(N8804), .A(N7696), .B(N9144), .S0(N10297));
MXI2XL inst_cellmath__203_0_I2655 (.Y(N10238), .A(N8766), .B(N10101), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2656 (.Y(N9165), .A(N7696), .B(N9144), .S0(N10238));
MXI2XL inst_cellmath__203_0_I2657 (.Y(N10176), .A(N9115), .B(N8766), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2658 (.Y(N9557), .A(N7696), .B(N9144), .S0(N10176));
MXI2XL inst_cellmath__203_0_I2659 (.Y(N10116), .A(N9507), .B(N9115), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2660 (.Y(N9934), .A(N7696), .B(N9144), .S0(N10116));
MXI2XL inst_cellmath__203_0_I2661 (.Y(N10055), .A(N9888), .B(N9507), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2662 (.Y(N10288), .A(N7696), .B(N9144), .S0(N10055));
MXI2XL inst_cellmath__203_0_I2663 (.Y(N9995), .A(N10248), .B(N9888), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2664 (.Y(N8946), .A(N7696), .B(N9144), .S0(N9995));
MXI2XL inst_cellmath__203_0_I2665 (.Y(N9935), .A(N8907), .B(N10248), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2666 (.Y(N9329), .A(N7696), .B(N9144), .S0(N9935));
MXI2XL inst_cellmath__203_0_I2667 (.Y(N9874), .A(N9277), .B(N8907), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2668 (.Y(N9719), .A(N7696), .B(N9144), .S0(N9874));
MXI2XL inst_cellmath__203_0_I2669 (.Y(N9810), .A(N9670), .B(N9277), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2670 (.Y(N10080), .A(N7696), .B(N9144), .S0(N9810));
MXI2XL inst_cellmath__203_0_I2671 (.Y(N9749), .A(N10038), .B(N9670), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2672 (.Y(N8750), .A(N7696), .B(N9144), .S0(N9749));
MXI2XL inst_cellmath__203_0_I2673 (.Y(N9682), .A(N8716), .B(N10038), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2674 (.Y(N9099), .A(N7696), .B(N9144), .S0(N9682));
MXI2XL inst_cellmath__203_0_I2675 (.Y(N9614), .A(N9055), .B(N8716), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2676 (.Y(N9488), .A(N7696), .B(N9144), .S0(N9614));
MXI2XL inst_cellmath__203_0_I2677 (.Y(N9550), .A(N9437), .B(N9055), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2678 (.Y(N9873), .A(N7696), .B(N9144), .S0(N9550));
MXI2XL inst_cellmath__203_0_I2679 (.Y(N9481), .A(N9825), .B(N9437), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2680 (.Y(N10232), .A(N7696), .B(N9144), .S0(N9481));
MXI2XL inst_cellmath__203_0_I2681 (.Y(N9415), .A(N10183), .B(N9825), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2682 (.Y(N8888), .A(N7696), .B(N9144), .S0(N9415));
MXI2XL inst_cellmath__203_0_I2683 (.Y(N9349), .A(N8842), .B(N10183), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2684 (.Y(N9261), .A(N7696), .B(N9144), .S0(N9349));
MXI2XL inst_cellmath__203_0_I2685 (.Y(N9281), .A(N9208), .B(N8842), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2686 (.Y(N9654), .A(N7696), .B(N9144), .S0(N9281));
MXI2XL inst_cellmath__203_0_I2687 (.Y(N9216), .A(N9599), .B(N9208), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2688 (.Y(N10018), .A(N7696), .B(N9144), .S0(N9216));
MXI2XL inst_cellmath__203_0_I2689 (.Y(N9150), .A(N9978), .B(N9599), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2690 (.Y(N8702), .A(N7696), .B(N9144), .S0(N9150));
MXI2XL inst_cellmath__203_0_I2691 (.Y(N9086), .A(N8664), .B(N9978), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2692 (.Y(N9040), .A(N7696), .B(N9144), .S0(N9086));
MXI2XL inst_cellmath__203_0_I2693 (.Y(N9026), .A(N8993), .B(N8664), .S0(N7958));
MXI2XL inst_cellmath__203_0_I2694 (.Y(N9421), .A(N7696), .B(N9144), .S0(N9026));
NOR2BX1 inst_cellmath__203_0_I2695 (.Y(N8962), .AN(N7958), .B(N8993));
MXI2XL inst_cellmath__203_0_I2696 (.Y(N9808), .A(N7696), .B(N9144), .S0(N8962));
XNOR2X1 inst_cellmath__203_0_I2697 (.Y(N9586), .A(inst_cellmath__61[3]), .B(inst_cellmath__61[2]));
NOR2XL inst_cellmath__203_0_I2698 (.Y(N9668), .A(inst_cellmath__61[3]), .B(inst_cellmath__61[2]));
OAI2BB1X1 inst_cellmath__203_0_I2699 (.Y(N9196), .A0N(inst_cellmath__61[3]), .A1N(inst_cellmath__61[2]), .B0(inst_cellmath__61[4]));
INVXL inst_cellmath__203_0_I2700 (.Y(N9918), .A(N9196));
OR2XL inst_cellmath__203_0_I2701 (.Y(N9306), .A(N9668), .B(inst_cellmath__61[4]));
INVXL inst_cellmath__203_0_I2702 (.Y(N9698), .A(N9918));
NOR2XL inst_cellmath__203_0_I2703 (.Y(N8662), .A(N9736), .B(N9586));
MXI2XL inst_cellmath__203_0_I2704 (.Y(N10112), .A(N9698), .B(N9306), .S0(N8662));
MXI2XL inst_cellmath__203_0_I2705 (.Y(N10269), .A(N10101), .B(N9736), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2706 (.Y(N8777), .A(N9698), .B(N9306), .S0(N10269));
MXI2XL inst_cellmath__203_0_I2707 (.Y(N10209), .A(N8766), .B(N10101), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2708 (.Y(N9130), .A(N9698), .B(N9306), .S0(N10209));
MXI2XL inst_cellmath__203_0_I2709 (.Y(N10145), .A(N9115), .B(N8766), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2710 (.Y(N9521), .A(N9698), .B(N9306), .S0(N10145));
MXI2XL inst_cellmath__203_0_I2711 (.Y(N10090), .A(N9507), .B(N9115), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2712 (.Y(N9897), .A(N9698), .B(N9306), .S0(N10090));
MXI2XL inst_cellmath__203_0_I2713 (.Y(N10028), .A(N9888), .B(N9507), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2714 (.Y(N10258), .A(N9698), .B(N9306), .S0(N10028));
MXI2XL inst_cellmath__203_0_I2715 (.Y(N9968), .A(N10248), .B(N9888), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2716 (.Y(N8917), .A(N9698), .B(N9306), .S0(N9968));
MXI2XL inst_cellmath__203_0_I2717 (.Y(N9906), .A(N8907), .B(N10248), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2718 (.Y(N9287), .A(N9698), .B(N9306), .S0(N9906));
MXI2XL inst_cellmath__203_0_I2719 (.Y(N9845), .A(N9277), .B(N8907), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2720 (.Y(N9681), .A(N9698), .B(N9306), .S0(N9845));
MXI2XL inst_cellmath__203_0_I2721 (.Y(N9780), .A(N9670), .B(N9277), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2722 (.Y(N10048), .A(N9698), .B(N9306), .S0(N9780));
MXI2XL inst_cellmath__203_0_I2723 (.Y(N9717), .A(N10038), .B(N9670), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2724 (.Y(N8727), .A(N9698), .B(N9306), .S0(N9717));
MXI2XL inst_cellmath__203_0_I2725 (.Y(N9651), .A(N8716), .B(N10038), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2726 (.Y(N9068), .A(N9698), .B(N9306), .S0(N9651));
MXI2XL inst_cellmath__203_0_I2727 (.Y(N9583), .A(N9055), .B(N8716), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2728 (.Y(N9451), .A(N9698), .B(N9306), .S0(N9583));
MXI2XL inst_cellmath__203_0_I2729 (.Y(N9519), .A(N9437), .B(N9055), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2730 (.Y(N9836), .A(N9698), .B(N9306), .S0(N9519));
MXI2XL inst_cellmath__203_0_I2731 (.Y(N9449), .A(N9825), .B(N9437), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2732 (.Y(N10195), .A(N9698), .B(N9306), .S0(N9449));
MXI2XL inst_cellmath__203_0_I2733 (.Y(N9384), .A(N10183), .B(N9825), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2734 (.Y(N8855), .A(N9698), .B(N9306), .S0(N9384));
MXI2XL inst_cellmath__203_0_I2735 (.Y(N9320), .A(N8842), .B(N10183), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2736 (.Y(N9223), .A(N9698), .B(N9306), .S0(N9320));
MXI2XL inst_cellmath__203_0_I2737 (.Y(N9250), .A(N9208), .B(N8842), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2738 (.Y(N9613), .A(N9698), .B(N9306), .S0(N9250));
MXI2XL inst_cellmath__203_0_I2739 (.Y(N9184), .A(N9599), .B(N9208), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2740 (.Y(N9986), .A(N9698), .B(N9306), .S0(N9184));
MXI2XL inst_cellmath__203_0_I2741 (.Y(N9119), .A(N9978), .B(N9599), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2742 (.Y(N8673), .A(N9698), .B(N9306), .S0(N9119));
MXI2XL inst_cellmath__203_0_I2743 (.Y(N9058), .A(N8664), .B(N9978), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2744 (.Y(N9007), .A(N9698), .B(N9306), .S0(N9058));
MXI2XL inst_cellmath__203_0_I2745 (.Y(N8997), .A(N8993), .B(N8664), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2746 (.Y(N9386), .A(N9698), .B(N9306), .S0(N8997));
NOR2BX1 inst_cellmath__203_0_I2747 (.Y(N8934), .AN(N9586), .B(N8993));
MXI2XL inst_cellmath__203_0_I2748 (.Y(N9774), .A(N9698), .B(N9306), .S0(N8934));
XNOR2X1 inst_cellmath__203_0_I2749 (.Y(N9549), .A(inst_cellmath__61[5]), .B(inst_cellmath__61[4]));
NOR2XL inst_cellmath__203_0_I2750 (.Y(N9634), .A(inst_cellmath__61[5]), .B(inst_cellmath__61[4]));
OAI2BB1X1 inst_cellmath__203_0_I2751 (.Y(N9157), .A0N(inst_cellmath__61[5]), .A1N(inst_cellmath__61[4]), .B0(inst_cellmath__61[6]));
INVXL inst_cellmath__203_0_I2752 (.Y(N10064), .A(N9157));
OR2XL inst_cellmath__203_0_I2753 (.Y(N9467), .A(N9634), .B(inst_cellmath__61[6]));
INVXL inst_cellmath__203_0_I2754 (.Y(N9857), .A(N10064));
NOR2XL inst_cellmath__203_0_I2755 (.Y(N10299), .A(N9736), .B(N9549));
MXI2XL inst_cellmath__203_0_I2756 (.Y(N10074), .A(N9857), .B(N9467), .S0(N10299));
MXI2XL inst_cellmath__203_0_I2757 (.Y(N10242), .A(N10101), .B(N9736), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2758 (.Y(N8746), .A(N9857), .B(N9467), .S0(N10242));
MXI2XL inst_cellmath__203_0_I2759 (.Y(N10178), .A(N8766), .B(N10101), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2760 (.Y(N9094), .A(N9857), .B(N9467), .S0(N10178));
MXI2XL inst_cellmath__203_0_I2761 (.Y(N10119), .A(N9115), .B(N8766), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2762 (.Y(N9479), .A(N9857), .B(N9467), .S0(N10119));
MXI2XL inst_cellmath__203_0_I2763 (.Y(N10057), .A(N9507), .B(N9115), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2764 (.Y(N9865), .A(N9857), .B(N9467), .S0(N10057));
MXI2XL inst_cellmath__203_0_I2765 (.Y(N9998), .A(N9888), .B(N9507), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2766 (.Y(N10224), .A(N9857), .B(N9467), .S0(N9998));
MXI2XL inst_cellmath__203_0_I2767 (.Y(N9939), .A(N10248), .B(N9888), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2768 (.Y(N8882), .A(N9857), .B(N9467), .S0(N9939));
MXI2XL inst_cellmath__203_0_I2769 (.Y(N9876), .A(N8907), .B(N10248), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2770 (.Y(N9252), .A(N9857), .B(N9467), .S0(N9876));
MXI2XL inst_cellmath__203_0_I2771 (.Y(N9813), .A(N9277), .B(N8907), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2772 (.Y(N9644), .A(N9857), .B(N9467), .S0(N9813));
MXI2XL inst_cellmath__203_0_I2773 (.Y(N9752), .A(N9670), .B(N9277), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2774 (.Y(N10012), .A(N9857), .B(N9467), .S0(N9752));
MXI2XL inst_cellmath__203_0_I2775 (.Y(N9684), .A(N10038), .B(N9670), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2776 (.Y(N8696), .A(N9857), .B(N9467), .S0(N9684));
MXI2XL inst_cellmath__203_0_I2777 (.Y(N9617), .A(N8716), .B(N10038), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2778 (.Y(N9032), .A(N9857), .B(N9467), .S0(N9617));
MXI2XL inst_cellmath__203_0_I2779 (.Y(N9554), .A(N9055), .B(N8716), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2780 (.Y(N9413), .A(N9857), .B(N9467), .S0(N9554));
MXI2XL inst_cellmath__203_0_I2781 (.Y(N9484), .A(N9437), .B(N9055), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2782 (.Y(N9800), .A(N9857), .B(N9467), .S0(N9484));
MXI2XL inst_cellmath__203_0_I2783 (.Y(N9418), .A(N9825), .B(N9437), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2784 (.Y(N10161), .A(N9857), .B(N9467), .S0(N9418));
MXI2XL inst_cellmath__203_0_I2785 (.Y(N9353), .A(N10183), .B(N9825), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2786 (.Y(N8823), .A(N9857), .B(N9467), .S0(N9353));
MXI2XL inst_cellmath__203_0_I2787 (.Y(N9283), .A(N8842), .B(N10183), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2788 (.Y(N9186), .A(N9857), .B(N9467), .S0(N9283));
MXI2XL inst_cellmath__203_0_I2789 (.Y(N9218), .A(N9208), .B(N8842), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2790 (.Y(N9576), .A(N9857), .B(N9467), .S0(N9218));
MXI2XL inst_cellmath__203_0_I2791 (.Y(N9152), .A(N9599), .B(N9208), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2792 (.Y(N9955), .A(N9857), .B(N9467), .S0(N9152));
MXI2XL inst_cellmath__203_0_I2793 (.Y(N9088), .A(N9978), .B(N9599), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2794 (.Y(N10307), .A(N9857), .B(N9467), .S0(N9088));
MXI2XL inst_cellmath__203_0_I2795 (.Y(N9028), .A(N8664), .B(N9978), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2796 (.Y(N8971), .A(N9857), .B(N9467), .S0(N9028));
MXI2XL inst_cellmath__203_0_I2797 (.Y(N8964), .A(N8993), .B(N8664), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2798 (.Y(N9347), .A(N9857), .B(N9467), .S0(N8964));
NOR2BX1 inst_cellmath__203_0_I2799 (.Y(N8906), .AN(N9549), .B(N8993));
MXI2XL inst_cellmath__203_0_I2800 (.Y(N9740), .A(N9857), .B(N9467), .S0(N8906));
XNOR2X1 inst_cellmath__203_0_I2801 (.Y(N9512), .A(inst_cellmath__61[7]), .B(inst_cellmath__61[6]));
NOR2XL inst_cellmath__203_0_I2802 (.Y(N9600), .A(inst_cellmath__61[7]), .B(inst_cellmath__61[6]));
OAI2BB1X1 inst_cellmath__203_0_I2803 (.Y(N9121), .A0N(inst_cellmath__61[7]), .A1N(inst_cellmath__61[6]), .B0(inst_cellmath__61[8]));
INVXL inst_cellmath__203_0_I2804 (.Y(N10213), .A(N9121));
OR2XL inst_cellmath__203_0_I2805 (.Y(N9632), .A(N9600), .B(inst_cellmath__61[8]));
INVXL inst_cellmath__203_0_I2806 (.Y(N10003), .A(N10213));
NOR2XL inst_cellmath__203_0_I2807 (.Y(N10272), .A(N9736), .B(N9512));
MXI2XL inst_cellmath__203_0_I2808 (.Y(N10041), .A(N10003), .B(N9632), .S0(N10272));
MXI2XL inst_cellmath__203_0_I2809 (.Y(N10212), .A(N10101), .B(N9736), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2810 (.Y(N8720), .A(N10003), .B(N9632), .S0(N10212));
MXI2XL inst_cellmath__203_0_I2811 (.Y(N10147), .A(N8766), .B(N10101), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2812 (.Y(N9060), .A(N10003), .B(N9632), .S0(N10147));
MXI2XL inst_cellmath__203_0_I2813 (.Y(N10093), .A(N9115), .B(N8766), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2814 (.Y(N9442), .A(N10003), .B(N9632), .S0(N10093));
MXI2XL inst_cellmath__203_0_I2815 (.Y(N10030), .A(N9507), .B(N9115), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2816 (.Y(N9828), .A(N10003), .B(N9632), .S0(N10030));
MXI2XL inst_cellmath__203_0_I2817 (.Y(N9971), .A(N9888), .B(N9507), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2818 (.Y(N10189), .A(N10003), .B(N9632), .S0(N9971));
MXI2XL inst_cellmath__203_0_I2819 (.Y(N9908), .A(N10248), .B(N9888), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2820 (.Y(N8848), .A(N10003), .B(N9632), .S0(N9908));
MXI2XL inst_cellmath__203_0_I2821 (.Y(N9848), .A(N8907), .B(N10248), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2822 (.Y(N9213), .A(N10003), .B(N9632), .S0(N9848));
MXI2XL inst_cellmath__203_0_I2823 (.Y(N9782), .A(N9277), .B(N8907), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2824 (.Y(N9605), .A(N10003), .B(N9632), .S0(N9782));
MXI2XL inst_cellmath__203_0_I2825 (.Y(N9720), .A(N9670), .B(N9277), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2826 (.Y(N9981), .A(N10003), .B(N9632), .S0(N9720));
MXI2XL inst_cellmath__203_0_I2827 (.Y(N9655), .A(N10038), .B(N9670), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2828 (.Y(N8667), .A(N10003), .B(N9632), .S0(N9655));
MXI2XL inst_cellmath__203_0_I2829 (.Y(N9587), .A(N8716), .B(N10038), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2830 (.Y(N8998), .A(N10003), .B(N9632), .S0(N9587));
MXI2XL inst_cellmath__203_0_I2831 (.Y(N9522), .A(N9055), .B(N8716), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2832 (.Y(N9377), .A(N10003), .B(N9632), .S0(N9522));
MXI2XL inst_cellmath__203_0_I2833 (.Y(N9452), .A(N9437), .B(N9055), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2834 (.Y(N9765), .A(N10003), .B(N9632), .S0(N9452));
MXI2XL inst_cellmath__203_0_I2835 (.Y(N9387), .A(N9825), .B(N9437), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2836 (.Y(N10129), .A(N10003), .B(N9632), .S0(N9387));
MXI2XL inst_cellmath__203_0_I2837 (.Y(N9322), .A(N10183), .B(N9825), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2838 (.Y(N8793), .A(N10003), .B(N9632), .S0(N9322));
MXI2XL inst_cellmath__203_0_I2839 (.Y(N9253), .A(N8842), .B(N10183), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2840 (.Y(N9148), .A(N10003), .B(N9632), .S0(N9253));
MXI2XL inst_cellmath__203_0_I2841 (.Y(N9187), .A(N9208), .B(N8842), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2842 (.Y(N9541), .A(N10003), .B(N9632), .S0(N9187));
MXI2XL inst_cellmath__203_0_I2843 (.Y(N9122), .A(N9599), .B(N9208), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2844 (.Y(N9923), .A(N10003), .B(N9632), .S0(N9122));
MXI2XL inst_cellmath__203_0_I2845 (.Y(N9061), .A(N9978), .B(N9599), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2846 (.Y(N10276), .A(N10003), .B(N9632), .S0(N9061));
MXI2XL inst_cellmath__203_0_I2847 (.Y(N8999), .A(N8664), .B(N9978), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2848 (.Y(N8936), .A(N10003), .B(N9632), .S0(N8999));
MXI2XL inst_cellmath__203_0_I2849 (.Y(N8937), .A(N8993), .B(N8664), .S0(N9512));
MXI2XL inst_cellmath__203_0_I2850 (.Y(N9313), .A(N10003), .B(N9632), .S0(N8937));
NOR2BX1 inst_cellmath__203_0_I2851 (.Y(N8875), .AN(N9512), .B(N8993));
MXI2XL inst_cellmath__203_0_I2852 (.Y(N9702), .A(N10003), .B(N9632), .S0(N8875));
XNOR2X1 inst_cellmath__203_0_I2853 (.Y(N9470), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
NOR2XL inst_cellmath__203_0_I2854 (.Y(N9569), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
OAI2BB1X1 inst_cellmath__203_0_I2855 (.Y(N9083), .A0N(inst_cellmath__61[9]), .A1N(inst_cellmath__61[8]), .B0(inst_cellmath__61[10]));
INVXL inst_cellmath__203_0_I2856 (.Y(N8687), .A(N9083));
OR2XL inst_cellmath__203_0_I2857 (.Y(N9790), .A(N9569), .B(inst_cellmath__61[10]));
INVXL inst_cellmath__203_0_I2858 (.Y(N10148), .A(N8687));
NOR2XL inst_cellmath__203_0_I2859 (.Y(N10246), .A(N9736), .B(N9470));
MXI2XL inst_cellmath__203_0_I2860 (.Y(N10007), .A(N10148), .B(N9790), .S0(N10246));
MXI2XL inst_cellmath__203_0_I2861 (.Y(N10181), .A(N10101), .B(N9736), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2862 (.Y(N8690), .A(N10148), .B(N9790), .S0(N10181));
MXI2XL inst_cellmath__203_0_I2863 (.Y(N10123), .A(N8766), .B(N10101), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2864 (.Y(N9025), .A(N10148), .B(N9790), .S0(N10123));
MXI2XL inst_cellmath__203_0_I2865 (.Y(N10061), .A(N9115), .B(N8766), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2866 (.Y(N9404), .A(N10148), .B(N9790), .S0(N10061));
MXI2XL inst_cellmath__203_0_I2867 (.Y(N10000), .A(N9507), .B(N9115), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2868 (.Y(N9793), .A(N10148), .B(N9790), .S0(N10000));
MXI2XL inst_cellmath__203_0_I2869 (.Y(N9943), .A(N9888), .B(N9507), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2870 (.Y(N10154), .A(N10148), .B(N9790), .S0(N9943));
MXI2XL inst_cellmath__203_0_I2871 (.Y(N9880), .A(N10248), .B(N9888), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2872 (.Y(N8814), .A(N10148), .B(N9790), .S0(N9880));
MXI2XL inst_cellmath__203_0_I2873 (.Y(N9817), .A(N8907), .B(N10248), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2874 (.Y(N9176), .A(N10148), .B(N9790), .S0(N9817));
MXI2XL inst_cellmath__203_0_I2875 (.Y(N9754), .A(N9277), .B(N8907), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2876 (.Y(N9568), .A(N10148), .B(N9790), .S0(N9754));
MXI2XL inst_cellmath__203_0_I2877 (.Y(N9688), .A(N9670), .B(N9277), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2878 (.Y(N9948), .A(N10148), .B(N9790), .S0(N9688));
MXI2XL inst_cellmath__203_0_I2879 (.Y(N9621), .A(N10038), .B(N9670), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2880 (.Y(N10300), .A(N10148), .B(N9790), .S0(N9621));
MXI2XL inst_cellmath__203_0_I2881 (.Y(N9556), .A(N8716), .B(N10038), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2882 (.Y(N8961), .A(N10148), .B(N9790), .S0(N9556));
MXI2XL inst_cellmath__203_0_I2883 (.Y(N9487), .A(N9055), .B(N8716), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2884 (.Y(N9338), .A(N10148), .B(N9790), .S0(N9487));
MXI2XL inst_cellmath__203_0_I2885 (.Y(N9420), .A(N9437), .B(N9055), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2886 (.Y(N9733), .A(N10148), .B(N9790), .S0(N9420));
MXI2XL inst_cellmath__203_0_I2887 (.Y(N9355), .A(N9825), .B(N9437), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2888 (.Y(N10098), .A(N10148), .B(N9790), .S0(N9355));
MXI2XL inst_cellmath__203_0_I2889 (.Y(N9286), .A(N10183), .B(N9825), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2890 (.Y(N8762), .A(N10148), .B(N9790), .S0(N9286));
MXI2XL inst_cellmath__203_0_I2891 (.Y(N9222), .A(N8842), .B(N10183), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2892 (.Y(N9111), .A(N10148), .B(N9790), .S0(N9222));
MXI2XL inst_cellmath__203_0_I2893 (.Y(N9155), .A(N9208), .B(N8842), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2894 (.Y(N9503), .A(N10148), .B(N9790), .S0(N9155));
MXI2XL inst_cellmath__203_0_I2895 (.Y(N9091), .A(N9599), .B(N9208), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2896 (.Y(N9885), .A(N10148), .B(N9790), .S0(N9091));
MXI2XL inst_cellmath__203_0_I2897 (.Y(N9031), .A(N9978), .B(N9599), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2898 (.Y(N10244), .A(N10148), .B(N9790), .S0(N9031));
MXI2XL inst_cellmath__203_0_I2899 (.Y(N8969), .A(N8664), .B(N9978), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2900 (.Y(N8904), .A(N10148), .B(N9790), .S0(N8969));
MXI2XL inst_cellmath__203_0_I2901 (.Y(N8910), .A(N8993), .B(N8664), .S0(N9470));
MXI2XL inst_cellmath__203_0_I2902 (.Y(N9271), .A(N10148), .B(N9790), .S0(N8910));
NOR2BX1 inst_cellmath__203_0_I2903 (.Y(N8846), .AN(N9470), .B(N8993));
MXI2XL inst_cellmath__203_0_I2904 (.Y(N9667), .A(N10148), .B(N9790), .S0(N8846));
XNOR2X1 inst_cellmath__203_0_I2905 (.Y(N9435), .A(inst_cellmath__61[11]), .B(inst_cellmath__61[10]));
NOR2XL inst_cellmath__203_0_I2906 (.Y(N9539), .A(inst_cellmath__61[11]), .B(inst_cellmath__61[10]));
OAI2BB1X1 inst_cellmath__203_0_I2907 (.Y(N9052), .A0N(inst_cellmath__61[11]), .A1N(inst_cellmath__61[10]), .B0(inst_cellmath__61[12]));
INVXL inst_cellmath__203_0_I2908 (.Y(N8812), .A(N9052));
OR2XL inst_cellmath__203_0_I2909 (.Y(N9945), .A(N9539), .B(inst_cellmath__61[12]));
INVXL inst_cellmath__203_0_I2910 (.Y(N10298), .A(N8812));
NOR2XL inst_cellmath__203_0_I2911 (.Y(N10217), .A(N9736), .B(N9435));
MXI2XL inst_cellmath__203_0_I2912 (.Y(N9975), .A(N10298), .B(N9945), .S0(N10217));
MXI2XL inst_cellmath__203_0_I2913 (.Y(N10151), .A(N10101), .B(N9736), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2914 (.Y(N8660), .A(N10298), .B(N9945), .S0(N10151));
MXI2XL inst_cellmath__203_0_I2915 (.Y(N10096), .A(N8766), .B(N10101), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2916 (.Y(N8989), .A(N10298), .B(N9945), .S0(N10096));
MXI2XL inst_cellmath__203_0_I2917 (.Y(N10033), .A(N9115), .B(N8766), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2918 (.Y(N9368), .A(N10298), .B(N9945), .S0(N10033));
MXI2XL inst_cellmath__203_0_I2919 (.Y(N9973), .A(N9507), .B(N9115), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2920 (.Y(N9758), .A(N10298), .B(N9945), .S0(N9973));
MXI2XL inst_cellmath__203_0_I2921 (.Y(N9911), .A(N9888), .B(N9507), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2922 (.Y(N10121), .A(N10298), .B(N9945), .S0(N9911));
MXI2XL inst_cellmath__203_0_I2923 (.Y(N9850), .A(N10248), .B(N9888), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2924 (.Y(N8787), .A(N10298), .B(N9945), .S0(N9850));
MXI2XL inst_cellmath__203_0_I2925 (.Y(N9786), .A(N8907), .B(N10248), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2926 (.Y(N9138), .A(N10298), .B(N9945), .S0(N9786));
MXI2XL inst_cellmath__203_0_I2927 (.Y(N9724), .A(N9277), .B(N8907), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2928 (.Y(N9531), .A(N10298), .B(N9945), .S0(N9724));
MXI2XL inst_cellmath__203_0_I2929 (.Y(N9658), .A(N9670), .B(N9277), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2930 (.Y(N9914), .A(N10298), .B(N9945), .S0(N9658));
MXI2XL inst_cellmath__203_0_I2931 (.Y(N9590), .A(N10038), .B(N9670), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2932 (.Y(N10267), .A(N10298), .B(N9945), .S0(N9590));
MXI2XL inst_cellmath__203_0_I2933 (.Y(N9525), .A(N8716), .B(N10038), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2934 (.Y(N8927), .A(N10298), .B(N9945), .S0(N9525));
MXI2XL inst_cellmath__203_0_I2935 (.Y(N9455), .A(N9055), .B(N8716), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2936 (.Y(N9302), .A(N10298), .B(N9945), .S0(N9455));
MXI2XL inst_cellmath__203_0_I2937 (.Y(N9390), .A(N9437), .B(N9055), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2938 (.Y(N9693), .A(N10298), .B(N9945), .S0(N9390));
MXI2XL inst_cellmath__203_0_I2939 (.Y(N9325), .A(N9825), .B(N9437), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2940 (.Y(N10059), .A(N10298), .B(N9945), .S0(N9325));
MXI2XL inst_cellmath__203_0_I2941 (.Y(N9256), .A(N10183), .B(N9825), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2942 (.Y(N8738), .A(N10298), .B(N9945), .S0(N9256));
MXI2XL inst_cellmath__203_0_I2943 (.Y(N9190), .A(N8842), .B(N10183), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2944 (.Y(N9075), .A(N10298), .B(N9945), .S0(N9190));
MXI2XL inst_cellmath__203_0_I2945 (.Y(N9126), .A(N9208), .B(N8842), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2946 (.Y(N9463), .A(N10298), .B(N9945), .S0(N9126));
MXI2XL inst_cellmath__203_0_I2947 (.Y(N9065), .A(N9599), .B(N9208), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2948 (.Y(N9853), .A(N10298), .B(N9945), .S0(N9065));
MXI2XL inst_cellmath__203_0_I2949 (.Y(N9002), .A(N9978), .B(N9599), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2950 (.Y(N10206), .A(N10298), .B(N9945), .S0(N9002));
MXI2XL inst_cellmath__203_0_I2951 (.Y(N8939), .A(N8664), .B(N9978), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2952 (.Y(N8867), .A(N10298), .B(N9945), .S0(N8939));
MXI2XL inst_cellmath__203_0_I2953 (.Y(N8877), .A(N8993), .B(N8664), .S0(N9435));
MXI2XL inst_cellmath__203_0_I2954 (.Y(N9238), .A(N10298), .B(N9945), .S0(N8877));
NOR2BX1 inst_cellmath__203_0_I2955 (.Y(N8818), .AN(N9435), .B(N8993));
MXI2XL inst_cellmath__203_0_I2956 (.Y(N9627), .A(N10298), .B(N9945), .S0(N8818));
XNOR2X1 inst_cellmath__203_0_I2957 (.Y(N9401), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
NOR2XL inst_cellmath__203_0_I2958 (.Y(N9506), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
OAI2BB1X1 inst_cellmath__203_0_I2959 (.Y(N9016), .A0N(inst_cellmath__61[13]), .A1N(inst_cellmath__61[12]), .B0(inst_cellmath__61[14]));
INVXL inst_cellmath__203_0_I2960 (.Y(N8956), .A(N9016));
OR2XL inst_cellmath__203_0_I2961 (.Y(N10094), .A(N9506), .B(inst_cellmath__61[14]));
INVXL inst_cellmath__203_0_I2962 (.Y(N8759), .A(N8956));
NOR2XL inst_cellmath__203_0_I2963 (.Y(N10184), .A(N9736), .B(N9401));
MXI2XL inst_cellmath__203_0_I2964 (.Y(N9941), .A(N8759), .B(N10094), .S0(N10184));
MXI2XL inst_cellmath__203_0_I2965 (.Y(N10125), .A(N10101), .B(N9736), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2966 (.Y(N10294), .A(N8759), .B(N10094), .S0(N10125));
MXI2XL inst_cellmath__203_0_I2967 (.Y(N10065), .A(N8766), .B(N10101), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2968 (.Y(N8951), .A(N8759), .B(N10094), .S0(N10065));
MXI2XL inst_cellmath__203_0_I2969 (.Y(N10004), .A(N9115), .B(N8766), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2970 (.Y(N9333), .A(N8759), .B(N10094), .S0(N10004));
MXI2XL inst_cellmath__203_0_I2971 (.Y(N9946), .A(N9507), .B(N9115), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2972 (.Y(N9727), .A(N8759), .B(N10094), .S0(N9946));
MXI2XL inst_cellmath__203_0_I2973 (.Y(N9883), .A(N9888), .B(N9507), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2974 (.Y(N10087), .A(N8759), .B(N10094), .S0(N9883));
MXI2XL inst_cellmath__203_0_I2975 (.Y(N9819), .A(N10248), .B(N9888), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2976 (.Y(N8756), .A(N8759), .B(N10094), .S0(N9819));
MXI2XL inst_cellmath__203_0_I2977 (.Y(N9756), .A(N8907), .B(N10248), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2978 (.Y(N9102), .A(N8759), .B(N10094), .S0(N9756));
MXI2XL inst_cellmath__203_0_I2979 (.Y(N9690), .A(N9277), .B(N8907), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2980 (.Y(N9493), .A(N8759), .B(N10094), .S0(N9690));
MXI2XL inst_cellmath__203_0_I2981 (.Y(N9624), .A(N9670), .B(N9277), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2982 (.Y(N9878), .A(N8759), .B(N10094), .S0(N9624));
MXI2XL inst_cellmath__203_0_I2983 (.Y(N9559), .A(N10038), .B(N9670), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2984 (.Y(N10235), .A(N8759), .B(N10094), .S0(N9559));
MXI2XL inst_cellmath__203_0_I2985 (.Y(N9490), .A(N8716), .B(N10038), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2986 (.Y(N8896), .A(N8759), .B(N10094), .S0(N9490));
MXI2XL inst_cellmath__203_0_I2987 (.Y(N9424), .A(N9055), .B(N8716), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2988 (.Y(N9266), .A(N8759), .B(N10094), .S0(N9424));
MXI2XL inst_cellmath__203_0_I2989 (.Y(N9357), .A(N9437), .B(N9055), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2990 (.Y(N9660), .A(N8759), .B(N10094), .S0(N9357));
MXI2XL inst_cellmath__203_0_I2991 (.Y(N9289), .A(N9825), .B(N9437), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2992 (.Y(N10027), .A(N8759), .B(N10094), .S0(N9289));
MXI2XL inst_cellmath__203_0_I2993 (.Y(N9225), .A(N10183), .B(N9825), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2994 (.Y(N8708), .A(N8759), .B(N10094), .S0(N9225));
MXI2XL inst_cellmath__203_0_I2995 (.Y(N9158), .A(N8842), .B(N10183), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2996 (.Y(N9044), .A(N8759), .B(N10094), .S0(N9158));
MXI2XL inst_cellmath__203_0_I2997 (.Y(N9095), .A(N9208), .B(N8842), .S0(N9401));
MXI2XL inst_cellmath__203_0_I2998 (.Y(N9429), .A(N8759), .B(N10094), .S0(N9095));
MXI2XL inst_cellmath__203_0_I2999 (.Y(N9033), .A(N9599), .B(N9208), .S0(N9401));
MXI2XL inst_cellmath__203_0_I3000 (.Y(N9814), .A(N8759), .B(N10094), .S0(N9033));
MXI2XL inst_cellmath__203_0_I3001 (.Y(N8972), .A(N9978), .B(N9599), .S0(N9401));
MXI2XL inst_cellmath__203_0_I3002 (.Y(N10171), .A(N8759), .B(N10094), .S0(N8972));
MXI2XL inst_cellmath__203_0_I3003 (.Y(N8912), .A(N8664), .B(N9978), .S0(N9401));
MXI2XL inst_cellmath__203_0_I3004 (.Y(N8836), .A(N8759), .B(N10094), .S0(N8912));
MXI2XL inst_cellmath__203_0_I3005 (.Y(N8849), .A(N8993), .B(N8664), .S0(N9401));
MXI2XL inst_cellmath__203_0_I3006 (.Y(N9200), .A(N8759), .B(N10094), .S0(N8849));
NOR2BX1 inst_cellmath__203_0_I3007 (.Y(N8794), .AN(N9401), .B(N8993));
MXI2XL inst_cellmath__203_0_I3008 (.Y(N9700), .A(N8759), .B(N10094), .S0(N8794));
XNOR2X1 inst_cellmath__203_0_I3009 (.Y(N9361), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
NOR2XL inst_cellmath__203_0_I3010 (.Y(N9472), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
OAI2BB1X1 inst_cellmath__203_0_I3011 (.Y(N8982), .A0N(inst_cellmath__61[15]), .A1N(inst_cellmath__61[14]), .B0(inst_cellmath__115__W1[0]));
INVXL inst_cellmath__203_0_I3012 (.Y(N9107), .A(N8982));
OR2XL inst_cellmath__203_0_I3013 (.Y(N10239), .A(N9472), .B(inst_cellmath__115__W1[0]));
INVXL inst_cellmath__203_0_I3014 (.Y(inst_cellmath__203__W0[42]), .A(N9107));
NOR2XL inst_cellmath__203_0_I3015 (.Y(N10155), .A(N9736), .B(N9361));
MXI2XL inst_cellmath__203_0_I3016 (.Y(N9905), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N10155));
MXI2XL inst_cellmath__203_0_I3017 (.Y(N10099), .A(N10101), .B(N9736), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3018 (.Y(N10261), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N10099));
MXI2XL inst_cellmath__203_0_I3019 (.Y(N10036), .A(N8766), .B(N10101), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3020 (.Y(N8920), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N10036));
MXI2XL inst_cellmath__203_0_I3021 (.Y(N9976), .A(N9115), .B(N8766), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3022 (.Y(N9295), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9976));
MXI2XL inst_cellmath__203_0_I3023 (.Y(N9915), .A(N9507), .B(N9115), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3024 (.Y(N9685), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9915));
MXI2XL inst_cellmath__203_0_I3025 (.Y(N9854), .A(N9888), .B(N9507), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3026 (.Y(N10051), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9854));
MXI2XL inst_cellmath__203_0_I3027 (.Y(N9788), .A(N10248), .B(N9888), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3028 (.Y(N8732), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9788));
MXI2XL inst_cellmath__203_0_I3029 (.Y(N9728), .A(N8907), .B(N10248), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3030 (.Y(N9070), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9728));
MXI2XL inst_cellmath__203_0_I3031 (.Y(N9662), .A(N9277), .B(N8907), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3032 (.Y(N9457), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9662));
MXI2XL inst_cellmath__203_0_I3033 (.Y(N9592), .A(N9670), .B(N9277), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3034 (.Y(N9844), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9592));
MXI2XL inst_cellmath__203_0_I3035 (.Y(N9528), .A(N10038), .B(N9670), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3036 (.Y(N10199), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9528));
MXI2XL inst_cellmath__203_0_I3037 (.Y(N9459), .A(N8716), .B(N10038), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3038 (.Y(N8859), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9459));
MXI2XL inst_cellmath__203_0_I3039 (.Y(N9394), .A(N9055), .B(N8716), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3040 (.Y(N9230), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9394));
MXI2XL inst_cellmath__203_0_I3041 (.Y(N9327), .A(N9437), .B(N9055), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3042 (.Y(N9618), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9327));
MXI2XL inst_cellmath__203_0_I3043 (.Y(N9259), .A(N9825), .B(N9437), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3044 (.Y(N9991), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9259));
MXI2XL inst_cellmath__203_0_I3045 (.Y(N9194), .A(N10183), .B(N9825), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3046 (.Y(N8679), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9194));
MXI2XL inst_cellmath__203_0_I3047 (.Y(N9128), .A(N8842), .B(N10183), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3048 (.Y(N9010), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9128));
MXI2XL inst_cellmath__203_0_I3049 (.Y(N9067), .A(N9208), .B(N8842), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3050 (.Y(N9392), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9067));
MXI2XL inst_cellmath__203_0_I3051 (.Y(N9005), .A(N9599), .B(N9208), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3052 (.Y(N9779), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N9005));
MXI2XL inst_cellmath__203_0_I3053 (.Y(N8941), .A(N9978), .B(N9599), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3054 (.Y(N10137), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N8941));
MXI2XL inst_cellmath__203_0_I3055 (.Y(N8881), .A(N8664), .B(N9978), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3056 (.Y(N8802), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N8881));
MXI2XL inst_cellmath__203_0_I3057 (.Y(N8822), .A(N8993), .B(N8664), .S0(N9361));
MXI2XL inst_cellmath__203_0_I3058 (.Y(N9163), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N8822));
NOR2BX1 inst_cellmath__203_0_I3059 (.Y(N8770), .AN(N9361), .B(N8993));
MXI2XL inst_cellmath__203_0_I3060 (.Y(inst_cellmath__203__W1[42]), .A(inst_cellmath__203__W0[42]), .B(N10239), .S0(N8770));
ADDHX1 inst_cellmath__203_0_I3061 (.CO(inst_cellmath__203__W0[2]), .S(inst_cellmath__203__W1[1]), .A(N10277), .B(inst_cellmath__198[19]));
ADDHX1 inst_cellmath__203_0_I3062 (.CO(N9546), .S(inst_cellmath__203__W1[2]), .A(N9311), .B(N9366));
ADDHX1 inst_cellmath__203_0_I3063 (.CO(N10281), .S(inst_cellmath__203__W0[3]), .A(N10069), .B(N9759));
ADDFX1 inst_cellmath__203_0_I3064 (.CO(inst_cellmath__203__W0[4]), .S(inst_cellmath__203__W1[3]), .A(N9942), .B(N9768), .CI(N9546));
ADDFX1 inst_cellmath__203_0_I3065 (.CO(N10072), .S(N9710), .A(N9084), .B(N9564), .CI(N10122));
ADDFX1 inst_cellmath__203_0_I3066 (.CO(N9090), .S(inst_cellmath__203__W1[4]), .A(N10281), .B(N10292), .CI(N9710));
ADDFX1 inst_cellmath__203_0_I3067 (.CO(N9863), .S(N9476), .A(N10296), .B(inst_cellmath__61[2]), .CI(N10138));
ADDFX1 inst_cellmath__203_0_I3068 (.CO(N8878), .S(N10222), .A(N9859), .B(N9476), .CI(N8786));
ADDFX1 inst_cellmath__203_0_I3069 (.CO(N9642), .S(inst_cellmath__203__W0[5]), .A(N8952), .B(N9925), .CI(N9133));
ADDFX1 inst_cellmath__203_0_I3070 (.CO(inst_cellmath__203__W0[6]), .S(inst_cellmath__203__W1[5]), .A(N10222), .B(N10072), .CI(N9090));
ADDFX1 inst_cellmath__203_0_I3071 (.CO(N9410), .S(N9030), .A(N8804), .B(N9336), .CI(N9863));
ADDFX1 inst_cellmath__203_0_I3072 (.CO(N10160), .S(N9797), .A(N8874), .B(N9030), .CI(N9139));
ADDFX1 inst_cellmath__203_0_I3073 (.CO(N9182), .S(N8819), .A(N9527), .B(N9334), .CI(N8878));
ADDFX1 inst_cellmath__203_0_I3074 (.CO(inst_cellmath__203__W0[7]), .S(inst_cellmath__203__W1[6]), .A(N9642), .B(N9797), .CI(N8819));
ADDFX1 inst_cellmath__203_0_I3075 (.CO(N8968), .S(N10304), .A(N10091), .B(N9918), .CI(N9165));
ADDFX1 inst_cellmath__203_0_I3076 (.CO(N9737), .S(N9344), .A(N10304), .B(N10112), .CI(N9410));
ADDFX1 inst_cellmath__203_0_I3077 (.CO(N8767), .S(N10104), .A(N9635), .B(N9344), .CI(N9532));
ADDFX1 inst_cellmath__203_0_I3078 (.CO(N9510), .S(N9117), .A(N9725), .B(N10071), .CI(N10078));
ADDFX1 inst_cellmath__203_0_I3079 (.CO(N10250), .S(N9889), .A(N10160), .B(N9903), .CI(N10104));
ADDFX1 inst_cellmath__203_0_I3080 (.CO(inst_cellmath__203__W0[8]), .S(inst_cellmath__203__W1[7]), .A(N9117), .B(N9182), .CI(N9889));
ADDFX1 inst_cellmath__203_0_I3081 (.CO(N10039), .S(N9671), .A(N9557), .B(N9106), .CI(N8777));
ADDFX1 inst_cellmath__203_0_I3082 (.CO(N9057), .S(N8717), .A(N9671), .B(N8968), .CI(N9737));
ADDFX1 inst_cellmath__203_0_I3083 (.CO(N9826), .S(N9440), .A(N8691), .B(N8717), .CI(N9912));
ADDFX1 inst_cellmath__203_0_I3084 (.CO(N8845), .S(N10186), .A(N8749), .B(N10088), .CI(N10262));
ADDFX1 inst_cellmath__203_0_I3085 (.CO(N9602), .S(N9209), .A(N9440), .B(N8767), .CI(N9510));
ADDFX1 inst_cellmath__203_0_I3086 (.CO(inst_cellmath__203__W0[9]), .S(inst_cellmath__203__W1[8]), .A(N10186), .B(N10250), .CI(N9209));
ADDFX1 inst_cellmath__203_0_I3087 (.CO(N9374), .S(N8995), .A(N9882), .B(N10064), .CI(N9934));
ADDFX1 inst_cellmath__203_0_I3088 (.CO(N10127), .S(N9764), .A(N10074), .B(N9130), .CI(N10039));
ADDFX1 inst_cellmath__203_0_I3089 (.CO(N9147), .S(N8791), .A(N9764), .B(N8995), .CI(N9057));
ADDFX1 inst_cellmath__203_0_I3090 (.CO(N9920), .S(N9536), .A(N8791), .B(N9405), .CI(N10268));
ADDFX1 inst_cellmath__203_0_I3091 (.CO(N8932), .S(N10274), .A(N8757), .B(N10219), .CI(N9285));
ADDFX1 inst_cellmath__203_0_I3092 (.CO(N9701), .S(N9308), .A(N8921), .B(N9097), .CI(N9826));
ADDFX1 inst_cellmath__203_0_I3093 (.CO(N8741), .S(N10066), .A(N8845), .B(N9536), .CI(N10274));
ADDFX1 inst_cellmath__203_0_I3094 (.CO(inst_cellmath__203__W0[10]), .S(inst_cellmath__203__W1[9]), .A(N9602), .B(N9308), .CI(N10066));
ADDFX1 inst_cellmath__203_0_I3095 (.CO(N10215), .S(N9858), .A(N9521), .B(N8897), .CI(N8746));
ADDFX1 inst_cellmath__203_0_I3096 (.CO(N9243), .S(N8872), .A(N9374), .B(N10288), .CI(N9858));
ADDFX1 inst_cellmath__203_0_I3097 (.CO(N10005), .S(N9633), .A(N8872), .B(N10127), .CI(N10152));
ADDFX1 inst_cellmath__203_0_I3098 (.CO(N9022), .S(N8688), .A(N9633), .B(N9147), .CI(N8928));
ADDFX1 inst_cellmath__203_0_I3099 (.CO(N9791), .S(N9403), .A(N9678), .B(N9103), .CI(N9485));
ADDFX1 inst_cellmath__203_0_I3100 (.CO(N8813), .S(N10150), .A(N9920), .B(N9293), .CI(N8688));
ADDFX1 inst_cellmath__203_0_I3101 (.CO(N9566), .S(N9172), .A(N9701), .B(N8932), .CI(N9403));
ADDFX1 inst_cellmath__203_0_I3102 (.CO(inst_cellmath__203__W0[11]), .S(inst_cellmath__203__W1[10]), .A(N8741), .B(N10150), .CI(N9172));
ADDFX1 inst_cellmath__203_0_I3103 (.CO(N9337), .S(N8958), .A(N9664), .B(N10213), .CI(N8946));
ADDFX1 inst_cellmath__203_0_I3104 (.CO(N10095), .S(N9730), .A(N9094), .B(N9897), .CI(N10041));
ADDFX1 inst_cellmath__203_0_I3105 (.CO(N9108), .S(N8760), .A(N8958), .B(N10215), .CI(N9730));
ADDFX1 inst_cellmath__203_0_I3106 (.CO(N9884), .S(N9499), .A(N8760), .B(N9243), .CI(N9177));
ADDFX1 inst_cellmath__203_0_I3107 (.CO(N8901), .S(N10240), .A(N9499), .B(N10005), .CI(N9300));
ADDFX1 inst_cellmath__203_0_I3108 (.CO(N9665), .S(N9269), .A(N9494), .B(N8693), .CI(N10046));
ADDFX1 inst_cellmath__203_0_I3109 (.CO(N8713), .S(N10032), .A(N10220), .B(N9870), .CI(N9686));
ADDFX1 inst_cellmath__203_0_I3110 (.CO(N9432), .S(N9048), .A(N10240), .B(N9022), .CI(N9791));
ADDFX1 inst_cellmath__203_0_I3111 (.CO(N10177), .S(N9820), .A(N9269), .B(N8813), .CI(N10032));
ADDFX1 inst_cellmath__203_0_I3112 (.CO(inst_cellmath__203__W0[12]), .S(inst_cellmath__203__W1[11]), .A(N9566), .B(N9048), .CI(N9820));
ADDFX1 inst_cellmath__203_0_I3113 (.CO(N9972), .S(N9594), .A(N9329), .B(N8712), .CI(N9479));
ADDFX1 inst_cellmath__203_0_I3114 (.CO(N8986), .S(N8658), .A(N8720), .B(N10258), .CI(N9337));
ADDFX1 inst_cellmath__203_0_I3115 (.CO(N9757), .S(N9364), .A(N9594), .B(N10095), .CI(N8658));
ADDFX1 inst_cellmath__203_0_I3116 (.CO(N8785), .S(N10117), .A(N9364), .B(N9108), .CI(N9949));
ADDFX1 inst_cellmath__203_0_I3117 (.CO(N9529), .S(N9136), .A(N10117), .B(N9884), .CI(N9694));
ADDFX1 inst_cellmath__203_0_I3118 (.CO(N10265), .S(N9910), .A(N8725), .B(N9879), .CI(N8879));
ADDFX1 inst_cellmath__203_0_I3119 (.CO(N9298), .S(N8924), .A(N10052), .B(N10227), .CI(N8901));
ADDFX1 inst_cellmath__203_0_I3120 (.CO(N10056), .S(N9691), .A(N9665), .B(N9136), .CI(N8713));
ADDFX1 inst_cellmath__203_0_I3121 (.CO(N9074), .S(N8735), .A(N8924), .B(N9910), .CI(N9432));
ADDFX1 inst_cellmath__203_0_I3122 (.CO(inst_cellmath__203__W0[13]), .S(inst_cellmath__203__W1[12]), .A(N10177), .B(N9691), .CI(N8735));
ADDFX1 inst_cellmath__203_0_I3123 (.CO(N8863), .S(N10203), .A(N9430), .B(N8687), .CI(N8917));
ADDFX1 inst_cellmath__203_0_I3124 (.CO(N9625), .S(N9234), .A(N9060), .B(N9865), .CI(N9719));
ADDFX1 inst_cellmath__203_0_I3125 (.CO(N8681), .S(N9996), .A(N9972), .B(N10007), .CI(N10203));
ADDFX1 inst_cellmath__203_0_I3126 (.CO(N9397), .S(N9015), .A(N8986), .B(N9234), .CI(N9996));
ADDFX1 inst_cellmath__203_0_I3127 (.CO(N10143), .S(N9784), .A(N9015), .B(N9757), .CI(N8960));
ADDFX1 inst_cellmath__203_0_I3128 (.CO(N9167), .S(N8806), .A(N9784), .B(N8785), .CI(N10060));
ADDFX1 inst_cellmath__203_0_I3129 (.CO(N9936), .S(N9562), .A(N9066), .B(N10236), .CI(N9249));
ADDFX1 inst_cellmath__203_0_I3130 (.CO(N8950), .S(N10290), .A(N8886), .B(N8817), .CI(N8729));
ADDFX1 inst_cellmath__203_0_I3131 (.CO(N9722), .S(N9330), .A(N9438), .B(N9529), .CI(N8806));
ADDFX1 inst_cellmath__203_0_I3132 (.CO(N8752), .S(N10085), .A(N9298), .B(N10265), .CI(N9562));
ADDFX1 inst_cellmath__203_0_I3133 (.CO(N9492), .S(N9101), .A(N10056), .B(N10290), .CI(N9330));
ADDFX1 inst_cellmath__203_0_I3134 (.CO(inst_cellmath__203__W0[14]), .S(inst_cellmath__203__W1[13]), .A(N10085), .B(N9074), .CI(N9101));
ADDFX1 inst_cellmath__203_0_I3135 (.CO(N9263), .S(N8892), .A(N9287), .B(N10175), .CI(N9442));
ADDFX1 inst_cellmath__203_0_I3136 (.CO(N10023), .S(N9657), .A(N8690), .B(N10224), .CI(N10080));
ADDFX1 inst_cellmath__203_0_I3137 (.CO(N9042), .S(N8705), .A(N9625), .B(N8863), .CI(N8892));
ADDFX1 inst_cellmath__203_0_I3138 (.CO(N9811), .S(N9426), .A(N8681), .B(N9657), .CI(N8705));
ADDFX1 inst_cellmath__203_0_I3139 (.CO(N8832), .S(N10169), .A(N9734), .B(N9397), .CI(N9426));
ADDFX1 inst_cellmath__203_0_I3140 (.CO(N9589), .S(N9198), .A(N10169), .B(N10143), .CI(N8736));
ADDFX1 inst_cellmath__203_0_I3141 (.CO(N8652), .S(N9964), .A(N9448), .B(N8893), .CI(N9640));
ADDFX1 inst_cellmath__203_0_I3142 (.CO(N9359), .S(N8980), .A(N9071), .B(N9258), .CI(N9167));
ADDFX1 inst_cellmath__203_0_I3143 (.CO(N10114), .S(N9750), .A(N9198), .B(N9827), .CI(N9936));
ADDFX1 inst_cellmath__203_0_I3144 (.CO(N9131), .S(N8780), .A(N9964), .B(N8950), .CI(N9722));
ADDFX1 inst_cellmath__203_0_I3145 (.CO(N9901), .S(N9524), .A(N9750), .B(N8980), .CI(N8752));
ADDFX1 inst_cellmath__203_0_I3146 (.CO(inst_cellmath__203__W0[15]), .S(inst_cellmath__203__W1[14]), .A(N8780), .B(N9492), .CI(N9524));
ADDHX1 inst_cellmath__203_0_I3147 (.CO(N9683), .S(N9292), .A(N8812), .B(N9203));
ADDFX1 inst_cellmath__203_0_I3148 (.CO(N8728), .S(N10049), .A(N8882), .B(N9292), .CI(N8750));
ADDFX1 inst_cellmath__203_0_I3149 (.CO(N9454), .S(N9069), .A(N9025), .B(N9828), .CI(N9681));
ADDFX1 inst_cellmath__203_0_I3150 (.CO(N10197), .S(N9840), .A(N9263), .B(N9975), .CI(N10023));
ADDFX1 inst_cellmath__203_0_I3151 (.CO(N9227), .S(N8857), .A(N9069), .B(N10049), .CI(N9042));
ADDFX1 inst_cellmath__203_0_I3152 (.CO(N9988), .S(N9615), .A(N8857), .B(N9840), .CI(N9811));
ADDFX1 inst_cellmath__203_0_I3153 (.CO(N9008), .S(N8675), .A(N8832), .B(N8763), .CI(N9615));
ADDFX1 inst_cellmath__203_0_I3154 (.CO(N9776), .S(N9389), .A(N10149), .B(N8675), .CI(N9076));
ADDFX1 inst_cellmath__203_0_I3155 (.CO(N8800), .S(N10135), .A(N9833), .B(N9267), .CI(N10010));
ADDFX1 inst_cellmath__203_0_I3156 (.CO(N9552), .S(N9160), .A(N9458), .B(N9649), .CI(N9589));
ADDFX1 inst_cellmath__203_0_I3157 (.CO(N10284), .S(N9930), .A(N9389), .B(N10187), .CI(N8652));
ADDFX1 inst_cellmath__203_0_I3158 (.CO(N9324), .S(N8943), .A(N10135), .B(N9359), .CI(N9160));
ADDFX1 inst_cellmath__203_0_I3159 (.CO(N10076), .S(N9714), .A(N9930), .B(N10114), .CI(N9131));
ADDFX1 inst_cellmath__203_0_I3160 (.CO(inst_cellmath__203__W0[16]), .S(inst_cellmath__203__W1[15]), .A(N9901), .B(N8943), .CI(N9714));
ADDFX1 inst_cellmath__203_0_I3161 (.CO(N9866), .S(N9482), .A(N9683), .B(N9969), .CI(N9252));
ADDFX1 inst_cellmath__203_0_I3162 (.CO(N8884), .S(N10226), .A(N9404), .B(N9099), .CI(N10048));
ADDFX1 inst_cellmath__203_0_I3163 (.CO(N9647), .S(N9254), .A(N8660), .B(N10189), .CI(N8728));
ADDFX1 inst_cellmath__203_0_I3164 (.CO(N8697), .S(N10015), .A(N9482), .B(N9454), .CI(N10226));
ADDFX1 inst_cellmath__203_0_I3165 (.CO(N9417), .S(N9035), .A(N9254), .B(N10197), .CI(N10015));
ADDFX1 inst_cellmath__203_0_I3166 (.CO(N10163), .S(N9802), .A(N9501), .B(N9227), .CI(N9035));
ADDFX1 inst_cellmath__203_0_I3167 (.CO(N9188), .S(N8826), .A(N9802), .B(N9988), .CI(N9008));
ADDFX1 inst_cellmath__203_0_I3168 (.CO(N9958), .S(N9579), .A(N9464), .B(N9173), .CI(N8826));
ADDFX1 inst_cellmath__203_0_I3169 (.CO(N8974), .S(N10308), .A(N10193), .B(N9661), .CI(N8695));
ADDFX1 inst_cellmath__203_0_I3170 (.CO(N9742), .S(N9351), .A(N9842), .B(N10016), .CI(N9776));
ADDFX1 inst_cellmath__203_0_I3171 (.CO(N8773), .S(N10106), .A(N9579), .B(N8843), .CI(N8800));
ADDFX1 inst_cellmath__203_0_I3172 (.CO(N9514), .S(N9123), .A(N10308), .B(N9552), .CI(N9351));
ADDFX1 inst_cellmath__203_0_I3173 (.CO(N10253), .S(N9893), .A(N10106), .B(N10284), .CI(N9324));
ADDFX1 inst_cellmath__203_0_I3174 (.CO(inst_cellmath__203__W0[17]), .S(inst_cellmath__203__W1[16]), .A(N10076), .B(N9123), .CI(N9893));
ADDFX1 inst_cellmath__203_0_I3175 (.CO(N10042), .S(N9674), .A(N8985), .B(N8956), .CI(N9488));
ADDFX1 inst_cellmath__203_0_I3176 (.CO(N9062), .S(N8723), .A(N8727), .B(N8848), .CI(N9793));
ADDFX1 inst_cellmath__203_0_I3177 (.CO(N9831), .S(N9444), .A(N9941), .B(N8989), .CI(N9644));
ADDFX1 inst_cellmath__203_0_I3178 (.CO(N8850), .S(N10190), .A(N8884), .B(N9866), .CI(N9674));
ADDFX1 inst_cellmath__203_0_I3179 (.CO(N9607), .S(N9217), .A(N9444), .B(N8723), .CI(N9647));
ADDFX1 inst_cellmath__203_0_I3180 (.CO(N8668), .S(N9982), .A(N10190), .B(N8697), .CI(N9217));
ADDFX1 inst_cellmath__203_0_I3181 (.CO(N9379), .S(N9000), .A(N10245), .B(N9417), .CI(N9982));
ADDFX1 inst_cellmath__203_0_I3182 (.CO(N10130), .S(N9767), .A(N9000), .B(N10163), .CI(N9947));
ADDFX1 inst_cellmath__203_0_I3183 (.CO(N9151), .S(N8795), .A(N9851), .B(N9188), .CI(N10025));
ADDFX1 inst_cellmath__203_0_I3184 (.CO(N9924), .S(N9543), .A(N8700), .B(N8853), .CI(N10200));
ADDFX1 inst_cellmath__203_0_I3185 (.CO(N8938), .S(N10279), .A(N9767), .B(N9029), .CI(N9958));
ADDFX1 inst_cellmath__203_0_I3186 (.CO(N9705), .S(N9315), .A(N8795), .B(N9210), .CI(N8974));
ADDFX1 inst_cellmath__203_0_I3187 (.CO(N8743), .S(N10070), .A(N10279), .B(N9742), .CI(N9543));
ADDFX1 inst_cellmath__203_0_I3188 (.CO(N9473), .S(N9087), .A(N9315), .B(N8773), .CI(N9514));
ADDFX1 inst_cellmath__203_0_I3189 (.CO(inst_cellmath__203__W0[18]), .S(inst_cellmath__203__W1[17]), .A(N10253), .B(N10070), .CI(N9087));
ADDFX1 inst_cellmath__203_0_I3190 (.CO(N9247), .S(N8876), .A(N9213), .B(N9755), .CI(N10154));
ADDFX1 inst_cellmath__203_0_I3191 (.CO(N10008), .S(N9638), .A(N9368), .B(N9068), .CI(N10294));
ADDFX1 inst_cellmath__203_0_I3192 (.CO(N9027), .S(N8692), .A(N10012), .B(N9873), .CI(N10042));
ADDFX1 inst_cellmath__203_0_I3193 (.CO(N9794), .S(N9408), .A(N9831), .B(N9062), .CI(N8876));
ADDFX1 inst_cellmath__203_0_I3194 (.CO(N8816), .S(N10156), .A(N8692), .B(N9638), .CI(N8850));
ADDFX1 inst_cellmath__203_0_I3195 (.CO(N9571), .S(N9179), .A(N9408), .B(N9607), .CI(N10156));
ADDFX1 inst_cellmath__203_0_I3196 (.CO(N10301), .S(N9951), .A(N9272), .B(N8668), .CI(N9179));
ADDFX1 inst_cellmath__203_0_I3197 (.CO(N9341), .S(N8963), .A(N9951), .B(N9379), .CI(N8957));
ADDFX1 inst_cellmath__203_0_I3198 (.CO(N10100), .S(N9735), .A(N8709), .B(N10207), .CI(N10130));
ADDFX1 inst_cellmath__203_0_I3199 (.CO(N9113), .S(N8765), .A(N9036), .B(N9220), .CI(N8860));
ADDFX1 inst_cellmath__203_0_I3200 (.CO(N9887), .S(N9505), .A(N8963), .B(N9411), .CI(N9603));
ADDFX1 inst_cellmath__203_0_I3201 (.CO(N8905), .S(N10247), .A(N8938), .B(N9151), .CI(N9735));
ADDFX1 inst_cellmath__203_0_I3202 (.CO(N9669), .S(N9276), .A(N8765), .B(N9924), .CI(N9505));
ADDFX1 inst_cellmath__203_0_I3203 (.CO(N8715), .S(N10037), .A(N8743), .B(N9705), .CI(N10247));
ADDFX1 inst_cellmath__203_0_I3204 (.CO(inst_cellmath__203__W0[19]), .S(inst_cellmath__203__W1[18]), .A(N9473), .B(N9276), .CI(N10037));
ADDFX1 inst_cellmath__203_0_I3205 (.CO(N10182), .S(N9824), .A(N8784), .B(N9107), .CI(N9451));
ADDFX1 inst_cellmath__203_0_I3206 (.CO(N9207), .S(N8841), .A(N8696), .B(N8814), .CI(N9758));
ADDFX1 inst_cellmath__203_0_I3207 (.CO(N9977), .S(N9598), .A(N10232), .B(N8951), .CI(N9605));
ADDFX1 inst_cellmath__203_0_I3208 (.CO(N8991), .S(N8663), .A(N9247), .B(N9905), .CI(N10008));
ADDFX1 inst_cellmath__203_0_I3209 (.CO(N9761), .S(N9370), .A(N8841), .B(N9824), .CI(N9027));
ADDFX1 inst_cellmath__203_0_I3210 (.CO(N8789), .S(N10124), .A(N9794), .B(N9598), .CI(N8663));
ADDFX1 inst_cellmath__203_0_I3211 (.CO(N9533), .S(N9143), .A(N8816), .B(N9370), .CI(N10124));
ADDFX1 inst_cellmath__203_0_I3212 (.CO(N10271), .S(N9917), .A(N9571), .B(N10034), .CI(N9143));
ADDFX1 inst_cellmath__203_0_I3213 (.CO(N9305), .S(N8930), .A(N9917), .B(N10301), .CI(N9731));
ADDFX1 inst_cellmath__203_0_I3214 (.CO(N10062), .S(N9697), .A(N9045), .B(N8868), .CI(N9341));
ADDFX1 inst_cellmath__203_0_I3215 (.CO(N9081), .S(N8740), .A(N9419), .B(N9609), .CI(N9228));
ADDFX1 inst_cellmath__203_0_I3216 (.CO(N9856), .S(N9465), .A(N8930), .B(N9798), .CI(N9979));
ADDFX1 inst_cellmath__203_0_I3217 (.CO(N8870), .S(N10211), .A(N9113), .B(N10100), .CI(N9697));
ADDFX1 inst_cellmath__203_0_I3218 (.CO(N9631), .S(N9241), .A(N8740), .B(N9887), .CI(N9465));
ADDFX1 inst_cellmath__203_0_I3219 (.CO(N8685), .S(N10001), .A(N10211), .B(N8905), .CI(N9669));
ADDFX1 inst_cellmath__203_0_I3220 (.CO(inst_cellmath__203__W0[20]), .S(inst_cellmath__203__W1[19]), .A(N8715), .B(N9241), .CI(N10001));
INVXL inst_cellmath__203_0_I3221 (.Y(N8719), .A(N9171));
ADDFX1 inst_cellmath__203_0_I3222 (.CO(N10146), .S(N9789), .A(N9032), .B(N9176), .CI(N8719));
ADDFX1 inst_cellmath__203_0_I3223 (.CO(N9944), .S(N9565), .A(N10121), .B(N9333), .CI(N9981));
ADDFX1 inst_cellmath__203_0_I3224 (.CO(N8955), .S(N10295), .A(N10261), .B(N8888), .CI(N9836));
ADDFX1 inst_cellmath__203_0_I3225 (.CO(N9729), .S(N9335), .A(N9207), .B(N10182), .CI(N9977));
ADDFX1 inst_cellmath__203_0_I3226 (.CO(N8758), .S(N10092), .A(N9565), .B(N9789), .CI(N10295));
ADDFX1 inst_cellmath__203_0_I3227 (.CO(N9497), .S(N9105), .A(N9761), .B(N8991), .CI(N9335));
ADDFX1 inst_cellmath__203_0_I3228 (.CO(N10237), .S(N9881), .A(N8789), .B(N10092), .CI(N9105));
ADDFX1 inst_cellmath__203_0_I3229 (.CO(N9268), .S(N8899), .A(N9533), .B(N9219), .CI(N9881));
ADDFX1 inst_cellmath__203_0_I3230 (.CO(N10029), .S(N9663), .A(N8899), .B(N10271), .CI(N8761));
ADDFX1 inst_cellmath__203_0_I3231 (.CO(N9047), .S(N8711), .A(N9427), .B(N9236), .CI(N9305));
ADDFX1 inst_cellmath__203_0_I3232 (.CO(N9818), .S(N9431), .A(N9805), .B(N9984), .CI(N9619));
ADDFX1 inst_cellmath__203_0_I3233 (.CO(N8838), .S(N10174), .A(N9663), .B(N10158), .CI(N8665));
ADDFX1 inst_cellmath__203_0_I3234 (.CO(N9593), .S(N9202), .A(N9081), .B(N10062), .CI(N8711));
ADDFX1 inst_cellmath__203_0_I3235 (.CO(N8657), .S(N9970), .A(N9431), .B(N9856), .CI(N10174));
ADDFX1 inst_cellmath__203_0_I3236 (.CO(N9362), .S(N8984), .A(N9202), .B(N8870), .CI(N9631));
ADDFX1 inst_cellmath__203_0_I3237 (.CO(inst_cellmath__203__W0[21]), .S(inst_cellmath__203__W1[20]), .A(N8685), .B(N9970), .CI(N8984));
INVXL inst_cellmath__203_0_I3238 (.Y(N8666), .A(N9907));
ADDFX1 inst_cellmath__203_0_I3239 (.CO(N9135), .S(N8783), .A(N9413), .B(N9171), .CI(N8666));
ADDFX1 inst_cellmath__203_0_I3240 (.CO(N8922), .S(N10264), .A(N9261), .B(N8787), .CI(N9727));
ADDFX1 inst_cellmath__203_0_I3241 (.CO(N9689), .S(N9296), .A(N8920), .B(N8667), .CI(N9568));
ADDFX1 inst_cellmath__203_0_I3242 (.CO(N8733), .S(N10054), .A(N10146), .B(N10195), .CI(N9944));
ADDFX1 inst_cellmath__203_0_I3243 (.CO(N9460), .S(N9073), .A(N8783), .B(N8955), .CI(N10264));
ADDFX1 inst_cellmath__203_0_I3244 (.CO(N10202), .S(N9846), .A(N9729), .B(N9296), .CI(N10054));
ADDFX1 inst_cellmath__203_0_I3245 (.CO(N9231), .S(N8861), .A(N9073), .B(N8758), .CI(N9497));
ADDFX1 inst_cellmath__203_0_I3246 (.CO(N9994), .S(N9623), .A(N8861), .B(N9846), .CI(N10237));
ADDFX1 inst_cellmath__203_0_I3247 (.CO(N9013), .S(N8680), .A(N9268), .B(N9623), .CI(N9498));
ADDFX1 inst_cellmath__203_0_I3248 (.CO(N9781), .S(N9395), .A(N9815), .B(N9628), .CI(N10029));
ADDFX1 inst_cellmath__203_0_I3249 (.CO(N8803), .S(N10139), .A(N10164), .B(N8670), .CI(N9992));
ADDFX1 inst_cellmath__203_0_I3250 (.CO(N9558), .S(N9164), .A(N8680), .B(N8820), .CI(N8996));
ADDFX1 inst_cellmath__203_0_I3251 (.CO(N10287), .S(N9933), .A(N9818), .B(N9047), .CI(N9395));
ADDFX1 inst_cellmath__203_0_I3252 (.CO(N9328), .S(N8947), .A(N10139), .B(N8838), .CI(N9164));
ADDFX1 inst_cellmath__203_0_I3253 (.CO(N10082), .S(N9718), .A(N9933), .B(N9593), .CI(N8657));
ADDFX1 inst_cellmath__203_0_I3254 (.CO(inst_cellmath__203__W0[22]), .S(inst_cellmath__203__W1[21]), .A(N9362), .B(N8947), .CI(N9718));
ADDFX1 inst_cellmath__203_0_I3255 (.CO(N9872), .S(N9489), .A(N9297), .B(N9907), .CI(N9654));
ADDFX1 inst_cellmath__203_0_I3256 (.CO(N8890), .S(N10231), .A(N8998), .B(N9138), .CI(N10087));
ADDFX1 inst_cellmath__203_0_I3257 (.CO(N9653), .S(N9260), .A(N8855), .B(N9295), .CI(N9948));
ADDFX1 inst_cellmath__203_0_I3258 (.CO(N8701), .S(N10021), .A(N9135), .B(N9800), .CI(N8922));
ADDFX1 inst_cellmath__203_0_I3259 (.CO(N9423), .S(N9039), .A(N9489), .B(N9689), .CI(N10231));
ADDFX1 inst_cellmath__203_0_I3260 (.CO(N10167), .S(N9807), .A(N8733), .B(N9260), .CI(N9460));
ADDFX1 inst_cellmath__203_0_I3261 (.CO(N9195), .S(N8830), .A(N9039), .B(N10021), .CI(N10202));
ADDFX1 inst_cellmath__203_0_I3262 (.CO(N9962), .S(N9585), .A(N9231), .B(N9807), .CI(N8830));
ADDFX1 inst_cellmath__203_0_I3263 (.CO(N8978), .S(N8650), .A(N9585), .B(N9994), .CI(N9001));
ADDFX1 inst_cellmath__203_0_I3264 (.CO(N9748), .S(N9356), .A(N8650), .B(N10241), .CI(N10172));
ADDFX1 inst_cellmath__203_0_I3265 (.CO(N8778), .S(N10111), .A(N9003), .B(N9013), .CI(N9183));
ADDFX1 inst_cellmath__203_0_I3266 (.CO(N9520), .S(N9129), .A(N8676), .B(N8827), .CI(N9375));
ADDFX1 inst_cellmath__203_0_I3267 (.CO(N10257), .S(N9899), .A(N9356), .B(N9781), .CI(N8803));
ADDFX1 inst_cellmath__203_0_I3268 (.CO(N9288), .S(N8916), .A(N10111), .B(N9558), .CI(N9129));
ADDFX1 inst_cellmath__203_0_I3269 (.CO(N10047), .S(N9680), .A(N9899), .B(N10287), .CI(N9328));
ADDFX1 inst_cellmath__203_0_I3270 (.CO(inst_cellmath__203__W0[23]), .S(inst_cellmath__203__W1[22]), .A(N10082), .B(N8916), .CI(N9680));
INVXL inst_cellmath__203_0_I3271 (.Y(N10275), .A(N8854));
ADDFX1 inst_cellmath__203_0_I3272 (.CO(N9838), .S(N9450), .A(N10018), .B(N9377), .CI(N10275));
ADDFX1 inst_cellmath__203_0_I3273 (.CO(N9612), .S(N9224), .A(N9223), .B(N8756), .CI(N9685));
ADDFX1 inst_cellmath__203_0_I3274 (.CO(N8672), .S(N9985), .A(N10161), .B(N10300), .CI(N9531));
ADDFX1 inst_cellmath__203_0_I3275 (.CO(N9385), .S(N9006), .A(N8890), .B(N9872), .CI(N9653));
ADDFX1 inst_cellmath__203_0_I3276 (.CO(N10134), .S(N9773), .A(N9224), .B(N9450), .CI(N9985));
ADDFX1 inst_cellmath__203_0_I3277 (.CO(N9156), .S(N8798), .A(N9423), .B(N8701), .CI(N9006));
ADDFX1 inst_cellmath__203_0_I3278 (.CO(N9928), .S(N9551), .A(N10167), .B(N9773), .CI(N8798));
ADDFX1 inst_cellmath__203_0_I3279 (.CO(N8942), .S(N10282), .A(N9551), .B(N9195), .CI(N9962));
ADDFX1 inst_cellmath__203_0_I3280 (.CO(N9711), .S(N9321), .A(N10282), .B(N9270), .CI(N8978));
ADDFX1 inst_cellmath__203_0_I3281 (.CO(N8745), .S(N10075), .A(N9383), .B(N8833), .CI(N9572));
ADDFX1 inst_cellmath__203_0_I3282 (.CO(N9480), .S(N9093), .A(N9011), .B(N9192), .CI(N9321));
ADDFX1 inst_cellmath__203_0_I3283 (.CO(N10223), .S(N9864), .A(N9748), .B(N9762), .CI(N8778));
ADDFX1 inst_cellmath__203_0_I3284 (.CO(N9251), .S(N8883), .A(N10075), .B(N9520), .CI(N9093));
ADDFX1 inst_cellmath__203_0_I3285 (.CO(N10013), .S(N9643), .A(N9864), .B(N10257), .CI(N9288));
ADDFX1 inst_cellmath__203_0_I3286 (.CO(inst_cellmath__203__W0[24]), .S(inst_cellmath__203__W1[23]), .A(N10047), .B(N8883), .CI(N9643));
INVXL inst_cellmath__203_0_I3287 (.Y(N10216), .A(N8824));
ADDFX1 inst_cellmath__203_0_I3288 (.CO(N9799), .S(N9414), .A(N8702), .B(N8854), .CI(N10216));
ADDFX1 inst_cellmath__203_0_I3289 (.CO(N9575), .S(N9185), .A(N9102), .B(N9613), .CI(N10051));
ADDFX1 inst_cellmath__203_0_I3290 (.CO(N10306), .S(N9956), .A(N8823), .B(N8961), .CI(N9914));
ADDFX1 inst_cellmath__203_0_I3291 (.CO(N9348), .S(N8970), .A(N9838), .B(N9765), .CI(N9612));
ADDFX1 inst_cellmath__203_0_I3292 (.CO(N10105), .S(N9739), .A(N9414), .B(N8672), .CI(N9185));
ADDFX1 inst_cellmath__203_0_I3293 (.CO(N9120), .S(N8771), .A(N9385), .B(N9956), .CI(N8970));
ADDFX1 inst_cellmath__203_0_I3294 (.CO(N9891), .S(N9511), .A(N9739), .B(N10134), .CI(N9156));
ADDFX1 inst_cellmath__203_0_I3295 (.CO(N8911), .S(N10252), .A(N9511), .B(N8771), .CI(N9928));
ADDFX1 inst_cellmath__203_0_I3296 (.CO(N9672), .S(N9280), .A(N8942), .B(N10252), .CI(N9153));
ADDFX1 inst_cellmath__203_0_I3297 (.CO(N8721), .S(N10040), .A(N9711), .B(N10031), .CI(N9280));
ADDFX1 inst_cellmath__203_0_I3298 (.CO(N9441), .S(N9059), .A(N9581), .B(N9769), .CI(N9393));
ADDFX1 inst_cellmath__203_0_I3299 (.CO(N10188), .S(N9829), .A(N10128), .B(N9953), .CI(N10040));
ADDFX1 inst_cellmath__203_0_I3300 (.CO(N9215), .S(N8847), .A(N9480), .B(N8745), .CI(N9059));
ADDFX1 inst_cellmath__203_0_I3301 (.CO(N9980), .S(N9604), .A(N9829), .B(N10223), .CI(N9251));
ADDFX1 inst_cellmath__203_0_I3302 (.CO(inst_cellmath__203__W0[25]), .S(inst_cellmath__203__W1[24]), .A(N10013), .B(N8847), .CI(N9604));
XNOR2X1 inst_cellmath__203_0_I3303 (.Y(N9376), .A(N9847), .B(N8824));
OR2XL inst_cellmath__203_0_I3304 (.Y(N9766), .A(N9847), .B(N8824));
ADDFX1 inst_cellmath__203_0_I3305 (.CO(N9540), .S(N9149), .A(N9338), .B(N9376), .CI(N8732));
ADDFX1 inst_cellmath__203_0_I3306 (.CO(N10278), .S(N9922), .A(N9986), .B(N9040), .CI(N9186));
ADDFX1 inst_cellmath__203_0_I3307 (.CO(N9312), .S(N8935), .A(N10129), .B(N10267), .CI(N9493));
ADDFX1 inst_cellmath__203_0_I3308 (.CO(N10068), .S(N9703), .A(N9575), .B(N9799), .CI(N10306));
ADDFX1 inst_cellmath__203_0_I3309 (.CO(N9085), .S(N8742), .A(N9922), .B(N9149), .CI(N8935));
ADDFX1 inst_cellmath__203_0_I3310 (.CO(N9860), .S(N9469), .A(N10105), .B(N9348), .CI(N9703));
ADDFX1 inst_cellmath__203_0_I3311 (.CO(N8873), .S(N10218), .A(N9120), .B(N8742), .CI(N9469));
ADDFX1 inst_cellmath__203_0_I3312 (.CO(N9636), .S(N9245), .A(N10218), .B(N9891), .CI(N8911));
ADDFX1 inst_cellmath__203_0_I3313 (.CO(N8689), .S(N10006), .A(N9245), .B(N9049), .CI(N9672));
ADDFX1 inst_cellmath__203_0_I3314 (.CO(N9407), .S(N9024), .A(N9959), .B(N10131), .CI(N9778));
ADDFX1 inst_cellmath__203_0_I3315 (.CO(N10153), .S(N9792), .A(N8792), .B(N10305), .CI(N10006));
ADDFX1 inst_cellmath__203_0_I3316 (.CO(N9175), .S(N8815), .A(N9441), .B(N8721), .CI(N9024));
ADDFX1 inst_cellmath__203_0_I3317 (.CO(N9950), .S(N9567), .A(N9792), .B(N10188), .CI(N9215));
ADDFX1 inst_cellmath__203_0_I3318 (.CO(inst_cellmath__203__W0[26]), .S(inst_cellmath__203__W1[25]), .A(N9980), .B(N8815), .CI(N9567));
ADDHX1 inst_cellmath__203_0_I3319 (.CO(N9732), .S(N9340), .A(N9766), .B(N9421));
ADDFX1 inst_cellmath__203_0_I3320 (.CO(N8764), .S(N10097), .A(N9576), .B(N8673), .CI(N9340));
ADDFX1 inst_cellmath__203_0_I3321 (.CO(N9502), .S(N9110), .A(N8927), .B(N9070), .CI(N8793));
ADDFX1 inst_cellmath__203_0_I3322 (.CO(N10243), .S(N9886), .A(N9878), .B(N9733), .CI(N9540));
ADDFX1 inst_cellmath__203_0_I3323 (.CO(N9274), .S(N8903), .A(N9312), .B(N10278), .CI(N10097));
ADDFX1 inst_cellmath__203_0_I3324 (.CO(N10035), .S(N9666), .A(N10068), .B(N9110), .CI(N9886));
ADDFX1 inst_cellmath__203_0_I3325 (.CO(N9051), .S(N8714), .A(N8903), .B(N9085), .CI(N9860));
ADDFX1 inst_cellmath__203_0_I3326 (.CO(N9823), .S(N9434), .A(N8873), .B(N9666), .CI(N8714));
ADDFX1 inst_cellmath__203_0_I3327 (.CO(N8840), .S(N10179), .A(N9636), .B(N9434), .CI(N9821));
ADDFX1 inst_cellmath__203_0_I3328 (.CO(N9597), .S(N9205), .A(N8797), .B(N9317), .CI(N8966));
ADDFX1 inst_cellmath__203_0_I3329 (.CO(N8661), .S(N9974), .A(N10179), .B(N8649), .CI(N8689));
ADDFX1 inst_cellmath__203_0_I3330 (.CO(N9367), .S(N8988), .A(N9407), .B(N9145), .CI(N9205));
ADDFX1 inst_cellmath__203_0_I3331 (.CO(N10120), .S(N9760), .A(N10153), .B(N9974), .CI(N9175));
ADDFX1 inst_cellmath__203_0_I3332 (.CO(inst_cellmath__203__W0[27]), .S(inst_cellmath__203__W1[26]), .A(N9950), .B(N8988), .CI(N9760));
XNOR2X1 inst_cellmath__203_0_I3333 (.Y(N9530), .A(N9808), .B(N9302));
OR2XL inst_cellmath__203_0_I3334 (.Y(N9913), .A(N9808), .B(N9302));
ADDFX1 inst_cellmath__203_0_I3335 (.CO(N9695), .S(N9301), .A(N9955), .B(N9007), .CI(N9148));
ADDFX1 inst_cellmath__203_0_I3336 (.CO(N8737), .S(N10058), .A(N10235), .B(N9732), .CI(N10098));
ADDFX1 inst_cellmath__203_0_I3337 (.CO(N9462), .S(N9078), .A(N9530), .B(N9457), .CI(N8764));
ADDFX1 inst_cellmath__203_0_I3338 (.CO(N10208), .S(N9852), .A(N9301), .B(N9502), .CI(N10058));
ADDFX1 inst_cellmath__203_0_I3339 (.CO(N9237), .S(N8866), .A(N9274), .B(N10243), .CI(N9078));
ADDFX1 inst_cellmath__203_0_I3340 (.CO(N9999), .S(N9629), .A(N10035), .B(N9852), .CI(N8866));
ADDFX1 inst_cellmath__203_0_I3341 (.CO(N9019), .S(N8683), .A(N9629), .B(N9051), .CI(N9823));
ADDFX1 inst_cellmath__203_0_I3342 (.CO(N9787), .S(N9400), .A(N8683), .B(N8839), .CI(N8840));
ADDFX1 inst_cellmath__203_0_I3343 (.CO(N8810), .S(N10144), .A(N8976), .B(N9154), .CI(N9345));
ADDFX1 inst_cellmath__203_0_I3344 (.CO(N9563), .S(N9169), .A(N9400), .B(N9537), .CI(N9597));
ADDFX1 inst_cellmath__203_0_I3345 (.CO(N10293), .S(N9940), .A(N10144), .B(N8661), .CI(N9169));
ADDFX1 inst_cellmath__203_0_I3346 (.CO(inst_cellmath__203__W0[28]), .S(inst_cellmath__203__W1[27]), .A(N10120), .B(N9367), .CI(N9940));
ADDFX1 inst_cellmath__203_0_I3348 (.CO(N10089), .S(N9726), .A(N10307), .B(N9386), .CI(N7517));
ADDFX1 inst_cellmath__203_0_I3349 (.CO(N9877), .S(N9496), .A(N8896), .B(N9541), .CI(N8762));
ADDFX1 inst_cellmath__203_0_I3350 (.CO(N8895), .S(N10234), .A(N9844), .B(N9693), .CI(N9913));
ADDFX1 inst_cellmath__203_0_I3351 (.CO(N9659), .S(N9265), .A(N8737), .B(N9695), .CI(N9726));
ADDFX1 inst_cellmath__203_0_I3352 (.CO(N8710), .S(N10026), .A(N10234), .B(N9496), .CI(N9462));
ADDFX1 inst_cellmath__203_0_I3353 (.CO(N9428), .S(N9043), .A(N9265), .B(N10208), .CI(N10026));
ADDFX1 inst_cellmath__203_0_I3354 (.CO(N10170), .S(N9816), .A(N9043), .B(N9237), .CI(N9999));
ADDFX1 inst_cellmath__203_0_I3355 (.CO(N9201), .S(N8835), .A(N9019), .B(N9816), .CI(N9475));
ADDFX1 inst_cellmath__203_0_I3356 (.CO(N9967), .S(N9591), .A(N8835), .B(N9595), .CI(N9547));
ADDFX1 inst_cellmath__203_0_I3357 (.CO(N8981), .S(N8656), .A(N9787), .B(N9738), .CI(N9921));
ADDFX1 inst_cellmath__203_0_I3358 (.CO(N9753), .S(N9360), .A(N9591), .B(N8810), .CI(N8656));
ADDFX1 inst_cellmath__203_0_I3359 (.CO(inst_cellmath__203__W0[29]), .S(inst_cellmath__203__W1[28]), .A(N10293), .B(N9563), .CI(N9360));
ADDFX1 inst_cellmath__203_0_I3360 (.CO(N9526), .S(N9134), .A(N9774), .B(N7696), .CI(N9266));
ADDFX1 inst_cellmath__203_0_I3361 (.CO(N10263), .S(N9904), .A(N9923), .B(N8971), .CI(N9111));
ADDFX1 inst_cellmath__203_0_I3362 (.CO(N9294), .S(N8919), .A(N10059), .B(N10199), .CI(N10089));
ADDFX1 inst_cellmath__203_0_I3363 (.CO(N10050), .S(N9687), .A(N8895), .B(N9877), .CI(N9134));
ADDFX1 inst_cellmath__203_0_I3364 (.CO(N9072), .S(N8731), .A(N9659), .B(N9904), .CI(N8919));
ADDFX1 inst_cellmath__203_0_I3365 (.CO(N9843), .S(N9456), .A(N8710), .B(N9687), .CI(N8731));
ADDFX1 inst_cellmath__203_0_I3366 (.CO(N8858), .S(N10201), .A(N9456), .B(N9428), .CI(N10170));
ADDFX1 inst_cellmath__203_0_I3367 (.CO(N9620), .S(N9229), .A(N10201), .B(N8659), .CI(N9201));
ADDFX1 inst_cellmath__203_0_I3368 (.CO(N8678), .S(N9990), .A(N10102), .B(N9927), .CI(N10273));
ADDFX1 inst_cellmath__203_0_I3369 (.CO(N9391), .S(N9012), .A(N9967), .B(N9229), .CI(N8981));
ADDFX1 inst_cellmath__203_0_I3370 (.CO(inst_cellmath__203__W0[30]), .S(inst_cellmath__203__W1[29]), .A(N9753), .B(N9990), .CI(N9012));
INVXL inst_cellmath__203_0_I3371 (.Y(N9433), .A(N9698));
ADDFX1 inst_cellmath__203_0_I3372 (.CO(N9162), .S(N8801), .A(N10276), .B(N9347), .CI(N9433));
ADDFX1 inst_cellmath__203_0_I3373 (.CO(N8945), .S(N10286), .A(N8859), .B(N9503), .CI(N8738));
ADDFX1 inst_cellmath__203_0_I3374 (.CO(N9716), .S(N9326), .A(N9526), .B(N9660), .CI(N10263));
ADDFX1 inst_cellmath__203_0_I3375 (.CO(N8748), .S(N10079), .A(N10286), .B(N8801), .CI(N9294));
ADDFX1 inst_cellmath__203_0_I3376 (.CO(N9486), .S(N9098), .A(N9326), .B(N10050), .CI(N10079));
ADDFX1 inst_cellmath__203_0_I3377 (.CO(N10229), .S(N9869), .A(N9098), .B(N9072), .CI(N9843));
ADDFX1 inst_cellmath__203_0_I3378 (.CO(N9257), .S(N8887), .A(N8858), .B(N9869), .CI(N9639));
ADDFX1 inst_cellmath__203_0_I3379 (.CO(N10017), .S(N9650), .A(N8887), .B(N9363), .CI(N8768));
ADDFX1 inst_cellmath__203_0_I3380 (.CO(N9037), .S(N8699), .A(N8933), .B(N9620), .CI(N9650));
ADDFX1 inst_cellmath__203_0_I3381 (.CO(inst_cellmath__203__W1[31]), .S(inst_cellmath__203__W1[30]), .A(N9391), .B(N8678), .CI(N8699));
ADDFX1 inst_cellmath__203_0_I3382 (.CO(N8828), .S(N10165), .A(N9740), .B(N9698), .CI(N9230));
ADDFX1 inst_cellmath__203_0_I3383 (.CO(N9582), .S(N9191), .A(N9885), .B(N8936), .CI(N9075));
ADDFX1 inst_cellmath__203_0_I3384 (.CO(N8648), .S(N9960), .A(N9162), .B(N10027), .CI(N8945));
ADDFX1 inst_cellmath__203_0_I3385 (.CO(N9354), .S(N8977), .A(N9191), .B(N10165), .CI(N9716));
ADDFX1 inst_cellmath__203_0_I3386 (.CO(N10109), .S(N9746), .A(N8748), .B(N9960), .CI(N8977));
ADDFX1 inst_cellmath__203_0_I3387 (.CO(N9127), .S(N8776), .A(N9746), .B(N9486), .CI(N10229));
ADDFX1 inst_cellmath__203_0_I3388 (.CO(N9896), .S(N9518), .A(N10118), .B(N8776), .CI(N9257));
ADDFX1 inst_cellmath__203_0_I3389 (.CO(N8915), .S(N10256), .A(N9309), .B(N9118), .CI(N9518));
ADDFX1 inst_cellmath__203_0_I3390 (.CO(inst_cellmath__203__W1[32]), .S(inst_cellmath__203__W0[31]), .A(N10256), .B(N10017), .CI(N9037));
INVXL inst_cellmath__203_0_I3391 (.Y(N9365), .A(N9857));
ADDFX1 inst_cellmath__203_0_I3392 (.CO(N8726), .S(N10045), .A(N10244), .B(N9313), .CI(N9365));
ADDFX1 inst_cellmath__203_0_I3393 (.CO(N10194), .S(N9835), .A(N8708), .B(N9463), .CI(N9618));
ADDFX1 inst_cellmath__203_0_I3394 (.CO(N9221), .S(N8852), .A(N9582), .B(N8828), .CI(N10045));
ADDFX1 inst_cellmath__203_0_I3395 (.CO(N9983), .S(N9611), .A(N8648), .B(N9835), .CI(N9354));
ADDFX1 inst_cellmath__203_0_I3396 (.CO(N9004), .S(N8671), .A(N9611), .B(N8852), .CI(N10109));
ADDFX1 inst_cellmath__203_0_I3397 (.CO(N9771), .S(N9382), .A(N9127), .B(N8671), .CI(N9137));
ADDFX1 inst_cellmath__203_0_I3398 (.CO(N8796), .S(N10132), .A(N9382), .B(N9795), .CI(N9896));
ADDFX1 inst_cellmath__203_0_I3399 (.CO(inst_cellmath__203__W1[33]), .S(inst_cellmath__203__W0[32]), .A(N10132), .B(N9699), .CI(N8915));
ADDFX1 inst_cellmath__203_0_I3400 (.CO(N10280), .S(N9926), .A(N9702), .B(N9857), .CI(N8904));
ADDFX1 inst_cellmath__203_0_I3401 (.CO(N9318), .S(N8940), .A(N9044), .B(N9853), .CI(N9991));
ADDFX1 inst_cellmath__203_0_I3402 (.CO(N10073), .S(N9709), .A(N10194), .B(N8726), .CI(N9926));
ADDFX1 inst_cellmath__203_0_I3403 (.CO(N9089), .S(N8744), .A(N9221), .B(N8940), .CI(N9709));
ADDFX1 inst_cellmath__203_0_I3404 (.CO(N9862), .S(N9478), .A(N8744), .B(N9983), .CI(N9004));
ADDFX1 inst_cellmath__203_0_I3405 (.CO(N8880), .S(N10221), .A(N9909), .B(N9478), .CI(N9771));
ADDFX1 inst_cellmath__203_0_I3406 (.CO(inst_cellmath__203__W1[34]), .S(inst_cellmath__203__W0[33]), .A(N10221), .B(N10067), .CI(N8796));
INVXL inst_cellmath__203_0_I3407 (.Y(N9299), .A(N10003));
ADDFX1 inst_cellmath__203_0_I3408 (.CO(N8694), .S(N10011), .A(N10206), .B(N9271), .CI(N9299));
ADDFX1 inst_cellmath__203_0_I3409 (.CO(N10159), .S(N9796), .A(N8679), .B(N9429), .CI(N10280));
ADDFX1 inst_cellmath__203_0_I3410 (.CO(N9181), .S(N8821), .A(N10011), .B(N9318), .CI(N9796));
ADDFX1 inst_cellmath__203_0_I3411 (.CO(N9954), .S(N9574), .A(N8821), .B(N10073), .CI(N9089));
ADDFX1 inst_cellmath__203_0_I3412 (.CO(N8967), .S(N10303), .A(N9862), .B(N9574), .CI(N8925));
ADDFX1 inst_cellmath__203_0_I3413 (.CO(inst_cellmath__203__W1[35]), .S(inst_cellmath__203__W0[34]), .A(N10303), .B(N9952), .CI(N8880));
ADDFX1 inst_cellmath__203_0_I3414 (.CO(N8769), .S(N10103), .A(N9667), .B(N10003), .CI(N8867));
ADDFX1 inst_cellmath__203_0_I3415 (.CO(N9509), .S(N9116), .A(N9010), .B(N9814), .CI(N8694));
ADDFX1 inst_cellmath__203_0_I3416 (.CO(N10249), .S(N9890), .A(N10159), .B(N10103), .CI(N9116));
ADDFX1 inst_cellmath__203_0_I3417 (.CO(N9279), .S(N8909), .A(N9890), .B(N9181), .CI(N9954));
ADDFX1 inst_cellmath__203_0_I3418 (.CO(inst_cellmath__203__W1[36]), .S(inst_cellmath__203__W0[35]), .A(N9692), .B(N8909), .CI(N8967));
INVXL inst_cellmath__203_0_I3419 (.Y(N9235), .A(N10148));
ADDFX1 inst_cellmath__203_0_I3420 (.CO(N9056), .S(N8718), .A(N10171), .B(N9238), .CI(N9235));
ADDFX1 inst_cellmath__203_0_I3421 (.CO(N8844), .S(N10185), .A(N8769), .B(N9392), .CI(N8718));
ADDFX1 inst_cellmath__203_0_I3422 (.CO(N9601), .S(N9212), .A(N10185), .B(N9509), .CI(N10249));
ADDFX1 inst_cellmath__203_0_I3423 (.CO(inst_cellmath__203__W1[37]), .S(inst_cellmath__203__W0[36]), .A(N9279), .B(N9212), .CI(N10192));
ADDFX1 inst_cellmath__203_0_I3424 (.CO(N9373), .S(N8994), .A(N9627), .B(N10148), .CI(N8836));
ADDFX1 inst_cellmath__203_0_I3425 (.CO(N10126), .S(N9763), .A(N9056), .B(N9779), .CI(N8994));
ADDFX1 inst_cellmath__203_0_I3426 (.CO(inst_cellmath__203__W1[38]), .S(inst_cellmath__203__W0[37]), .A(N9763), .B(N8844), .CI(N9601));
ADDFX1 inst_cellmath__203_0_I3427 (.CO(N9919), .S(N9538), .A(N9200), .B(N10298), .CI(N10137));
ADDFX1 inst_cellmath__203_0_I3428 (.CO(inst_cellmath__203__W1[39]), .S(inst_cellmath__203__W0[38]), .A(N9538), .B(N9373), .CI(N10126));
INVXL inst_cellmath__203_0_I3429 (.Y(N9307), .A(N9700));
ADDFX1 inst_cellmath__203_0_I3430 (.CO(inst_cellmath__203__W1[40]), .S(inst_cellmath__203__W0[39]), .A(N8802), .B(N9307), .CI(N9919));
ADDFX1 inst_cellmath__203_0_I3431 (.CO(inst_cellmath__203__W1[41]), .S(inst_cellmath__203__W0[40]), .A(N9700), .B(N8759), .CI(N9163));
INVXL inst_cellmath__203_0_I3432 (.Y(inst_cellmath__203__W0[41]), .A(inst_cellmath__203__W1[42]));
ADDHX1 cynw_cm_float_sin_I3435 (.CO(N12120), .S(N11989), .A(inst_cellmath__195[0]), .B(inst_cellmath__203__W0[18]));
ADDFX1 cynw_cm_float_sin_I3436 (.CO(N12405), .S(N12259), .A(inst_cellmath__203__W0[19]), .B(inst_cellmath__195[1]), .CI(inst_cellmath__203__W1[19]));
ADDFX1 cynw_cm_float_sin_I3437 (.CO(N12044), .S(N11906), .A(inst_cellmath__203__W0[20]), .B(inst_cellmath__195[2]), .CI(inst_cellmath__203__W1[20]));
ADDFX1 cynw_cm_float_sin_I3438 (.CO(N12317), .S(N12178), .A(inst_cellmath__203__W0[21]), .B(inst_cellmath__195[3]), .CI(inst_cellmath__203__W1[21]));
ADDFX1 cynw_cm_float_sin_I3439 (.CO(N11966), .S(N12458), .A(inst_cellmath__203__W0[22]), .B(inst_cellmath__195[4]), .CI(inst_cellmath__203__W1[22]));
ADDFX1 cynw_cm_float_sin_I3440 (.CO(N12235), .S(N12094), .A(inst_cellmath__203__W0[23]), .B(inst_cellmath__195[5]), .CI(inst_cellmath__203__W1[23]));
ADDFX1 cynw_cm_float_sin_I3441 (.CO(N12512), .S(N12381), .A(inst_cellmath__203__W0[24]), .B(inst_cellmath__195[6]), .CI(inst_cellmath__203__W1[24]));
ADDFX1 cynw_cm_float_sin_I3442 (.CO(N12155), .S(N12022), .A(inst_cellmath__203__W0[25]), .B(inst_cellmath__195[7]), .CI(inst_cellmath__203__W1[25]));
ADDFX1 cynw_cm_float_sin_I3443 (.CO(N12436), .S(N12294), .A(inst_cellmath__203__W0[26]), .B(inst_cellmath__195[8]), .CI(inst_cellmath__203__W1[26]));
ADDFX1 cynw_cm_float_sin_I3444 (.CO(N12072), .S(N11942), .A(inst_cellmath__203__W0[27]), .B(inst_cellmath__195[9]), .CI(inst_cellmath__203__W1[27]));
ADDFX1 cynw_cm_float_sin_I3445 (.CO(N12354), .S(N12212), .A(inst_cellmath__203__W0[28]), .B(inst_cellmath__195[10]), .CI(inst_cellmath__203__W1[28]));
ADDFX1 cynw_cm_float_sin_I3446 (.CO(N12000), .S(N12491), .A(inst_cellmath__203__W0[29]), .B(inst_cellmath__195[11]), .CI(inst_cellmath__203__W1[29]));
ADDFX1 cynw_cm_float_sin_I3447 (.CO(N12272), .S(N12132), .A(inst_cellmath__203__W0[30]), .B(inst_cellmath__195[12]), .CI(inst_cellmath__203__W1[30]));
ADDFX1 cynw_cm_float_sin_I3448 (.CO(N11919), .S(N12416), .A(inst_cellmath__203__W0[31]), .B(inst_cellmath__195[13]), .CI(inst_cellmath__203__W1[31]));
ADDFX1 cynw_cm_float_sin_I3449 (.CO(N12189), .S(N12054), .A(inst_cellmath__203__W0[32]), .B(inst_cellmath__195[14]), .CI(inst_cellmath__203__W1[32]));
ADDFX1 cynw_cm_float_sin_I3450 (.CO(N12469), .S(N12329), .A(inst_cellmath__203__W0[33]), .B(inst_cellmath__195[15]), .CI(inst_cellmath__203__W1[33]));
ADDFX1 cynw_cm_float_sin_I3451 (.CO(N12108), .S(N11977), .A(inst_cellmath__203__W0[34]), .B(inst_cellmath__195[16]), .CI(inst_cellmath__203__W1[34]));
ADDFX1 cynw_cm_float_sin_I3452 (.CO(N12392), .S(N12245), .A(inst_cellmath__203__W1[35]), .B(inst_cellmath__195[17]), .CI(inst_cellmath__203__W0[35]));
ADDFX1 cynw_cm_float_sin_I3453 (.CO(N12033), .S(N12522), .A(inst_cellmath__203__W0[36]), .B(inst_cellmath__195[18]), .CI(inst_cellmath__203__W1[36]));
ADDFX1 cynw_cm_float_sin_I3454 (.CO(N12305), .S(N12164), .A(inst_cellmath__203__W0[37]), .B(inst_cellmath__195[19]), .CI(inst_cellmath__203__W1[37]));
ADDFX1 cynw_cm_float_sin_I3455 (.CO(N11951), .S(N12446), .A(inst_cellmath__203__W0[38]), .B(inst_cellmath__195[20]), .CI(inst_cellmath__203__W1[38]));
ADDFX1 cynw_cm_float_sin_I3456 (.CO(N12222), .S(N12080), .A(inst_cellmath__203__W0[39]), .B(inst_cellmath__195[21]), .CI(inst_cellmath__203__W1[39]));
ADDFX1 cynw_cm_float_sin_I3457 (.CO(N12501), .S(N12365), .A(inst_cellmath__203__W0[40]), .B(inst_cellmath__195[22]), .CI(inst_cellmath__203__W1[40]));
ADDFX1 cynw_cm_float_sin_I3458 (.CO(N12140), .S(N12008), .A(inst_cellmath__203__W0[41]), .B(inst_cellmath__195[23]), .CI(inst_cellmath__203__W1[41]));
ADDFX1 cynw_cm_float_sin_I3459 (.CO(N12424), .S(N12283), .A(inst_cellmath__203__W1[42]), .B(inst_cellmath__203__W0[42]), .CI(inst_cellmath__195[24]));
ADDHX1 cynw_cm_float_sin_I3460 (.CO(N12059), .S(N11929), .A(1'B1), .B(inst_cellmath__195[25]));
ADDHX1 cynw_cm_float_sin_I3461 (.CO(N12337), .S(N12197), .A(1'B1), .B(inst_cellmath__195[26]));
ADDHX1 cynw_cm_float_sin_I3462 (.CO(N11984), .S(N12476), .A(1'B1), .B(inst_cellmath__195[27]));
INVXL hap1_A_I23833 (.Y(N12117), .A(inst_cellmath__195[28]));
OR2XL hap1_A_I8522 (.Y(N12255), .A(1'B0), .B(inst_cellmath__195[28]));
NOR3BXL cynw_cm_float_sin_I8507 (.Y(N12400), .AN(N6248), .B(N6355), .C(N6521));
AND2XL cynw_cm_float_sin_I3469 (.Y(N12230), .A(inst_cellmath__203__W0[2]), .B(inst_cellmath__203__W1[2]));
NOR2XL cynw_cm_float_sin_I3470 (.Y(N12376), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
NAND2XL cynw_cm_float_sin_I3471 (.Y(N12509), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
AND2XL cynw_cm_float_sin_I3473 (.Y(N12151), .A(inst_cellmath__203__W0[4]), .B(inst_cellmath__203__W1[4]));
NOR2XL cynw_cm_float_sin_I3474 (.Y(N12291), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
NAND2XL cynw_cm_float_sin_I3475 (.Y(N12432), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
AND2XL cynw_cm_float_sin_I3477 (.Y(N12069), .A(inst_cellmath__203__W0[6]), .B(inst_cellmath__203__W1[6]));
NOR2XL cynw_cm_float_sin_I3478 (.Y(N12207), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
NAND2XL cynw_cm_float_sin_I3479 (.Y(N12350), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
AND2XL cynw_cm_float_sin_I3481 (.Y(N11996), .A(inst_cellmath__203__W0[8]), .B(inst_cellmath__203__W1[8]));
NOR2XL cynw_cm_float_sin_I3482 (.Y(N12128), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
NAND2XL cynw_cm_float_sin_I3483 (.Y(N12270), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
AND2XL cynw_cm_float_sin_I3485 (.Y(N11915), .A(inst_cellmath__203__W0[10]), .B(inst_cellmath__203__W1[10]));
NOR2XL cynw_cm_float_sin_I3486 (.Y(N12052), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
NAND2XL cynw_cm_float_sin_I3487 (.Y(N12185), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
AND2XL cynw_cm_float_sin_I3489 (.Y(N12467), .A(inst_cellmath__203__W0[12]), .B(inst_cellmath__203__W1[12]));
NOR2XL cynw_cm_float_sin_I3490 (.Y(N11973), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NAND2XL cynw_cm_float_sin_I3491 (.Y(N12104), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NOR2XL cynw_cm_float_sin_I3492 (.Y(N12243), .A(inst_cellmath__203__W0[14]), .B(inst_cellmath__203__W1[14]));
NOR2XL cynw_cm_float_sin_I3494 (.Y(N12519), .A(inst_cellmath__203__W0[15]), .B(inst_cellmath__203__W1[15]));
NAND2XL cynw_cm_float_sin_I3495 (.Y(N12031), .A(inst_cellmath__203__W0[15]), .B(inst_cellmath__203__W1[15]));
NOR2XL cynw_cm_float_sin_I3496 (.Y(N12161), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
NOR2XL cynw_cm_float_sin_I3498 (.Y(N12444), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
NAND2XL cynw_cm_float_sin_I3499 (.Y(N11948), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
AND2XL cynw_cm_float_sin_I3501 (.Y(N12220), .A(inst_cellmath__203__W1[18]), .B(N11989));
AND2XL cynw_cm_float_sin_I3503 (.Y(N12498), .A(N12120), .B(N12259));
AND2XL cynw_cm_float_sin_I23834 (.Y(N12278), .A(inst_cellmath__203__W0[1]), .B(inst_cellmath__203__W1[1]));
OAI22XL cynw_cm_float_sin_I8470 (.Y(N12112), .A0(N12230), .A1(N12278), .B0(inst_cellmath__203__W0[2]), .B1(inst_cellmath__203__W1[2]));
AOI21XL cynw_cm_float_sin_I3508 (.Y(N11958), .A0(N12509), .A1(N12112), .B0(N12376));
OAI22XL cynw_cm_float_sin_I8471 (.Y(N12346), .A0(N12151), .A1(N11958), .B0(inst_cellmath__203__W0[4]), .B1(inst_cellmath__203__W1[4]));
AOI21XL cynw_cm_float_sin_I3512 (.Y(N12101), .A0(N12432), .A1(N12346), .B0(N12291));
OAI22XL cynw_cm_float_sin_I8472 (.Y(N12421), .A0(N12069), .A1(N12101), .B0(inst_cellmath__203__W0[6]), .B1(inst_cellmath__203__W1[6]));
AOI21XL cynw_cm_float_sin_I3516 (.Y(N12083), .A0(N12350), .A1(N12421), .B0(N12207));
OAI22XL cynw_cm_float_sin_I8473 (.Y(N12320), .A0(N11996), .A1(N12083), .B0(inst_cellmath__203__W0[8]), .B1(inst_cellmath__203__W1[8]));
AOI21XL cynw_cm_float_sin_I3520 (.Y(N11920), .A0(N12270), .A1(N12320), .B0(N12128));
OAI22XL cynw_cm_float_sin_I8474 (.Y(N12061), .A0(N11915), .A1(N11920), .B0(inst_cellmath__203__W0[10]), .B1(inst_cellmath__203__W1[10]));
AOI21XL cynw_cm_float_sin_I3524 (.Y(N12210), .A0(N12185), .A1(N12061), .B0(N12052));
OAI22XL cynw_cm_float_sin_I8475 (.Y(N12281), .A0(N12467), .A1(N12210), .B0(inst_cellmath__203__W0[12]), .B1(inst_cellmath__203__W1[12]));
AOI21XL cynw_cm_float_sin_I3528 (.Y(N12348), .A0(N12104), .A1(N12281), .B0(N11973));
AOI21XL cynw_cm_float_sin_I3529 (.Y(N12266), .A0(N12031), .A1(N12243), .B0(N12519));
OAI2BB1X1 cynw_cm_float_sin_I8476 (.Y(N12410), .A0N(inst_cellmath__203__W0[14]), .A1N(inst_cellmath__203__W1[14]), .B0(N12031));
OAI21XL cynw_cm_float_sin_I3531 (.Y(N12250), .A0(N12410), .A1(N12348), .B0(N12266));
AOI21XL cynw_cm_float_sin_I3532 (.Y(N12169), .A0(N11948), .A1(N12161), .B0(N12444));
OAI2BB1X1 cynw_cm_float_sin_I8477 (.Y(N12310), .A0N(inst_cellmath__203__W0[16]), .A1N(inst_cellmath__203__W1[16]), .B0(N11948));
OAI22XL cynw_cm_float_sin_I8478 (.Y(N12014), .A0(N12220), .A1(N12169), .B0(inst_cellmath__203__W1[18]), .B1(N11989));
NOR2XL cynw_cm_float_sin_I3539 (.Y(N12148), .A(N12220), .B(N12310));
AOI21XL cynw_cm_float_sin_I3544 (.Y(N12192), .A0(N12148), .A1(N12250), .B0(N12014));
OAI22XL cynw_cm_float_sin_I8479 (.Y(N12360), .A0(N12498), .A1(N12192), .B0(N12120), .B1(N12259));
NOR2XL cynw_cm_float_sin_I3587 (.Y(N12007), .A(N12405), .B(N11906));
NAND2XL cynw_cm_float_sin_I3588 (.Y(N12137), .A(N12405), .B(N11906));
NOR2XL cynw_cm_float_sin_I3589 (.Y(N12279), .A(N12044), .B(N12178));
NAND2XL cynw_cm_float_sin_I3590 (.Y(N12423), .A(N12044), .B(N12178));
NOR2XL cynw_cm_float_sin_I3591 (.Y(N11925), .A(N12317), .B(N12458));
NAND2XL cynw_cm_float_sin_I3592 (.Y(N12057), .A(N12317), .B(N12458));
NOR2XL cynw_cm_float_sin_I3593 (.Y(N12196), .A(N11966), .B(N12094));
NAND2XL cynw_cm_float_sin_I3594 (.Y(N12333), .A(N11966), .B(N12094));
NOR2XL cynw_cm_float_sin_I3595 (.Y(N12473), .A(N12235), .B(N12381));
NAND2XL cynw_cm_float_sin_I3596 (.Y(N11983), .A(N12235), .B(N12381));
NOR2XL cynw_cm_float_sin_I3597 (.Y(N12113), .A(N12512), .B(N12022));
NAND2XL cynw_cm_float_sin_I3598 (.Y(N12252), .A(N12512), .B(N12022));
NOR2XL cynw_cm_float_sin_I3599 (.Y(N12399), .A(N12155), .B(N12294));
NAND2XL cynw_cm_float_sin_I3600 (.Y(N11899), .A(N12155), .B(N12294));
NOR2XL cynw_cm_float_sin_I3601 (.Y(N12037), .A(N12436), .B(N11942));
NAND2XL cynw_cm_float_sin_I3602 (.Y(N12172), .A(N12436), .B(N11942));
NOR2XL cynw_cm_float_sin_I3603 (.Y(N12311), .A(N12072), .B(N12212));
NAND2XL cynw_cm_float_sin_I3604 (.Y(N12451), .A(N12072), .B(N12212));
NOR2XL cynw_cm_float_sin_I3605 (.Y(N11959), .A(N12354), .B(N12491));
NAND2XL cynw_cm_float_sin_I3606 (.Y(N12087), .A(N12354), .B(N12491));
NOR2XL cynw_cm_float_sin_I3607 (.Y(N12227), .A(N12000), .B(N12132));
NAND2XL cynw_cm_float_sin_I3608 (.Y(N12374), .A(N12000), .B(N12132));
NOR2XL cynw_cm_float_sin_I3609 (.Y(N12506), .A(N12272), .B(N12416));
NAND2XL cynw_cm_float_sin_I3610 (.Y(N12015), .A(N12272), .B(N12416));
NOR2XL cynw_cm_float_sin_I3611 (.Y(N12149), .A(N11919), .B(N12054));
NAND2XL cynw_cm_float_sin_I3612 (.Y(N12288), .A(N11919), .B(N12054));
NOR2XL cynw_cm_float_sin_I3613 (.Y(N12429), .A(N12189), .B(N12329));
NAND2XL cynw_cm_float_sin_I3614 (.Y(N11936), .A(N12189), .B(N12329));
NOR2XL cynw_cm_float_sin_I3615 (.Y(N12066), .A(N12469), .B(N11977));
NAND2XL cynw_cm_float_sin_I3616 (.Y(N12204), .A(N12469), .B(N11977));
NOR2XL cynw_cm_float_sin_I3617 (.Y(N12347), .A(N12108), .B(N12245));
NAND2XL cynw_cm_float_sin_I3618 (.Y(N12485), .A(N12108), .B(N12245));
NOR2XL cynw_cm_float_sin_I3619 (.Y(N11993), .A(N12522), .B(N12392));
NAND2XL cynw_cm_float_sin_I3620 (.Y(N12126), .A(N12522), .B(N12392));
NOR2XL cynw_cm_float_sin_I3621 (.Y(N12265), .A(N12164), .B(N12033));
NAND2XL cynw_cm_float_sin_I3622 (.Y(N12408), .A(N12164), .B(N12033));
NOR2XL cynw_cm_float_sin_I3623 (.Y(N11912), .A(N12446), .B(N12305));
NAND2XL cynw_cm_float_sin_I3624 (.Y(N12048), .A(N12446), .B(N12305));
NOR2XL cynw_cm_float_sin_I3625 (.Y(N12182), .A(N12080), .B(N11951));
NAND2XL cynw_cm_float_sin_I3626 (.Y(N12323), .A(N12080), .B(N11951));
NOR2XL cynw_cm_float_sin_I3627 (.Y(N12464), .A(N12365), .B(N12222));
NAND2XL cynw_cm_float_sin_I3628 (.Y(N11970), .A(N12365), .B(N12222));
NOR2XL cynw_cm_float_sin_I3629 (.Y(N12102), .A(N12008), .B(N12501));
NAND2XL cynw_cm_float_sin_I3630 (.Y(N12240), .A(N12008), .B(N12501));
NOR2XL cynw_cm_float_sin_I3631 (.Y(N12385), .A(N12283), .B(N12140));
NAND2XL cynw_cm_float_sin_I3632 (.Y(N12517), .A(N12283), .B(N12140));
NOR2XL cynw_cm_float_sin_I3633 (.Y(N12028), .A(N12424), .B(N11929));
NAND2XL cynw_cm_float_sin_I3634 (.Y(N12158), .A(N12424), .B(N11929));
NOR2XL cynw_cm_float_sin_I3635 (.Y(N12300), .A(N12059), .B(N12197));
NAND2XL cynw_cm_float_sin_I3636 (.Y(N12441), .A(N12059), .B(N12197));
NOR2XL cynw_cm_float_sin_I3637 (.Y(N11946), .A(N12337), .B(N12476));
NAND2XL cynw_cm_float_sin_I3638 (.Y(N12077), .A(N12337), .B(N12476));
NOR2XL cynw_cm_float_sin_I3639 (.Y(N12218), .A(N11984), .B(N12117));
NAND2XL cynw_cm_float_sin_I3640 (.Y(N12357), .A(N11984), .B(N12117));
NOR2XL cynw_cm_float_sin_I3641 (.Y(N12497), .A(N12400), .B(N12255));
NAND2XL cynw_cm_float_sin_I3642 (.Y(N12005), .A(N12400), .B(N12255));
AO21XL cynw_cm_float_sin_I3643 (.Y(N11923), .A0(N12137), .A1(N12360), .B0(N12007));
AO21XL cynw_cm_float_sin_I3644 (.Y(N12194), .A0(N12423), .A1(N12007), .B0(N12279));
AND2XL cynw_cm_float_sin_I3645 (.Y(N12331), .A(N12423), .B(N12137));
AO21XL cynw_cm_float_sin_I3646 (.Y(N12472), .A0(N12057), .A1(N12279), .B0(N11925));
AND2XL cynw_cm_float_sin_I3647 (.Y(N11981), .A(N12057), .B(N12423));
AO21XL cynw_cm_float_sin_I3648 (.Y(N12110), .A0(N12333), .A1(N11925), .B0(N12196));
AND2XL cynw_cm_float_sin_I3649 (.Y(N12249), .A(N12333), .B(N12057));
AO21XL cynw_cm_float_sin_I3650 (.Y(N12397), .A0(N11983), .A1(N12196), .B0(N12473));
AND2XL cynw_cm_float_sin_I3651 (.Y(N12524), .A(N11983), .B(N12333));
AO21XL cynw_cm_float_sin_I3652 (.Y(N12036), .A0(N12252), .A1(N12473), .B0(N12113));
AND2XL cynw_cm_float_sin_I3653 (.Y(N12168), .A(N12252), .B(N11983));
AO21XL cynw_cm_float_sin_I3654 (.Y(N12308), .A0(N11899), .A1(N12113), .B0(N12399));
AND2XL cynw_cm_float_sin_I3655 (.Y(N12449), .A(N11899), .B(N12252));
AO21XL cynw_cm_float_sin_I3656 (.Y(N11956), .A0(N12172), .A1(N12399), .B0(N12037));
AND2XL cynw_cm_float_sin_I3657 (.Y(N12084), .A(N12172), .B(N11899));
AO21XL cynw_cm_float_sin_I3658 (.Y(N12226), .A0(N12451), .A1(N12037), .B0(N12311));
AND2XL cynw_cm_float_sin_I3659 (.Y(N12371), .A(N12451), .B(N12172));
AO21XL cynw_cm_float_sin_I3660 (.Y(N12504), .A0(N12087), .A1(N12311), .B0(N11959));
AND2XL cynw_cm_float_sin_I3661 (.Y(N12013), .A(N12087), .B(N12451));
AO21XL cynw_cm_float_sin_I3662 (.Y(N12146), .A0(N12374), .A1(N11959), .B0(N12227));
AND2XL cynw_cm_float_sin_I3663 (.Y(N12286), .A(N12374), .B(N12087));
AO21XL cynw_cm_float_sin_I3664 (.Y(N12427), .A0(N12015), .A1(N12227), .B0(N12506));
AND2XL cynw_cm_float_sin_I3665 (.Y(N11933), .A(N12015), .B(N12374));
AO21XL cynw_cm_float_sin_I3666 (.Y(N12063), .A0(N12288), .A1(N12506), .B0(N12149));
AND2XL cynw_cm_float_sin_I3667 (.Y(N12202), .A(N12288), .B(N12015));
AO21XL cynw_cm_float_sin_I3668 (.Y(N12344), .A0(N11936), .A1(N12149), .B0(N12429));
AND2XL cynw_cm_float_sin_I3669 (.Y(N12481), .A(N11936), .B(N12288));
AO21XL cynw_cm_float_sin_I3670 (.Y(N11991), .A0(N12204), .A1(N12429), .B0(N12066));
AND2XL cynw_cm_float_sin_I3671 (.Y(N12123), .A(N12204), .B(N11936));
AO21XL cynw_cm_float_sin_I3672 (.Y(N12261), .A0(N12485), .A1(N12066), .B0(N12347));
AND2XL cynw_cm_float_sin_I3673 (.Y(N12406), .A(N12485), .B(N12204));
AO21XL cynw_cm_float_sin_I3674 (.Y(N11910), .A0(N12126), .A1(N12347), .B0(N11993));
AND2XL cynw_cm_float_sin_I3675 (.Y(N12045), .A(N12126), .B(N12485));
AO21XL cynw_cm_float_sin_I3676 (.Y(N12180), .A0(N12408), .A1(N11993), .B0(N12265));
AND2XL cynw_cm_float_sin_I3677 (.Y(N12321), .A(N12408), .B(N12126));
AO21XL cynw_cm_float_sin_I3678 (.Y(N12460), .A0(N12048), .A1(N12265), .B0(N11912));
AND2XL cynw_cm_float_sin_I3679 (.Y(N11968), .A(N12048), .B(N12408));
AO21XL cynw_cm_float_sin_I3680 (.Y(N12099), .A0(N12323), .A1(N11912), .B0(N12182));
AND2XL cynw_cm_float_sin_I3681 (.Y(N12236), .A(N12323), .B(N12048));
AO21XL cynw_cm_float_sin_I3682 (.Y(N12383), .A0(N11970), .A1(N12182), .B0(N12464));
AND2XL cynw_cm_float_sin_I3683 (.Y(N12515), .A(N11970), .B(N12323));
AO21XL cynw_cm_float_sin_I3684 (.Y(N12024), .A0(N12240), .A1(N12464), .B0(N12102));
AND2XL cynw_cm_float_sin_I3685 (.Y(N12156), .A(N12240), .B(N11970));
AO21XL cynw_cm_float_sin_I3686 (.Y(N12298), .A0(N12517), .A1(N12102), .B0(N12385));
AND2XL cynw_cm_float_sin_I3687 (.Y(N12437), .A(N12517), .B(N12240));
AO21XL cynw_cm_float_sin_I3688 (.Y(N11944), .A0(N12158), .A1(N12385), .B0(N12028));
AND2XL cynw_cm_float_sin_I3689 (.Y(N12075), .A(N12158), .B(N12517));
AO21XL cynw_cm_float_sin_I3690 (.Y(N12214), .A0(N12441), .A1(N12028), .B0(N12300));
AND2XL cynw_cm_float_sin_I3691 (.Y(N12355), .A(N12441), .B(N12158));
AO21XL cynw_cm_float_sin_I3692 (.Y(N12495), .A0(N12077), .A1(N12300), .B0(N11946));
AND2XL cynw_cm_float_sin_I3693 (.Y(N12002), .A(N12077), .B(N12441));
AO21XL cynw_cm_float_sin_I3694 (.Y(N12135), .A0(N12357), .A1(N11946), .B0(N12218));
AND2XL cynw_cm_float_sin_I3695 (.Y(N12276), .A(N12357), .B(N12077));
AO21XL cynw_cm_float_sin_I3696 (.Y(N12418), .A0(N12005), .A1(N12218), .B0(N12497));
AND2XL cynw_cm_float_sin_I3697 (.Y(N11921), .A(N12005), .B(N12357));
AND2XL cynw_cm_float_sin_I3698 (.Y(N12330), .A(N12400), .B(N12005));
AO21XL cynw_cm_float_sin_I3699 (.Y(N12394), .A0(N12331), .A1(N12360), .B0(N12194));
AO21XL cynw_cm_float_sin_I3700 (.Y(N12035), .A0(N11981), .A1(N11923), .B0(N12472));
AO21XL cynw_cm_float_sin_I3701 (.Y(N12307), .A0(N12249), .A1(N12194), .B0(N12110));
AND2XL cynw_cm_float_sin_I3702 (.Y(N12448), .A(N12249), .B(N12331));
AO21XL cynw_cm_float_sin_I3703 (.Y(N11953), .A0(N12524), .A1(N12472), .B0(N12397));
AND2XL cynw_cm_float_sin_I3704 (.Y(N12082), .A(N12524), .B(N11981));
AO21XL cynw_cm_float_sin_I3705 (.Y(N12225), .A0(N12168), .A1(N12110), .B0(N12036));
AND2XL cynw_cm_float_sin_I3706 (.Y(N12367), .A(N12168), .B(N12249));
AO21XL cynw_cm_float_sin_I3707 (.Y(N12503), .A0(N12449), .A1(N12397), .B0(N12308));
AND2XL cynw_cm_float_sin_I3708 (.Y(N12011), .A(N12449), .B(N12524));
AO21XL cynw_cm_float_sin_I3709 (.Y(N12143), .A0(N12084), .A1(N12036), .B0(N11956));
AND2XL cynw_cm_float_sin_I3710 (.Y(N12285), .A(N12084), .B(N12168));
AO21XL cynw_cm_float_sin_I3711 (.Y(N12426), .A0(N12371), .A1(N12308), .B0(N12226));
AND2XL cynw_cm_float_sin_I3712 (.Y(N11931), .A(N12371), .B(N12449));
AO21XL cynw_cm_float_sin_I3713 (.Y(N12062), .A0(N12013), .A1(N11956), .B0(N12504));
AND2XL cynw_cm_float_sin_I3714 (.Y(N12201), .A(N12013), .B(N12084));
AO21XL cynw_cm_float_sin_I3715 (.Y(N12341), .A0(N12286), .A1(N12226), .B0(N12146));
AND2XL cynw_cm_float_sin_I3716 (.Y(N12479), .A(N12286), .B(N12371));
AO21XL cynw_cm_float_sin_I3717 (.Y(N11988), .A0(N11933), .A1(N12504), .B0(N12427));
AND2XL cynw_cm_float_sin_I3718 (.Y(N12121), .A(N11933), .B(N12013));
AO21XL cynw_cm_float_sin_I3719 (.Y(N12258), .A0(N12202), .A1(N12146), .B0(N12063));
AND2XL cynw_cm_float_sin_I3720 (.Y(N12404), .A(N12202), .B(N12286));
AO21XL cynw_cm_float_sin_I3721 (.Y(N11907), .A0(N12481), .A1(N12427), .B0(N12344));
AND2XL cynw_cm_float_sin_I3722 (.Y(N12043), .A(N12481), .B(N11933));
AO21XL cynw_cm_float_sin_I3723 (.Y(N12177), .A0(N12123), .A1(N12063), .B0(N11991));
AND2XL cynw_cm_float_sin_I3724 (.Y(N12318), .A(N12123), .B(N12202));
AO21XL cynw_cm_float_sin_I3725 (.Y(N12457), .A0(N12406), .A1(N12344), .B0(N12261));
AND2XL cynw_cm_float_sin_I3726 (.Y(N11965), .A(N12406), .B(N12481));
AO21XL cynw_cm_float_sin_I3727 (.Y(N12095), .A0(N12045), .A1(N11991), .B0(N11910));
AND2XL cynw_cm_float_sin_I3728 (.Y(N12234), .A(N12045), .B(N12123));
AO21XL cynw_cm_float_sin_I3729 (.Y(N12380), .A0(N12321), .A1(N12261), .B0(N12180));
AND2XL cynw_cm_float_sin_I3730 (.Y(N12513), .A(N12321), .B(N12406));
AO21XL cynw_cm_float_sin_I3731 (.Y(N12021), .A0(N11968), .A1(N11910), .B0(N12460));
AND2XL cynw_cm_float_sin_I3732 (.Y(N12154), .A(N11968), .B(N12045));
AO21XL cynw_cm_float_sin_I3733 (.Y(N12295), .A0(N12236), .A1(N12180), .B0(N12099));
AND2XL cynw_cm_float_sin_I3734 (.Y(N12435), .A(N12236), .B(N12321));
AO21XL cynw_cm_float_sin_I3735 (.Y(N11941), .A0(N12515), .A1(N12460), .B0(N12383));
AND2XL cynw_cm_float_sin_I3736 (.Y(N12073), .A(N12515), .B(N11968));
AO21XL cynw_cm_float_sin_I3737 (.Y(N12211), .A0(N12156), .A1(N12099), .B0(N12024));
AND2XL cynw_cm_float_sin_I3738 (.Y(N12353), .A(N12156), .B(N12236));
AO21XL cynw_cm_float_sin_I3739 (.Y(N12492), .A0(N12437), .A1(N12383), .B0(N12298));
AND2XL cynw_cm_float_sin_I3740 (.Y(N11999), .A(N12437), .B(N12515));
AO21XL cynw_cm_float_sin_I3741 (.Y(N12131), .A0(N12075), .A1(N12024), .B0(N11944));
AND2XL cynw_cm_float_sin_I3742 (.Y(N12273), .A(N12075), .B(N12156));
AO21XL cynw_cm_float_sin_I3743 (.Y(N12415), .A0(N12355), .A1(N12298), .B0(N12214));
AND2XL cynw_cm_float_sin_I3744 (.Y(N11918), .A(N12355), .B(N12437));
AO21XL cynw_cm_float_sin_I3745 (.Y(N12055), .A0(N12002), .A1(N11944), .B0(N12495));
AND2XL cynw_cm_float_sin_I3746 (.Y(N12188), .A(N12002), .B(N12075));
AO21XL cynw_cm_float_sin_I3747 (.Y(N12328), .A0(N12276), .A1(N12214), .B0(N12135));
AND2XL cynw_cm_float_sin_I3748 (.Y(N12470), .A(N12276), .B(N12355));
AO21XL cynw_cm_float_sin_I3749 (.Y(N11976), .A0(N11921), .A1(N12495), .B0(N12418));
AND2XL cynw_cm_float_sin_I3750 (.Y(N12107), .A(N11921), .B(N12002));
AO22XL cynw_cm_float_sin_I3751 (.Y(N12246), .A0(N12400), .A1(N12497), .B0(N12330), .B1(N12135));
AND2XL cynw_cm_float_sin_I3752 (.Y(N12391), .A(N12330), .B(N12276));
AO21XL cynw_cm_float_sin_I3753 (.Y(N12364), .A0(N12448), .A1(N12360), .B0(N12307));
AO21XL cynw_cm_float_sin_I3754 (.Y(N12009), .A0(N12082), .A1(N11923), .B0(N11953));
AO21XL cynw_cm_float_sin_I3755 (.Y(N12282), .A0(N12367), .A1(N12394), .B0(N12225));
AO21XL cynw_cm_float_sin_I3756 (.Y(N11928), .A0(N12011), .A1(N12035), .B0(N12503));
AO21XL cynw_cm_float_sin_I3757 (.Y(N12198), .A0(N12285), .A1(N12307), .B0(N12143));
AND2XL cynw_cm_float_sin_I3758 (.Y(N12336), .A(N12285), .B(N12448));
AO21XL cynw_cm_float_sin_I3759 (.Y(N12475), .A0(N11931), .A1(N11953), .B0(N12426));
AND2XL cynw_cm_float_sin_I3760 (.Y(N11985), .A(N11931), .B(N12082));
AO21XL cynw_cm_float_sin_I3761 (.Y(N12116), .A0(N12201), .A1(N12225), .B0(N12062));
AND2XL cynw_cm_float_sin_I3762 (.Y(N12254), .A(N12201), .B(N12367));
AO21XL cynw_cm_float_sin_I3763 (.Y(N12401), .A0(N12479), .A1(N12503), .B0(N12341));
AND2XL cynw_cm_float_sin_I3764 (.Y(N11902), .A(N12479), .B(N12011));
AO21XL cynw_cm_float_sin_I3765 (.Y(N12040), .A0(N12121), .A1(N12143), .B0(N11988));
AND2XL cynw_cm_float_sin_I3766 (.Y(N12174), .A(N12121), .B(N12285));
AO21XL cynw_cm_float_sin_I3767 (.Y(N12313), .A0(N12404), .A1(N12426), .B0(N12258));
AND2XL cynw_cm_float_sin_I3768 (.Y(N12453), .A(N12404), .B(N11931));
AO21XL cynw_cm_float_sin_I3769 (.Y(N11961), .A0(N12043), .A1(N12062), .B0(N11907));
AND2XL cynw_cm_float_sin_I3770 (.Y(N12090), .A(N12043), .B(N12201));
AO21XL cynw_cm_float_sin_I3771 (.Y(N12229), .A0(N12318), .A1(N12341), .B0(N12177));
AND2XL cynw_cm_float_sin_I3772 (.Y(N12375), .A(N12318), .B(N12479));
AO21XL cynw_cm_float_sin_I3773 (.Y(N12508), .A0(N11965), .A1(N11988), .B0(N12457));
AND2XL cynw_cm_float_sin_I3774 (.Y(N12017), .A(N11965), .B(N12121));
AO21XL cynw_cm_float_sin_I3775 (.Y(N12150), .A0(N12234), .A1(N12258), .B0(N12095));
AND2XL cynw_cm_float_sin_I3776 (.Y(N12290), .A(N12234), .B(N12404));
AO21XL cynw_cm_float_sin_I3777 (.Y(N12431), .A0(N12513), .A1(N11907), .B0(N12380));
AND2XL cynw_cm_float_sin_I3778 (.Y(N11937), .A(N12513), .B(N12043));
AO21XL cynw_cm_float_sin_I3779 (.Y(N12068), .A0(N12154), .A1(N12177), .B0(N12021));
AND2XL cynw_cm_float_sin_I3780 (.Y(N12206), .A(N12154), .B(N12318));
AO21XL cynw_cm_float_sin_I3781 (.Y(N12349), .A0(N12435), .A1(N12457), .B0(N12295));
AND2XL cynw_cm_float_sin_I3782 (.Y(N12487), .A(N12435), .B(N11965));
AO21XL cynw_cm_float_sin_I3783 (.Y(N11995), .A0(N12073), .A1(N12095), .B0(N11941));
AND2XL cynw_cm_float_sin_I3784 (.Y(N12127), .A(N12073), .B(N12234));
AO21XL cynw_cm_float_sin_I3785 (.Y(N12269), .A0(N12353), .A1(N12380), .B0(N12211));
AND2XL cynw_cm_float_sin_I3786 (.Y(N12411), .A(N12353), .B(N12513));
AO21XL cynw_cm_float_sin_I3787 (.Y(N11914), .A0(N11999), .A1(N12021), .B0(N12492));
AND2XL cynw_cm_float_sin_I3788 (.Y(N12051), .A(N11999), .B(N12154));
AO21XL cynw_cm_float_sin_I3789 (.Y(N12184), .A0(N12273), .A1(N12295), .B0(N12131));
AND2XL cynw_cm_float_sin_I3790 (.Y(N12324), .A(N12273), .B(N12435));
AO21XL cynw_cm_float_sin_I3791 (.Y(N12466), .A0(N11918), .A1(N11941), .B0(N12415));
AND2XL cynw_cm_float_sin_I3792 (.Y(N11972), .A(N11918), .B(N12073));
AO21XL cynw_cm_float_sin_I3793 (.Y(N12103), .A0(N12188), .A1(N12211), .B0(N12055));
AND2XL cynw_cm_float_sin_I3794 (.Y(N12242), .A(N12188), .B(N12353));
AO21XL cynw_cm_float_sin_I3795 (.Y(N12387), .A0(N12470), .A1(N12492), .B0(N12328));
AND2XL cynw_cm_float_sin_I3796 (.Y(N12518), .A(N12470), .B(N11999));
AO21XL cynw_cm_float_sin_I3797 (.Y(N12030), .A0(N12107), .A1(N12131), .B0(N11976));
AND2XL cynw_cm_float_sin_I3798 (.Y(N12160), .A(N12107), .B(N12273));
AO21XL cynw_cm_float_sin_I3799 (.Y(N12302), .A0(N12391), .A1(N12415), .B0(N12246));
AND2XL cynw_cm_float_sin_I3800 (.Y(N12443), .A(N12391), .B(N11918));
AO21XL cynw_cm_float_sin_I3801 (.Y(N12251), .A0(N12336), .A1(N12360), .B0(N12198));
AO21XL cynw_cm_float_sin_I3802 (.Y(N11898), .A0(N11985), .A1(N11923), .B0(N12475));
AO21XL cynw_cm_float_sin_I3803 (.Y(N12171), .A0(N12254), .A1(N12394), .B0(N12116));
AO21XL cynw_cm_float_sin_I3804 (.Y(N12450), .A0(N11902), .A1(N12035), .B0(N12401));
AO21XL cynw_cm_float_sin_I3805 (.Y(N12086), .A0(N12174), .A1(N12364), .B0(N12040));
AO21XL cynw_cm_float_sin_I3806 (.Y(N12373), .A0(N12453), .A1(N12009), .B0(N12313));
AO21XL cynw_cm_float_sin_I3807 (.Y(N11935), .A0(N12017), .A1(N12198), .B0(N12508));
AND2XL cynw_cm_float_sin_I3808 (.Y(N12065), .A(N12017), .B(N12336));
AO21XL cynw_cm_float_sin_I3809 (.Y(N12203), .A0(N12290), .A1(N12475), .B0(N12150));
AND2XL cynw_cm_float_sin_I3810 (.Y(N12345), .A(N12290), .B(N11985));
AO21XL cynw_cm_float_sin_I3811 (.Y(N12484), .A0(N11937), .A1(N12116), .B0(N12431));
AND2XL cynw_cm_float_sin_I3812 (.Y(N11992), .A(N11937), .B(N12254));
AO21XL cynw_cm_float_sin_I3813 (.Y(N12125), .A0(N12206), .A1(N12401), .B0(N12068));
AND2XL cynw_cm_float_sin_I3814 (.Y(N12263), .A(N12206), .B(N11902));
AO21XL cynw_cm_float_sin_I3815 (.Y(N12407), .A0(N12487), .A1(N12040), .B0(N12349));
AND2XL cynw_cm_float_sin_I3816 (.Y(N11911), .A(N12487), .B(N12174));
AO21XL cynw_cm_float_sin_I3817 (.Y(N12047), .A0(N12127), .A1(N12313), .B0(N11995));
AND2XL cynw_cm_float_sin_I3818 (.Y(N12181), .A(N12127), .B(N12453));
AO21XL cynw_cm_float_sin_I3819 (.Y(N12322), .A0(N12411), .A1(N11961), .B0(N12269));
AND2XL cynw_cm_float_sin_I3820 (.Y(N12463), .A(N12411), .B(N12090));
AO21XL cynw_cm_float_sin_I3821 (.Y(N11969), .A0(N12051), .A1(N12229), .B0(N11914));
AND2XL cynw_cm_float_sin_I3822 (.Y(N12100), .A(N12051), .B(N12375));
AO21XL cynw_cm_float_sin_I3823 (.Y(N12239), .A0(N12324), .A1(N12508), .B0(N12184));
AND2XL cynw_cm_float_sin_I3824 (.Y(N12384), .A(N12324), .B(N12017));
AO21XL cynw_cm_float_sin_I3825 (.Y(N12516), .A0(N11972), .A1(N12150), .B0(N12466));
AND2XL cynw_cm_float_sin_I3826 (.Y(N12027), .A(N11972), .B(N12290));
AO21XL cynw_cm_float_sin_I3827 (.Y(N12157), .A0(N12242), .A1(N12431), .B0(N12103));
AND2XL cynw_cm_float_sin_I3828 (.Y(N12299), .A(N12242), .B(N11937));
AO21XL cynw_cm_float_sin_I3829 (.Y(N12440), .A0(N12518), .A1(N12068), .B0(N12387));
AND2XL cynw_cm_float_sin_I3830 (.Y(N11945), .A(N12518), .B(N12206));
AO21XL cynw_cm_float_sin_I3831 (.Y(N12076), .A0(N12160), .A1(N12349), .B0(N12030));
AND2XL cynw_cm_float_sin_I3832 (.Y(N12217), .A(N12160), .B(N12487));
AO21XL cynw_cm_float_sin_I3833 (.Y(N12356), .A0(N12443), .A1(N11995), .B0(N12302));
AOI21XL cynw_cm_float_sin_I3835 (.Y(N12124), .A0(N12090), .A1(N12282), .B0(N11961));
AOI21XL cynw_cm_float_sin_I3836 (.Y(N12264), .A0(N12375), .A1(N11928), .B0(N12229));
AO21XL cynw_cm_float_sin_I3837 (.Y(N11990), .A0(N12065), .A1(N12360), .B0(N11935));
AO21XL cynw_cm_float_sin_I3838 (.Y(N12260), .A0(N12345), .A1(N11923), .B0(N12203));
AO21XL cynw_cm_float_sin_I3839 (.Y(N11909), .A0(N11992), .A1(N12394), .B0(N12484));
AO21XL cynw_cm_float_sin_I3840 (.Y(N12179), .A0(N12263), .A1(N12035), .B0(N12125));
AO21XL cynw_cm_float_sin_I3841 (.Y(N12459), .A0(N11911), .A1(N12364), .B0(N12407));
AO21XL cynw_cm_float_sin_I3842 (.Y(N12097), .A0(N12181), .A1(N12009), .B0(N12047));
AO21XL cynw_cm_float_sin_I3843 (.Y(N12382), .A0(N12463), .A1(N12282), .B0(N12322));
AO21XL cynw_cm_float_sin_I3844 (.Y(N12023), .A0(N12100), .A1(N11928), .B0(N11969));
AO21XL cynw_cm_float_sin_I3845 (.Y(N12297), .A0(N12384), .A1(N12251), .B0(N12239));
AO21XL cynw_cm_float_sin_I3846 (.Y(N11943), .A0(N12027), .A1(N11898), .B0(N12516));
AO21XL cynw_cm_float_sin_I3847 (.Y(N12213), .A0(N12299), .A1(N12171), .B0(N12157));
AO21XL cynw_cm_float_sin_I3848 (.Y(N12494), .A0(N11945), .A1(N12450), .B0(N12440));
AO21XL cynw_cm_float_sin_I3849 (.Y(N12133), .A0(N12217), .A1(N12086), .B0(N12076));
NAND2BXL cynw_cm_float_sin_I3856 (.Y(N12284), .AN(N12113), .B(N12252));
NAND2BXL cynw_cm_float_sin_I3857 (.Y(N12060), .AN(N12399), .B(N11899));
NAND2BXL cynw_cm_float_sin_I3858 (.Y(N12478), .AN(N12037), .B(N12172));
NAND2BXL cynw_cm_float_sin_I3859 (.Y(N12257), .AN(N12311), .B(N12451));
NAND2BXL cynw_cm_float_sin_I3860 (.Y(N12042), .AN(N11959), .B(N12087));
NAND2BXL cynw_cm_float_sin_I3861 (.Y(N12456), .AN(N12227), .B(N12374));
NAND2BXL cynw_cm_float_sin_I3862 (.Y(N12232), .AN(N12506), .B(N12015));
NAND2BXL cynw_cm_float_sin_I3863 (.Y(N12020), .AN(N12149), .B(N12288));
NAND2BXL cynw_cm_float_sin_I3864 (.Y(N12434), .AN(N12429), .B(N11936));
NAND2BXL cynw_cm_float_sin_I3865 (.Y(N12209), .AN(N12066), .B(N12204));
NAND2BXL cynw_cm_float_sin_I3866 (.Y(N11998), .AN(N12347), .B(N12485));
NAND2BXL cynw_cm_float_sin_I3867 (.Y(N12414), .AN(N11993), .B(N12126));
NAND2BXL cynw_cm_float_sin_I3868 (.Y(N12187), .AN(N12265), .B(N12408));
NAND2BXL cynw_cm_float_sin_I3869 (.Y(N11975), .AN(N11912), .B(N12048));
NAND2BXL cynw_cm_float_sin_I3870 (.Y(N12390), .AN(N12182), .B(N12323));
NAND2BXL cynw_cm_float_sin_I3871 (.Y(N12163), .AN(N12464), .B(N11970));
NAND2BXL cynw_cm_float_sin_I3872 (.Y(N11950), .AN(N12102), .B(N12240));
NAND2BXL cynw_cm_float_sin_I3873 (.Y(N12362), .AN(N12385), .B(N12517));
NAND2BXL cynw_cm_float_sin_I3874 (.Y(N12138), .AN(N12028), .B(N12158));
NAND2BXL cynw_cm_float_sin_I3875 (.Y(N11927), .AN(N12300), .B(N12441));
NAND2BXL cynw_cm_float_sin_I3876 (.Y(N12335), .AN(N11946), .B(N12077));
NAND2BXL cynw_cm_float_sin_I3877 (.Y(N12115), .AN(N12218), .B(N12357));
NAND2BXL cynw_cm_float_sin_I3878 (.Y(N11901), .AN(N12497), .B(N12005));
XOR2XL cynw_cm_float_sin_I3884 (.Y(inst_cellmath__201[25]), .A(N12009), .B(N12284));
XOR2XL cynw_cm_float_sin_I3885 (.Y(inst_cellmath__201[26]), .A(N12282), .B(N12060));
XOR2XL cynw_cm_float_sin_I3886 (.Y(inst_cellmath__201[27]), .A(N11928), .B(N12478));
XOR2XL cynw_cm_float_sin_I3887 (.Y(inst_cellmath__201[28]), .A(N12251), .B(N12257));
XOR2XL cynw_cm_float_sin_I3888 (.Y(inst_cellmath__201[29]), .A(N11898), .B(N12042));
XOR2XL cynw_cm_float_sin_I3889 (.Y(inst_cellmath__201[30]), .A(N12171), .B(N12456));
XOR2XL cynw_cm_float_sin_I3890 (.Y(inst_cellmath__201[31]), .A(N12450), .B(N12232));
XOR2XL cynw_cm_float_sin_I3891 (.Y(inst_cellmath__201[32]), .A(N12086), .B(N12020));
XOR2XL cynw_cm_float_sin_I3892 (.Y(inst_cellmath__201[33]), .A(N12373), .B(N12434));
XNOR2X1 cynw_cm_float_sin_I3893 (.Y(inst_cellmath__201[34]), .A(N12124), .B(N12209));
XNOR2X1 cynw_cm_float_sin_I3894 (.Y(inst_cellmath__201[35]), .A(N12264), .B(N11998));
XOR2XL cynw_cm_float_sin_I3895 (.Y(inst_cellmath__201[36]), .A(N11990), .B(N12414));
XOR2XL cynw_cm_float_sin_I3896 (.Y(inst_cellmath__201[37]), .A(N12260), .B(N12187));
XOR2XL cynw_cm_float_sin_I3897 (.Y(inst_cellmath__201[38]), .A(N11909), .B(N11975));
XOR2XL cynw_cm_float_sin_I3898 (.Y(inst_cellmath__201[39]), .A(N12179), .B(N12390));
XOR2XL cynw_cm_float_sin_I3899 (.Y(inst_cellmath__201[40]), .A(N12459), .B(N12163));
XOR2XL cynw_cm_float_sin_I3900 (.Y(inst_cellmath__201[41]), .A(N12097), .B(N11950));
XOR2XL cynw_cm_float_sin_I3901 (.Y(inst_cellmath__201[42]), .A(N12382), .B(N12362));
XOR2XL cynw_cm_float_sin_I3902 (.Y(inst_cellmath__201[43]), .A(N12023), .B(N12138));
XOR2XL cynw_cm_float_sin_I3903 (.Y(inst_cellmath__201[44]), .A(N12297), .B(N11927));
XOR2XL cynw_cm_float_sin_I3904 (.Y(inst_cellmath__201[45]), .A(N11943), .B(N12335));
XOR2XL cynw_cm_float_sin_I3905 (.Y(inst_cellmath__201[46]), .A(N12213), .B(N12115));
XOR2XL cynw_cm_float_sin_I3906 (.Y(inst_cellmath__201[47]), .A(N12494), .B(N11901));
XNOR2X1 cynw_cm_float_sin_I3907 (.Y(inst_cellmath__201[48]), .A(N12133), .B(N12400));
AOI31X1 inst_cellmath__200_0_I8508 (.Y(N13041), .A0(N12443), .A1(N12127), .A2(N12373), .B0(N12356));
AND2XL inst_cellmath__200_0_I3934 (.Y(inst_cellmath__210[0]), .A(N13041), .B(inst_cellmath__201[25]));
AND2XL inst_cellmath__200_0_I3935 (.Y(inst_cellmath__210[1]), .A(N13041), .B(inst_cellmath__201[26]));
AND2XL inst_cellmath__200_0_I3936 (.Y(inst_cellmath__210[2]), .A(N13041), .B(inst_cellmath__201[27]));
AND2XL inst_cellmath__200_0_I3937 (.Y(inst_cellmath__210[3]), .A(N13041), .B(inst_cellmath__201[28]));
AND2XL inst_cellmath__200_0_I3938 (.Y(inst_cellmath__210[4]), .A(N13041), .B(inst_cellmath__201[29]));
AND2XL inst_cellmath__200_0_I3939 (.Y(inst_cellmath__210[5]), .A(N13041), .B(inst_cellmath__201[30]));
AND2XL inst_cellmath__200_0_I3940 (.Y(inst_cellmath__210[6]), .A(N13041), .B(inst_cellmath__201[31]));
AND2XL inst_cellmath__200_0_I3941 (.Y(inst_cellmath__210[7]), .A(N13041), .B(inst_cellmath__201[32]));
AND2XL inst_cellmath__200_0_I3942 (.Y(inst_cellmath__210[8]), .A(N13041), .B(inst_cellmath__201[33]));
AND2XL inst_cellmath__200_0_I3943 (.Y(inst_cellmath__210[9]), .A(N13041), .B(inst_cellmath__201[34]));
AND2XL inst_cellmath__200_0_I3944 (.Y(inst_cellmath__210[10]), .A(N13041), .B(inst_cellmath__201[35]));
AND2XL inst_cellmath__200_0_I3945 (.Y(inst_cellmath__210[11]), .A(N13041), .B(inst_cellmath__201[36]));
AND2XL inst_cellmath__200_0_I3946 (.Y(inst_cellmath__210[12]), .A(N13041), .B(inst_cellmath__201[37]));
AND2XL inst_cellmath__200_0_I3947 (.Y(inst_cellmath__210[13]), .A(N13041), .B(inst_cellmath__201[38]));
AND2XL inst_cellmath__200_0_I3948 (.Y(inst_cellmath__210[14]), .A(N13041), .B(inst_cellmath__201[39]));
AND2XL inst_cellmath__200_0_I3949 (.Y(inst_cellmath__210[15]), .A(N13041), .B(inst_cellmath__201[40]));
AND2XL inst_cellmath__200_0_I3950 (.Y(inst_cellmath__210[16]), .A(N13041), .B(inst_cellmath__201[41]));
AND2XL inst_cellmath__200_0_I3951 (.Y(inst_cellmath__210[17]), .A(N13041), .B(inst_cellmath__201[42]));
AND2XL inst_cellmath__200_0_I3952 (.Y(inst_cellmath__210[18]), .A(N13041), .B(inst_cellmath__201[43]));
AND2XL inst_cellmath__200_0_I3953 (.Y(inst_cellmath__210[19]), .A(N13041), .B(inst_cellmath__201[44]));
AND2XL inst_cellmath__200_0_I3954 (.Y(inst_cellmath__210[20]), .A(N13041), .B(inst_cellmath__201[45]));
AND2XL inst_cellmath__200_0_I3955 (.Y(inst_cellmath__210[21]), .A(N13041), .B(inst_cellmath__201[46]));
AND2XL inst_cellmath__200_0_I3956 (.Y(inst_cellmath__210[22]), .A(N13041), .B(inst_cellmath__201[47]));
NAND2XL inst_cellmath__19_0_I3958 (.Y(N13185), .A(a_exp[7]), .B(a_exp[0]));
AND4XL inst_cellmath__19_0_I23835 (.Y(N13187), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL hyperpropagate_4_1_A_I8523 (.Y(N19047), .A(a_exp[6]), .B(a_exp[5]), .C(N13187));
NOR2XL hyperpropagate_4_1_A_I8524 (.Y(inst_cellmath__19), .A(N13185), .B(N19047));
NOR2XL inst_cellmath__24_0_I3971 (.Y(N13208), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__24_0_I3972 (.Y(N13216), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__24_0_I3973 (.Y(N13227), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__24_0_I3974 (.Y(N13236), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__24_0_I23836 (.Y(N13221), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__24_0_I23837 (.Y(N13230), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__24_0_I23838 (.Y(N13240), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__24_0_I3978 (.Y(N13225), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N13221));
NAND4XL inst_cellmath__24_0_I3980 (.Y(N13219), .A(N13208), .B(N13227), .C(N13216), .D(N13236));
NOR4BX1 inst_cellmath__24_0_I23839 (.Y(inst_cellmath__24), .AN(N13225), .B(N13219), .C(N13230), .D(N13240));
AND2XL cynw_cm_float_sin_I23840 (.Y(inst_cellmath__68), .A(inst_cellmath__19), .B(inst_cellmath__24));
INVXL buf1_A_I8525 (.Y(N19054), .A(inst_cellmath__19));
INVXL buf1_A_I8526 (.Y(inst_cellmath__82), .A(N19054));
OR4X1 inst_cellmath__17_0_I23841 (.Y(N13288), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 inst_cellmath__17_0_I23842 (.Y(N13292), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NOR2XL inst_cellmath__17_0_I3995 (.Y(inst_cellmath__17), .A(N13288), .B(N13292));
OR2XL cynw_cm_float_sin_I3996 (.Y(N487), .A(inst_cellmath__17), .B(inst_cellmath__68));
OR3XL cynw_cm_float_sin_I3997 (.Y(N759), .A(inst_cellmath__82), .B(inst_cellmath__68), .C(N487));
AND4XL inst_cellmath__216__184__I3998 (.Y(N13316), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[5]), .D(a_exp[6]));
NOR2X1 inst_cellmath__216__184__I3999 (.Y(N639), .A(a_exp[7]), .B(N13316));
AND3XL cynw_cm_float_sin_I8483 (.Y(inst_cellmath__219), .A(N13041), .B(inst_cellmath__61[22]), .C(inst_cellmath__201[48]));
INVXL inst_cellmath__211__182__I4001 (.Y(N13398), .A(inst_cellmath__210[22]));
INVXL inst_cellmath__211__182__I4002 (.Y(N13340), .A(inst_cellmath__210[0]));
INVXL inst_cellmath__211__182__I4003 (.Y(N13376), .A(inst_cellmath__210[2]));
OAI21XL inst_cellmath__211__182__I4004 (.Y(N13393), .A0(inst_cellmath__210[1]), .A1(N13340), .B0(N13376));
OR2XL inst_cellmath__211__182__I4005 (.Y(N13397), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[1]));
NOR2BX1 inst_cellmath__211__182__I4006 (.Y(N13384), .AN(inst_cellmath__210[3]), .B(inst_cellmath__210[4]));
INVXL inst_cellmath__211__182__I4007 (.Y(N13402), .A(inst_cellmath__210[6]));
OAI21XL inst_cellmath__211__182__I4008 (.Y(N13337), .A0(inst_cellmath__210[5]), .A1(N13384), .B0(N13402));
NOR2XL inst_cellmath__211__182__I4009 (.Y(N13355), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[3]));
NOR2XL inst_cellmath__211__182__I4010 (.Y(N13371), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[5]));
NOR2BX1 inst_cellmath__211__182__I4011 (.Y(N13409), .AN(inst_cellmath__210[7]), .B(inst_cellmath__210[8]));
INVXL inst_cellmath__211__182__I4012 (.Y(N13343), .A(inst_cellmath__210[10]));
OAI21XL inst_cellmath__211__182__I4013 (.Y(N13362), .A0(inst_cellmath__210[9]), .A1(N13409), .B0(N13343));
NOR2XL inst_cellmath__211__182__I4014 (.Y(N13380), .A(inst_cellmath__210[8]), .B(inst_cellmath__210[7]));
NOR2XL inst_cellmath__211__182__I4015 (.Y(N13399), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[9]));
NOR2BX1 inst_cellmath__211__182__I4016 (.Y(N13352), .AN(inst_cellmath__210[11]), .B(inst_cellmath__210[12]));
INVXL inst_cellmath__211__182__I4017 (.Y(N13368), .A(inst_cellmath__210[14]));
OAI21XL inst_cellmath__211__182__I4018 (.Y(N13388), .A0(inst_cellmath__210[13]), .A1(N13352), .B0(N13368));
NOR2XL inst_cellmath__211__182__I4019 (.Y(N13407), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[11]));
NOR2XL inst_cellmath__211__182__I4020 (.Y(N13341), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[13]));
NOR2BX1 inst_cellmath__211__182__I4021 (.Y(N13377), .AN(inst_cellmath__210[15]), .B(inst_cellmath__210[16]));
INVXL inst_cellmath__211__182__I4022 (.Y(N13395), .A(inst_cellmath__210[18]));
OAI21XL inst_cellmath__211__182__I4023 (.Y(N13332), .A0(inst_cellmath__210[17]), .A1(N13377), .B0(N13395));
NOR2XL inst_cellmath__211__182__I4024 (.Y(N13348), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[15]));
NOR2XL inst_cellmath__211__182__I4025 (.Y(N13365), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[17]));
NOR2BX1 inst_cellmath__211__182__I4026 (.Y(N13404), .AN(inst_cellmath__210[19]), .B(inst_cellmath__210[20]));
OAI21XL inst_cellmath__211__182__I4027 (.Y(N13358), .A0(inst_cellmath__210[21]), .A1(N13404), .B0(N13398));
NOR2XL inst_cellmath__211__182__I4028 (.Y(N13373), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[19]));
NOR2XL inst_cellmath__211__182__I4029 (.Y(N13391), .A(inst_cellmath__210[22]), .B(inst_cellmath__210[21]));
INVXL inst_cellmath__211__182__I4030 (.Y(N13349), .A(N13371));
AOI21XL inst_cellmath__211__182__I4031 (.Y(N13367), .A0(N13355), .A1(N13397), .B0(N13349));
NAND2XL inst_cellmath__211__182__I4032 (.Y(N13405), .A(N13371), .B(N13355));
NAND2BXL inst_cellmath__211__182__I4033 (.Y(N13359), .AN(N13380), .B(N13399));
INVXL inst_cellmath__211__182__I4034 (.Y(N13375), .A(N13341));
AOI21XL inst_cellmath__211__182__I4035 (.Y(N13392), .A0(N13407), .A1(N13359), .B0(N13375));
NAND2XL inst_cellmath__211__182__I4036 (.Y(N13411), .A(N13399), .B(N13380));
NAND2XL inst_cellmath__211__182__I4037 (.Y(N13346), .A(N13341), .B(N13407));
NAND2BXL inst_cellmath__211__182__I4038 (.Y(N13383), .AN(N13348), .B(N13365));
NAND2XL inst_cellmath__211__182__I4039 (.Y(N13354), .A(N13365), .B(N13348));
NAND2XL inst_cellmath__211__182__I4040 (.Y(N13370), .A(N13391), .B(N13373));
INVXL inst_cellmath__211__182__I4041 (.Y(N13351), .A(N13405));
INVXL inst_cellmath__211__182__I4042 (.Y(N13387), .A(N13346));
OAI21XL inst_cellmath__211__182__I4043 (.Y(N13406), .A0(N13411), .A1(N13351), .B0(N13387));
NOR2XL inst_cellmath__211__182__I4044 (.Y(N13356), .A(N13346), .B(N13411));
NAND2BXL inst_cellmath__211__182__I4045 (.Y(N13347), .AN(N13370), .B(N13354));
OR2XL inst_cellmath__211__182__I4046 (.Y(N13386), .A(N13370), .B(N13354));
OR2XL inst_cellmath__211__182__I4047 (.Y(N544), .A(N13386), .B(N13356));
OAI21XL inst_cellmath__211__182__I4049 (.Y(N543), .A0(N13386), .A1(N13406), .B0(N13347));
AOI21XL inst_cellmath__211__182__I4050 (.Y(N13339), .A0(N13356), .A1(N13367), .B0(N13392));
OAI2BB1X1 inst_cellmath__211__182__I4051 (.Y(N13374), .A0N(N13373), .A1N(N13383), .B0(N13391));
OAI21XL inst_cellmath__211__182__I4052 (.Y(N542), .A0(N13386), .A1(N13339), .B0(N13374));
OAI21XL inst_cellmath__211__182__I4053 (.Y(N13379), .A0(N13405), .A1(N13393), .B0(N13337));
OAI21XL inst_cellmath__211__182__I4054 (.Y(N13334), .A0(N13346), .A1(N13362), .B0(N13388));
AOI21XL inst_cellmath__211__182__I4055 (.Y(N13360), .A0(N13356), .A1(N13379), .B0(N13334));
OA21X1 inst_cellmath__211__182__I4056 (.Y(N13394), .A0(N13332), .A1(N13370), .B0(N13358));
OAI21XL inst_cellmath__211__182__I4057 (.Y(N541), .A0(N13386), .A1(N13360), .B0(N13394));
INVXL inst_cellmath__215_0_I4058 (.Y(inst_cellmath__215[0]), .A(N541));
NAND2XL inst_cellmath__215_0_I4059 (.Y(N13472), .A(N542), .B(N541));
NAND3XL inst_cellmath__215_0_I4060 (.Y(N13470), .A(N543), .B(N542), .C(N541));
NAND2BXL inst_cellmath__215_0_I4061 (.Y(N13475), .AN(N544), .B(N13470));
XOR2XL inst_cellmath__215_0_I4064 (.Y(inst_cellmath__215[3]), .A(N13470), .B(N544));
INVXL inst_cellmath__220__188__I4066 (.Y(N13601), .A(inst_cellmath__215[0]));
AND2XL inst_cellmath__220__188__I4067 (.Y(N13639), .A(N13601), .B(inst_cellmath__210[0]));
MX2XL inst_cellmath__220__188__I4068 (.Y(N13555), .A(inst_cellmath__210[0]), .B(inst_cellmath__210[1]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4069 (.Y(N13589), .A(inst_cellmath__210[1]), .B(inst_cellmath__210[2]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4070 (.Y(N13623), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[3]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4071 (.Y(N13503), .A(inst_cellmath__210[3]), .B(inst_cellmath__210[4]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4072 (.Y(N13534), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[5]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4073 (.Y(N13571), .A(inst_cellmath__210[5]), .B(inst_cellmath__210[6]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4074 (.Y(N13604), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[7]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4075 (.Y(N13635), .A(inst_cellmath__210[7]), .B(inst_cellmath__210[8]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4076 (.Y(N13518), .A(inst_cellmath__210[8]), .B(inst_cellmath__210[9]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4077 (.Y(N13548), .A(inst_cellmath__210[9]), .B(inst_cellmath__210[10]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4078 (.Y(N13583), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[11]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4079 (.Y(N13617), .A(inst_cellmath__210[11]), .B(inst_cellmath__210[12]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4080 (.Y(N13497), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[13]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4081 (.Y(N13527), .A(inst_cellmath__210[13]), .B(inst_cellmath__210[14]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4082 (.Y(N13565), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[15]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4083 (.Y(N13598), .A(inst_cellmath__210[15]), .B(inst_cellmath__210[16]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4084 (.Y(N13629), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[17]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4085 (.Y(N13512), .A(inst_cellmath__210[17]), .B(inst_cellmath__210[18]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4086 (.Y(N13541), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[19]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4087 (.Y(N13577), .A(inst_cellmath__210[19]), .B(inst_cellmath__210[20]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4088 (.Y(N13612), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[21]), .S0(N13601));
MX2XL inst_cellmath__220__188__I4089 (.Y(N13492), .A(inst_cellmath__210[21]), .B(inst_cellmath__210[22]), .S0(N13601));
XOR2XL inst_cellmath__220__188__I8484 (.Y(N13594), .A(inst_cellmath__215[0]), .B(N542));
INVXL inst_cellmath__220__188__I4091 (.Y(N13609), .A(N13594));
NAND2XL inst_cellmath__220__188__I4092 (.Y(N13507), .A(N13639), .B(N13594));
NAND2XL inst_cellmath__220__188__I4093 (.Y(N13574), .A(N13555), .B(N13594));
AOI22XL inst_cellmath__220__188__I4094 (.Y(N13638), .A0(N13609), .A1(N13639), .B0(N13589), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4095 (.Y(N13521), .A0(N13609), .A1(N13555), .B0(N13623), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4096 (.Y(N13554), .A0(N13609), .A1(N13589), .B0(N13503), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4097 (.Y(N13587), .A0(N13609), .A1(N13623), .B0(N13534), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4098 (.Y(N13621), .A0(N13609), .A1(N13503), .B0(N13571), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4099 (.Y(N13502), .A0(N13609), .A1(N13534), .B0(N13604), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4100 (.Y(N13533), .A0(N13609), .A1(N13571), .B0(N13635), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4101 (.Y(N13570), .A0(N13609), .A1(N13604), .B0(N13518), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4102 (.Y(N13603), .A0(N13609), .A1(N13635), .B0(N13548), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4103 (.Y(N13634), .A0(N13609), .A1(N13518), .B0(N13583), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4104 (.Y(N13517), .A0(N13609), .A1(N13548), .B0(N13617), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4105 (.Y(N13547), .A0(N13609), .A1(N13583), .B0(N13497), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4106 (.Y(N13582), .A0(N13609), .A1(N13617), .B0(N13527), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4107 (.Y(N13616), .A0(N13609), .A1(N13497), .B0(N13565), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4108 (.Y(N13496), .A0(N13609), .A1(N13527), .B0(N13598), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4109 (.Y(N13526), .A0(N13609), .A1(N13565), .B0(N13629), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4110 (.Y(N13563), .A0(N13609), .A1(N13598), .B0(N13512), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4111 (.Y(N13596), .A0(N13609), .A1(N13629), .B0(N13541), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4112 (.Y(N13628), .A0(N13609), .A1(N13512), .B0(N13577), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4113 (.Y(N13511), .A0(N13609), .A1(N13541), .B0(N13612), .B1(N13594));
AOI22XL inst_cellmath__220__188__I4114 (.Y(N13540), .A0(N13609), .A1(N13577), .B0(N13492), .B1(N13594));
XOR2XL inst_cellmath__220__188__I8485 (.Y(N13549), .A(N13472), .B(N543));
INVXL inst_cellmath__220__188__I4116 (.Y(N13566), .A(N13549));
NOR2XL inst_cellmath__220__188__I4117 (.Y(N13560), .A(N13566), .B(N13507));
NOR2XL inst_cellmath__220__188__I4118 (.Y(N13506), .A(N13566), .B(N13574));
NOR2XL inst_cellmath__220__188__I4119 (.Y(N13608), .A(N13566), .B(N13638));
NOR2XL inst_cellmath__220__188__I4120 (.Y(N13553), .A(N13566), .B(N13521));
AOI22XL inst_cellmath__220__188__I4121 (.Y(N13501), .A0(N13549), .A1(N13554), .B0(N13507), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4122 (.Y(N13532), .A0(N13549), .A1(N13587), .B0(N13574), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4123 (.Y(N13569), .A0(N13549), .A1(N13621), .B0(N13638), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4124 (.Y(N13602), .A0(N13549), .A1(N13502), .B0(N13521), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4125 (.Y(N13633), .A0(N13549), .A1(N13533), .B0(N13554), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4126 (.Y(N13516), .A0(N13549), .A1(N13570), .B0(N13587), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4127 (.Y(N13546), .A0(N13549), .A1(N13603), .B0(N13621), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4128 (.Y(N13581), .A0(N13549), .A1(N13634), .B0(N13502), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4129 (.Y(N13615), .A0(N13549), .A1(N13517), .B0(N13533), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4130 (.Y(N13495), .A0(N13549), .A1(N13547), .B0(N13570), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4131 (.Y(N13525), .A0(N13549), .A1(N13582), .B0(N13603), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4132 (.Y(N13562), .A0(N13549), .A1(N13616), .B0(N13634), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4133 (.Y(N13595), .A0(N13549), .A1(N13496), .B0(N13517), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4134 (.Y(N13627), .A0(N13549), .A1(N13526), .B0(N13547), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4135 (.Y(N13510), .A0(N13549), .A1(N13563), .B0(N13582), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4136 (.Y(N13539), .A0(N13549), .A1(N13596), .B0(N13616), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4137 (.Y(N13576), .A0(N13549), .A1(N13628), .B0(N13496), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4138 (.Y(N13610), .A0(N13549), .A1(N13511), .B0(N13526), .B1(N13566));
AOI22XL inst_cellmath__220__188__I4139 (.Y(N13490), .A0(N13549), .A1(N13540), .B0(N13563), .B1(N13566));
INVXL inst_cellmath__220__188__I4140 (.Y(N13551), .A(inst_cellmath__215[3]));
NAND2XL inst_cellmath__220__188__I4141 (.Y(N13509), .A(N13560), .B(N13551));
NAND2XL inst_cellmath__220__188__I4142 (.Y(N13575), .A(N13506), .B(N13551));
NAND2XL inst_cellmath__220__188__I4143 (.Y(N13640), .A(N13608), .B(N13551));
NAND2XL inst_cellmath__220__188__I4144 (.Y(N13556), .A(N13553), .B(N13551));
NAND2XL inst_cellmath__220__188__I4145 (.Y(N13622), .A(N13501), .B(N13551));
NAND2XL inst_cellmath__220__188__I4146 (.Y(N13535), .A(N13532), .B(N13551));
NAND2XL inst_cellmath__220__188__I4147 (.Y(N13605), .A(N13569), .B(N13551));
AOI22XL inst_cellmath__220__188__I4148 (.Y(N13584), .A0(inst_cellmath__215[3]), .A1(N13560), .B0(N13633), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4149 (.Y(N13618), .A0(inst_cellmath__215[3]), .A1(N13506), .B0(N13516), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4150 (.Y(N13498), .A0(inst_cellmath__215[3]), .A1(N13608), .B0(N13546), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4151 (.Y(N13528), .A0(inst_cellmath__215[3]), .A1(N13553), .B0(N13581), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4152 (.Y(N13564), .A0(inst_cellmath__215[3]), .A1(N13501), .B0(N13615), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4153 (.Y(N13597), .A0(inst_cellmath__215[3]), .A1(N13532), .B0(N13495), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4154 (.Y(N13630), .A0(inst_cellmath__215[3]), .A1(N13569), .B0(N13525), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4155 (.Y(N13513), .A0(inst_cellmath__215[3]), .A1(N13602), .B0(N13562), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4156 (.Y(N13542), .A0(inst_cellmath__215[3]), .A1(N13633), .B0(N13595), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4157 (.Y(N13578), .A0(inst_cellmath__215[3]), .A1(N13516), .B0(N13627), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4158 (.Y(N13611), .A0(inst_cellmath__215[3]), .A1(N13546), .B0(N13510), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4159 (.Y(N13491), .A0(inst_cellmath__215[3]), .A1(N13581), .B0(N13539), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4160 (.Y(N13522), .A0(inst_cellmath__215[3]), .A1(N13615), .B0(N13576), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4161 (.Y(N13558), .A0(inst_cellmath__215[3]), .A1(N13495), .B0(N13610), .B1(N13551));
AOI22XL inst_cellmath__220__188__I4162 (.Y(N13591), .A0(inst_cellmath__215[3]), .A1(N13525), .B0(N13490), .B1(N13551));
XNOR2X1 inst_cellmath__220__188__I8486 (.Y(N13531), .A(N13475), .B(N13386));
INVXL inst_cellmath__220__188__I4164 (.Y(N13545), .A(N13531));
NOR2XL inst_cellmath__220__188__I4165 (.Y(N679), .A(N13545), .B(N13509));
NOR2XL inst_cellmath__220__188__I4166 (.Y(N680), .A(N13545), .B(N13575));
NOR2XL inst_cellmath__220__188__I4167 (.Y(N681), .A(N13545), .B(N13640));
NOR2XL inst_cellmath__220__188__I4168 (.Y(N682), .A(N13545), .B(N13556));
NOR2XL inst_cellmath__220__188__I4169 (.Y(N683), .A(N13545), .B(N13622));
NOR2XL inst_cellmath__220__188__I4170 (.Y(N684), .A(N13545), .B(N13535));
NOR2XL inst_cellmath__220__188__I4171 (.Y(N685), .A(N13545), .B(N13605));
NAND2XL inst_cellmath__220__188__I4172 (.Y(N13588), .A(N13602), .B(N13551));
NOR2XL inst_cellmath__220__188__I4173 (.Y(N686), .A(N13545), .B(N13588));
NOR2XL inst_cellmath__220__188__I4174 (.Y(N687), .A(N13545), .B(N13584));
NOR2XL inst_cellmath__220__188__I4175 (.Y(N688), .A(N13545), .B(N13618));
NOR2XL inst_cellmath__220__188__I4176 (.Y(N689), .A(N13545), .B(N13498));
NOR2XL inst_cellmath__220__188__I4177 (.Y(N690), .A(N13545), .B(N13528));
NOR2XL inst_cellmath__220__188__I4178 (.Y(N691), .A(N13545), .B(N13564));
NOR2XL inst_cellmath__220__188__I4179 (.Y(N692), .A(N13545), .B(N13597));
NOR2XL inst_cellmath__220__188__I4180 (.Y(N693), .A(N13545), .B(N13630));
NOR2XL inst_cellmath__220__188__I4181 (.Y(N694), .A(N13545), .B(N13513));
AOI22XL inst_cellmath__220__188__I4182 (.Y(N695), .A0(N13531), .A1(N13542), .B0(N13509), .B1(N13545));
AOI22XL inst_cellmath__220__188__I4183 (.Y(N696), .A0(N13531), .A1(N13578), .B0(N13575), .B1(N13545));
AOI22XL inst_cellmath__220__188__I4184 (.Y(N697), .A0(N13531), .A1(N13611), .B0(N13640), .B1(N13545));
AOI22XL inst_cellmath__220__188__I4185 (.Y(N698), .A0(N13531), .A1(N13491), .B0(N13556), .B1(N13545));
AOI22XL inst_cellmath__220__188__I4186 (.Y(N699), .A0(N13531), .A1(N13522), .B0(N13622), .B1(N13545));
AOI22XL inst_cellmath__220__188__I4187 (.Y(N700), .A0(N13531), .A1(N13558), .B0(N13535), .B1(N13545));
AOI22XL inst_cellmath__220__188__I4188 (.Y(N701), .A0(N13531), .A1(N13591), .B0(N13605), .B1(N13545));
NOR2X1 inst_cellmath__220_2WWMM_I4194 (.Y(N13822), .A(inst_cellmath__219), .B(N639));
AOI22XL inst_cellmath__220_2WWMM_I4195 (.Y(N13800), .A0(a_exp[0]), .A1(N639), .B0(N13822), .B1(N13601));
AOI22XL inst_cellmath__220_2WWMM_I4196 (.Y(N13845), .A0(a_exp[1]), .A1(N639), .B0(N13822), .B1(N13594));
AOI22XL inst_cellmath__220_2WWMM_I4197 (.Y(N13786), .A0(a_exp[2]), .A1(N639), .B0(N13822), .B1(N13549));
AOI22XL inst_cellmath__220_2WWMM_I4198 (.Y(N13832), .A0(a_exp[3]), .A1(N639), .B0(N13822), .B1(N13551));
AOI22XL inst_cellmath__220_2WWMM_I4199 (.Y(N13877), .A0(a_exp[4]), .A1(N639), .B0(N13822), .B1(N13531));
AOI21XL inst_cellmath__220_2WWMM_I4200 (.Y(N13818), .A0(a_exp[5]), .A1(N639), .B0(N13822));
AOI21XL inst_cellmath__220_2WWMM_I4201 (.Y(N13863), .A0(a_exp[6]), .A1(N639), .B0(N13822));
AND2XL inst_cellmath__220_2WWMM_I4202 (.Y(N647), .A(a_exp[7]), .B(N639));
AO22XL inst_cellmath__220_2WWMM_I4203 (.Y(N648), .A0(N639), .A1(a_man[0]), .B0(N13822), .B1(N679));
AO22XL inst_cellmath__220_2WWMM_I4204 (.Y(N649), .A0(N639), .A1(a_man[1]), .B0(N13822), .B1(N680));
AO22XL inst_cellmath__220_2WWMM_I4205 (.Y(N650), .A0(N639), .A1(a_man[2]), .B0(N13822), .B1(N681));
AO22XL inst_cellmath__220_2WWMM_I4206 (.Y(N651), .A0(N639), .A1(a_man[3]), .B0(N13822), .B1(N682));
AO22XL inst_cellmath__220_2WWMM_I4207 (.Y(N652), .A0(N639), .A1(a_man[4]), .B0(N13822), .B1(N683));
AO22XL inst_cellmath__220_2WWMM_I4208 (.Y(N653), .A0(N639), .A1(a_man[5]), .B0(N13822), .B1(N684));
AO22XL inst_cellmath__220_2WWMM_I4209 (.Y(N654), .A0(N639), .A1(a_man[6]), .B0(N13822), .B1(N685));
AO22XL inst_cellmath__220_2WWMM_I4210 (.Y(N655), .A0(N639), .A1(a_man[7]), .B0(N13822), .B1(N686));
AO22XL inst_cellmath__220_2WWMM_I4211 (.Y(N656), .A0(N639), .A1(a_man[8]), .B0(N13822), .B1(N687));
AO22XL inst_cellmath__220_2WWMM_I4212 (.Y(N657), .A0(N639), .A1(a_man[9]), .B0(N13822), .B1(N688));
AO22XL inst_cellmath__220_2WWMM_I4213 (.Y(N658), .A0(N639), .A1(a_man[10]), .B0(N13822), .B1(N689));
AO22XL inst_cellmath__220_2WWMM_I4214 (.Y(N659), .A0(N639), .A1(a_man[11]), .B0(N13822), .B1(N690));
AO22XL inst_cellmath__220_2WWMM_I4215 (.Y(N660), .A0(N639), .A1(a_man[12]), .B0(N13822), .B1(N691));
AO22XL inst_cellmath__220_2WWMM_I4216 (.Y(N661), .A0(N639), .A1(a_man[13]), .B0(N13822), .B1(N692));
AO22XL inst_cellmath__220_2WWMM_I4217 (.Y(N662), .A0(N639), .A1(a_man[14]), .B0(N13822), .B1(N693));
AO22XL inst_cellmath__220_2WWMM_I4218 (.Y(N663), .A0(N639), .A1(a_man[15]), .B0(N13822), .B1(N694));
AO22XL inst_cellmath__220_2WWMM_I4219 (.Y(N664), .A0(N639), .A1(a_man[16]), .B0(N13822), .B1(N695));
AO22XL inst_cellmath__220_2WWMM_I4220 (.Y(N665), .A0(N639), .A1(a_man[17]), .B0(N13822), .B1(N696));
AO22XL inst_cellmath__220_2WWMM_I4221 (.Y(N666), .A0(N639), .A1(a_man[18]), .B0(N13822), .B1(N697));
AO22XL inst_cellmath__220_2WWMM_I4222 (.Y(N667), .A0(N639), .A1(a_man[19]), .B0(N13822), .B1(N698));
AO22XL inst_cellmath__220_2WWMM_I4223 (.Y(N668), .A0(N639), .A1(a_man[20]), .B0(N13822), .B1(N699));
AO22XL inst_cellmath__220_2WWMM_I4224 (.Y(N669), .A0(N639), .A1(a_man[21]), .B0(N13822), .B1(N700));
AO22XL inst_cellmath__220_2WWMM_I4225 (.Y(N670), .A0(N639), .A1(a_man[22]), .B0(N13822), .B1(N701));
NAND2BXL inst_cellmath__220_2WWMM_I4226 (.Y(N13809), .AN(N639), .B(inst_cellmath__219));
NAND2XL inst_cellmath__220_2WWMM_I4227 (.Y(N640), .A(N13809), .B(N13800));
NAND2XL inst_cellmath__220_2WWMM_I4228 (.Y(N641), .A(N13809), .B(N13845));
NAND2XL inst_cellmath__220_2WWMM_I4229 (.Y(N642), .A(N13809), .B(N13786));
NAND2XL inst_cellmath__220_2WWMM_I4230 (.Y(N643), .A(N13809), .B(N13832));
NAND2XL inst_cellmath__220_2WWMM_I4231 (.Y(N644), .A(N13809), .B(N13877));
NAND2XL inst_cellmath__220_2WWMM_I4232 (.Y(N645), .A(N13809), .B(N13818));
NAND2XL inst_cellmath__220_2WWMM_I4233 (.Y(N646), .A(N13809), .B(N13863));
OR4X1 inst_cellmath__223__208__I4234 (.Y(N13925), .A(N647), .B(N645), .C(N646), .D(N640));
NOR3XL inst_cellmath__223__208__I4235 (.Y(N13957), .A(N13925), .B(N641), .C(N642));
NOR2XL inst_cellmath__223__208__I4236 (.Y(N13969), .A(N643), .B(N644));
NAND3BXL inst_cellmath__223__208__I4237 (.Y(N13939), .AN(N648), .B(N13957), .C(N13969));
NOR4X1 inst_cellmath__223__208__I4238 (.Y(N13955), .A(N649), .B(N650), .C(N13939), .D(N654));
NOR3XL inst_cellmath__223__208__I4239 (.Y(N13937), .A(N651), .B(N655), .C(N658));
NOR3XL inst_cellmath__223__208__I4242 (.Y(N13943), .A(N653), .B(N652), .C(N663));
NOR3BXL inst_cellmath__223__208__I4246 (.Y(N13934), .AN(N13955), .B(N657), .C(N662));
OR4X1 inst_cellmath__223__208__I23843 (.Y(N13947), .A(N659), .B(N656), .C(N661), .D(N660));
NOR4BX1 inst_cellmath__223__208__I23845 (.Y(N13940), .AN(N13937), .B(N669), .C(N13947), .D(N664));
OR4X1 inst_cellmath__223__208__I23844 (.Y(N13970), .A(N667), .B(N665), .C(N668), .D(N666));
NAND4BXL inst_cellmath__223__208__I23846 (.Y(N578), .AN(N13970), .B(N13943), .C(N13940), .D(N13934));
XOR2XL cynw_cm_float_sin_I4254 (.Y(N577), .A(a_sign), .B(N757));
NOR4BBX1 cynw_cm_float_sin_I8487 (.Y(N579), .AN(N577), .BN(N578), .C(inst_cellmath__82), .D(N487));
MX2XL cynw_cm_float_sin_I4257 (.Y(x[31]), .A(N579), .B(a_sign), .S0(N639));
NAND2BXL cynw_cm_float_sin_I4258 (.Y(N580), .AN(inst_cellmath__82), .B(N487));
INVXL inst_cellmath__228_0_I4259 (.Y(N14019), .A(N759));
INVXL inst_cellmath__228_0_I4260 (.Y(N14026), .A(N14019));
MX2XL inst_cellmath__228_0_I4261 (.Y(x[23]), .A(N640), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4262 (.Y(x[24]), .A(N641), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4263 (.Y(x[25]), .A(N642), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4264 (.Y(x[26]), .A(N643), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4265 (.Y(x[27]), .A(N644), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4266 (.Y(x[28]), .A(N645), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4267 (.Y(x[29]), .A(N646), .B(N580), .S0(N14026));
MX2XL inst_cellmath__228_0_I4268 (.Y(x[30]), .A(N647), .B(N580), .S0(N14026));
MX2XL inst_cellmath__231_0_I4269 (.Y(x[0]), .A(N648), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4270 (.Y(x[1]), .A(N649), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4271 (.Y(x[2]), .A(N650), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4272 (.Y(x[3]), .A(N651), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4273 (.Y(x[4]), .A(N652), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4274 (.Y(x[5]), .A(N653), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4275 (.Y(x[6]), .A(N654), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4276 (.Y(x[7]), .A(N655), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4277 (.Y(x[8]), .A(N656), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4278 (.Y(x[9]), .A(N657), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4279 (.Y(x[10]), .A(N658), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4280 (.Y(x[11]), .A(N659), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4281 (.Y(x[12]), .A(N660), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4282 (.Y(x[13]), .A(N661), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4283 (.Y(x[14]), .A(N662), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4284 (.Y(x[15]), .A(N663), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4285 (.Y(x[16]), .A(N664), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4286 (.Y(x[17]), .A(N665), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4287 (.Y(x[18]), .A(N666), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4288 (.Y(x[19]), .A(N667), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4289 (.Y(x[20]), .A(N668), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4290 (.Y(x[21]), .A(N669), .B(inst_cellmath__82), .S0(N759));
MX2XL inst_cellmath__231_0_I4291 (.Y(x[22]), .A(N670), .B(inst_cellmath__82), .S0(N759));
assign inst_cellmath__42[2] = 1'B0;
assign inst_cellmath__42[3] = 1'B0;
assign inst_cellmath__42[6] = 1'B0;
assign inst_cellmath__42[7] = 1'B0;
assign inst_cellmath__42[8] = 1'B0;
assign inst_cellmath__61[0] = 1'B0;
assign inst_cellmath__61[16] = 1'B0;
assign inst_cellmath__195[29] = 1'B0;
assign inst_cellmath__198[0] = 1'B0;
assign inst_cellmath__198[1] = 1'B0;
assign inst_cellmath__198[2] = 1'B0;
assign inst_cellmath__198[3] = 1'B0;
assign inst_cellmath__198[4] = 1'B0;
assign inst_cellmath__198[5] = 1'B0;
assign inst_cellmath__198[6] = 1'B0;
assign inst_cellmath__198[7] = 1'B0;
assign inst_cellmath__198[8] = 1'B0;
assign inst_cellmath__198[9] = 1'B0;
assign inst_cellmath__198[10] = 1'B0;
assign inst_cellmath__198[11] = 1'B0;
assign inst_cellmath__198[12] = 1'B0;
assign inst_cellmath__198[13] = 1'B0;
assign inst_cellmath__198[14] = 1'B0;
assign inst_cellmath__198[15] = 1'B0;
assign inst_cellmath__198[16] = 1'B0;
assign inst_cellmath__198[17] = 1'B0;
assign inst_cellmath__201[0] = 1'B0;
assign inst_cellmath__201[1] = 1'B0;
assign inst_cellmath__201[2] = 1'B0;
assign inst_cellmath__201[3] = 1'B0;
assign inst_cellmath__201[4] = 1'B0;
assign inst_cellmath__201[5] = 1'B0;
assign inst_cellmath__201[6] = 1'B0;
assign inst_cellmath__201[7] = 1'B0;
assign inst_cellmath__201[8] = 1'B0;
assign inst_cellmath__201[9] = 1'B0;
assign inst_cellmath__201[10] = 1'B0;
assign inst_cellmath__201[11] = 1'B0;
assign inst_cellmath__201[12] = 1'B0;
assign inst_cellmath__201[13] = 1'B0;
assign inst_cellmath__201[14] = 1'B0;
assign inst_cellmath__201[15] = 1'B0;
assign inst_cellmath__201[16] = 1'B0;
assign inst_cellmath__201[17] = 1'B0;
assign inst_cellmath__201[18] = 1'B0;
assign inst_cellmath__201[19] = 1'B0;
assign inst_cellmath__201[20] = 1'B0;
assign inst_cellmath__201[21] = 1'B0;
assign inst_cellmath__201[22] = 1'B0;
assign inst_cellmath__201[23] = 1'B0;
assign inst_cellmath__201[24] = 1'B0;
assign inst_cellmath__201[49] = 1'B0;
assign inst_cellmath__203__W0[0] = 1'B0;
assign inst_cellmath__203__W0[43] = 1'B1;
assign inst_cellmath__203__W0[44] = 1'B1;
assign inst_cellmath__203__W0[45] = 1'B1;
assign inst_cellmath__203__W0[46] = 1'B1;
assign inst_cellmath__203__W1[0] = 1'B0;
assign inst_cellmath__203__W1[43] = 1'B0;
assign inst_cellmath__203__W1[44] = 1'B0;
assign inst_cellmath__203__W1[45] = 1'B0;
assign inst_cellmath__203__W1[46] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign inst_cellmath__215[1] = 1'B0;
assign inst_cellmath__215[2] = 1'B0;
assign inst_cellmath__215[4] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  v7L3SgnXoxk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



