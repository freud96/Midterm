/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:12 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_div_ieee_E8_M23_0 (
	clk,
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	accept,
	x
	); /* architecture "gate_level" */ 
input  clk;
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input  accept;
output [31:0] x;
wire [31:0] inst_cellmath__8,
	inst_cellmath__9;
wire  inst_cellmath__11;
wire [3:0] inst_cellmath__12,
	inst_cellmath__13;
wire [25:0] inst_cellmath__14,
	inst_cellmath__16,
	inst_cellmath__17;
wire [4:0] inst_cellmath__22,
	inst_cellmath__23;
wire [6:0] inst_lookup0_cellmath__27;
wire [2:0] inst_lookup0_cellmath__29;
wire [25:0] inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__34,
	inst_cellmath__35,
	inst_cellmath__38__W0,
	inst_cellmath__38__W1,
	inst_cellmath__39__W0,
	inst_cellmath__39__W1;
wire [28:0] inst_cellmath__40,
	inst_cellmath__41,
	inst_cellmath__42,
	inst_cellmath__43,
	inst_cellmath__44,
	inst_cellmath__45,
	inst_cellmath__46,
	inst_cellmath__47;
wire [6:0] inst_it2_lookup1_cellmath__53;
wire [2:0] inst_it2_lookup1_cellmath__55;
wire [25:0] inst_it2_cellmath__56,
	inst_it2_cellmath__57,
	inst_it2_cellmath__60,
	inst_it2_cellmath__61,
	inst_it2_cellmath__62__W0,
	inst_it2_cellmath__62__W1,
	inst_it2_cellmath__63__W1;
wire [9:0] inst_cellmath__67,
	inst_cellmath__68;
wire  inst_cellmath__69,
	inst_cellmath__70,
	inst_cellmath__71,
	inst_cellmath__72,
	inst_cellmath__73,
	inst_cellmath__74,
	inst_cellmath__75,
	inst_cellmath__76,
	inst_cellmath__77,
	inst_cellmath__78,
	inst_cellmath__79,
	inst_cellmath__80,
	inst_cellmath__83,
	inst_cellmath__84,
	inst_cellmath__85,
	inst_cellmath__86,
	inst_cellmath__87,
	inst_cellmath__88,
	inst_cellmath__89,
	inst_cellmath__91,
	inst_cellmath__96,
	inst_cellmath__100,
	inst_cellmath__101,
	inst_cellmath__102,
	inst_cellmath__103,
	inst_cellmath__104,
	inst_cellmath__105,
	inst_cellmath__106,
	inst_cellmath__109;
wire [7:0] inst_cellmath__110,
	inst_cellmath__111;
wire [21:0] inst_cellmath__112;
wire [31:0] inst_cellmath__113;
wire [25:0] inst_cellmath__120;
wire  inst_cellmath__122;
wire [28:0] inst_cellmath__124;
wire [22:0] inst_cellmath__125;
wire  inst_cellmath__126,
	inst_cellmath__127;
wire [22:0] inst_cellmath__129;
wire  inst_cellmath__135,
	inst_cellmath__136,
	inst_cellmath__137;
wire N1322,N1324,N1325,N1326,N1327,N1386,N1387 
	,N1388,N1417,N1555,N1675,N1677,N1678,N1679,N1680 
	,N1681,N1682,N1750,N1751,N1752,N1753,N1754,N1755 
	,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763 
	,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771 
	,N1772,N1922,N2045,N2046,N2047,N2048,N2049,N2050 
	,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058 
	,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066 
	,N2067,N2068,N2150,N2151,N2152,N2153,N2154,N2155 
	,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163 
	,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171 
	,N2172,N2173,N2201,N2202,N2203,N2204,N2205,N2206 
	,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214 
	,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222 
	,N2223,N2224,N2254,N2255,N2256,N2257,N2258,N2259 
	,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267 
	,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275 
	,N2276,N2277,N4587,N4594,N12283,N12286,N12290,N12294 
	,N12297,N12310,N12313,N12314,N12315,N12318,N12322,N12323 
	,N12326,N12362,N12363,N12364,N12365,N12366,N12368,N12369 
	,N12371,N12373,N12375,N12376,N12377,N12378,N12379,N12380 
	,N12381,N12383,N12384,N12385,N12386,N12387,N12389,N12392 
	,N12394,N12395,N12396,N12397,N12399,N12400,N12401,N12403 
	,N12404,N12405,N12407,N12408,N12409,N12410,N12411,N12414 
	,N12417,N12418,N12419,N12421,N12573,N12658,N12720,N12723 
	,N12729,N12732,N12736,N12738,N12740,N12744,N12751,N12754 
	,N12761,N12764,N12771,N12774,N12782,N12785,N12791,N12794 
	,N12797,N12803,N12806,N12811,N12813,N12870,N12983,N13206 
	,N13373,N13376,N13380,N13384,N13387,N13401,N13402,N13403 
	,N13404,N13405,N13408,N13410,N13412,N13414,N13415,N13417 
	,N13419,N13420,N13422,N13423,N13424,N13425,N13426,N13428 
	,N13431,N13433,N13434,N13435,N13436,N13438,N13439,N13440 
	,N13442,N13444,N13447,N13448,N13449,N13450,N13453,N13456 
	,N13457,N13458,N13460,N13614,N13658,N13661,N13665,N13667 
	,N13673,N13677,N13680,N13685,N13689,N13692,N13697,N13704 
	,N13705,N13712,N13716,N13719,N13722,N13725,N13730,N13737 
	,N13738,N13745,N13750,N13753,N13758,N13935,N13952,N14010 
	,N14012,N14016,N14018,N14020,N14025,N14027,N14030,N14033 
	,N14035,N14038,N14043,N14045,N14047,N14053,N14055,N14058 
	,N14061,N14063,N14070,N14072,N14077,N14146,N14149,N14153 
	,N14158,N14160,N14165,N14169,N14173,N14177,N14179,N14181 
	,N14182,N14185,N14213,N14214,N14594,N14648,N14981,N15334 
	,N15398,N15400,N15401,N15403,N15404,N15406,N15409,N15411 
	,N15412,N15413,N15415,N15417,N15418,N15421,N15423,N15424 
	,N15426,N15429,N15430,N15431,N15432,N15434,N15435,N15436 
	,N15440,N15443,N15444,N15486,N15491,N15495,N15497,N15503 
	,N15504,N15506,N15511,N15518,N15523,N15552,N15554,N15560 
	,N15579,N15582,N15583,N15585,N15589,N15605,N15608,N15618 
	,N15631,N15636,N15640,N15656,N15660,N15663,N15666,N15679 
	,N15681,N15699,N15702,N15710,N15711,N15720,N15722,N15724 
	,N15726,N15728,N15730,N15732,N15733,N15736,N15758,N15759 
	,N15762,N15770,N15779,N15780,N15782,N15784,N15786,N15788 
	,N15790,N15792,N15795,N15830,N15834,N15837,N15840,N15848 
	,N15852,N15855,N15858,N15898,N15943,N15964,N16014,N16016 
	,N16019,N16030,N16033,N16051,N16052,N16055,N16059,N16064 
	,N16067,N16070,N16076,N16080,N16083,N16086,N16122,N16178 
	,N18408,N18417,N28016,N28021,N28027;
EDFFHQX1 inst_cellmath__0_0_0__I0 (.Q(x[0]), .D(inst_cellmath__113[0]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_1__I1 (.Q(x[1]), .D(inst_cellmath__113[1]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_2__I2 (.Q(x[2]), .D(inst_cellmath__113[2]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_3__I3 (.Q(x[3]), .D(inst_cellmath__113[3]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_4__I4 (.Q(x[4]), .D(inst_cellmath__113[4]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_5__I5 (.Q(x[5]), .D(inst_cellmath__113[5]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_6__I6 (.Q(x[6]), .D(inst_cellmath__113[6]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_7__I7 (.Q(x[7]), .D(inst_cellmath__113[7]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_8__I8 (.Q(x[8]), .D(inst_cellmath__113[8]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_9__I9 (.Q(x[9]), .D(inst_cellmath__113[9]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_10__I10 (.Q(x[10]), .D(inst_cellmath__113[10]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_11__I11 (.Q(x[11]), .D(inst_cellmath__113[11]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_12__I12 (.Q(x[12]), .D(inst_cellmath__113[12]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_13__I13 (.Q(x[13]), .D(inst_cellmath__113[13]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_14__I14 (.Q(x[14]), .D(inst_cellmath__113[14]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_15__I15 (.Q(x[15]), .D(inst_cellmath__113[15]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_16__I16 (.Q(x[16]), .D(inst_cellmath__113[16]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_17__I17 (.Q(x[17]), .D(inst_cellmath__113[17]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_18__I18 (.Q(x[18]), .D(inst_cellmath__113[18]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_19__I19 (.Q(x[19]), .D(inst_cellmath__113[19]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_20__I20 (.Q(x[20]), .D(inst_cellmath__113[20]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_21__I21 (.Q(x[21]), .D(inst_cellmath__113[21]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_22__I22 (.Q(x[22]), .D(inst_cellmath__113[22]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_23__I23 (.Q(x[23]), .D(inst_cellmath__113[23]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_24__I24 (.Q(x[24]), .D(inst_cellmath__113[24]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_25__I25 (.Q(x[25]), .D(inst_cellmath__113[25]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_26__I26 (.Q(x[26]), .D(inst_cellmath__113[26]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_27__I27 (.Q(x[27]), .D(inst_cellmath__113[27]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_28__I28 (.Q(x[28]), .D(inst_cellmath__113[28]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_29__I29 (.Q(x[29]), .D(inst_cellmath__113[29]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_30__I30 (.Q(x[30]), .D(inst_cellmath__113[30]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_31__I31 (.Q(x[31]), .D(inst_cellmath__113[31]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_0__I32 (.Q(inst_cellmath__9[0]), .D(b_man[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_1__I33 (.Q(inst_cellmath__9[1]), .D(b_man[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_2__I34 (.Q(inst_cellmath__9[2]), .D(b_man[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_3__I35 (.Q(inst_cellmath__9[3]), .D(b_man[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_4__I36 (.Q(inst_cellmath__9[4]), .D(b_man[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_5__I37 (.Q(inst_cellmath__9[5]), .D(b_man[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_6__I38 (.Q(inst_cellmath__9[6]), .D(b_man[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_7__I39 (.Q(inst_cellmath__9[7]), .D(b_man[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_8__I40 (.Q(inst_cellmath__9[8]), .D(b_man[8]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_9__I41 (.Q(inst_cellmath__9[9]), .D(b_man[9]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_10__I42 (.Q(inst_cellmath__9[10]), .D(b_man[10]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_11__I43 (.Q(inst_cellmath__9[11]), .D(b_man[11]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_12__I44 (.Q(inst_cellmath__9[12]), .D(b_man[12]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_13__I45 (.Q(inst_cellmath__9[13]), .D(b_man[13]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_14__I46 (.Q(inst_cellmath__9[14]), .D(b_man[14]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_15__I47 (.Q(inst_cellmath__9[15]), .D(b_man[15]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_16__I48 (.Q(inst_cellmath__9[16]), .D(b_man[16]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_17__I49 (.Q(inst_cellmath__9[17]), .D(b_man[17]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_18__I50 (.Q(inst_cellmath__9[18]), .D(b_man[18]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_19__I51 (.Q(inst_cellmath__9[19]), .D(b_man[19]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_20__I52 (.Q(inst_cellmath__9[20]), .D(b_man[20]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_21__I53 (.Q(inst_it2_lookup1_cellmath__53[0]), .D(b_man[21]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_22__I54 (.Q(inst_it2_lookup1_cellmath__53[1]), .D(b_man[22]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_23__I55 (.Q(inst_cellmath__9[23]), .D(b_exp[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_24__I56 (.Q(inst_cellmath__9[24]), .D(b_exp[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_25__I57 (.Q(inst_cellmath__9[25]), .D(b_exp[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_26__I58 (.Q(inst_cellmath__9[26]), .D(b_exp[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_27__I59 (.Q(inst_cellmath__9[27]), .D(b_exp[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_28__I60 (.Q(inst_cellmath__9[28]), .D(b_exp[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_29__I61 (.Q(inst_cellmath__9[29]), .D(b_exp[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_30__I62 (.Q(inst_cellmath__9[30]), .D(b_exp[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_31__I63 (.Q(inst_cellmath__9[31]), .D(b_sign), .E(accept), .CK(clk));
DFFQXL inst_cellmath__11_0_I64 (.Q(inst_cellmath__11), .D(accept), .CK(clk));
DFFQXL inst_cellmath__16_0_1__I65 (.Q(inst_cellmath__16[1]), .D(inst_cellmath__14[1]), .CK(clk));
DFFQXL inst_cellmath__16_0_2__I66 (.Q(inst_cellmath__16[2]), .D(inst_cellmath__14[2]), .CK(clk));
DFFQXL inst_cellmath__16_0_3__I67 (.Q(inst_cellmath__16[3]), .D(inst_cellmath__14[3]), .CK(clk));
DFFQXL inst_cellmath__16_0_4__I68 (.Q(inst_cellmath__16[4]), .D(inst_cellmath__14[4]), .CK(clk));
DFFQXL inst_cellmath__16_0_5__I69 (.Q(inst_cellmath__16[5]), .D(inst_cellmath__14[5]), .CK(clk));
DFFQXL inst_cellmath__16_0_6__I70 (.Q(inst_cellmath__16[6]), .D(inst_cellmath__14[6]), .CK(clk));
DFFQXL inst_cellmath__16_0_7__I71 (.Q(inst_cellmath__16[7]), .D(inst_cellmath__14[7]), .CK(clk));
DFFQXL inst_cellmath__16_0_8__I72 (.Q(inst_cellmath__16[8]), .D(inst_cellmath__14[8]), .CK(clk));
DFFQXL inst_cellmath__16_0_9__I73 (.Q(inst_cellmath__16[9]), .D(inst_cellmath__14[9]), .CK(clk));
DFFQXL inst_cellmath__16_0_10__I74 (.Q(inst_cellmath__16[10]), .D(inst_cellmath__14[10]), .CK(clk));
DFFQXL inst_cellmath__16_0_11__I75 (.Q(inst_cellmath__16[11]), .D(inst_cellmath__14[11]), .CK(clk));
DFFQXL inst_cellmath__16_0_12__I76 (.Q(inst_cellmath__16[12]), .D(inst_cellmath__14[12]), .CK(clk));
DFFQXL inst_cellmath__16_0_13__I77 (.Q(inst_cellmath__16[13]), .D(inst_cellmath__14[13]), .CK(clk));
DFFQXL inst_cellmath__16_0_14__I78 (.Q(inst_cellmath__16[14]), .D(inst_cellmath__14[14]), .CK(clk));
DFFQXL inst_cellmath__16_0_15__I79 (.Q(inst_cellmath__16[15]), .D(inst_cellmath__14[15]), .CK(clk));
DFFQXL inst_cellmath__16_0_16__I80 (.Q(inst_cellmath__16[16]), .D(inst_cellmath__14[16]), .CK(clk));
DFFQXL inst_cellmath__16_0_17__I81 (.Q(inst_cellmath__16[17]), .D(inst_cellmath__14[17]), .CK(clk));
DFFQXL inst_cellmath__16_0_18__I82 (.Q(inst_cellmath__16[18]), .D(inst_cellmath__14[18]), .CK(clk));
DFFQXL inst_cellmath__16_0_19__I83 (.Q(inst_cellmath__16[19]), .D(inst_cellmath__14[19]), .CK(clk));
DFFQXL inst_cellmath__16_0_20__I84 (.Q(inst_cellmath__16[20]), .D(inst_cellmath__14[20]), .CK(clk));
DFFQXL inst_cellmath__16_0_21__I85 (.Q(inst_cellmath__16[21]), .D(inst_cellmath__14[21]), .CK(clk));
DFFQXL inst_cellmath__16_0_22__I86 (.Q(inst_cellmath__16[22]), .D(inst_cellmath__14[22]), .CK(clk));
DFFQXL inst_cellmath__16_0_23__I87 (.Q(inst_cellmath__16[23]), .D(inst_cellmath__14[23]), .CK(clk));
DFFQXL inst_cellmath__16_0_24__I88 (.Q(inst_cellmath__16[24]), .D(inst_cellmath__14[24]), .CK(clk));
DFFQXL inst_cellmath__16_0_25__I89 (.Q(inst_cellmath__16[25]), .D(inst_cellmath__14[25]), .CK(clk));
DFFQXL inst_cellmath__17_0_1__I91 (.Q(inst_cellmath__17[1]), .D(inst_it2_cellmath__63__W1[1]), .CK(clk));
DFFQXL inst_cellmath__17_0_2__I92 (.Q(inst_cellmath__17[2]), .D(inst_it2_cellmath__63__W1[2]), .CK(clk));
DFFQXL inst_cellmath__17_0_3__I93 (.Q(inst_cellmath__17[3]), .D(inst_it2_cellmath__63__W1[3]), .CK(clk));
DFFQXL inst_cellmath__17_0_4__I94 (.Q(inst_cellmath__17[4]), .D(inst_it2_cellmath__63__W1[4]), .CK(clk));
DFFQXL inst_cellmath__17_0_5__I95 (.Q(inst_cellmath__17[5]), .D(inst_it2_cellmath__63__W1[5]), .CK(clk));
DFFQXL inst_cellmath__17_0_6__I96 (.Q(inst_cellmath__17[6]), .D(inst_it2_cellmath__63__W1[6]), .CK(clk));
DFFQXL inst_cellmath__17_0_7__I97 (.Q(inst_cellmath__17[7]), .D(inst_it2_cellmath__63__W1[7]), .CK(clk));
DFFQXL inst_cellmath__17_0_8__I98 (.Q(inst_cellmath__17[8]), .D(inst_it2_cellmath__63__W1[8]), .CK(clk));
DFFQXL inst_cellmath__17_0_9__I99 (.Q(inst_cellmath__17[9]), .D(inst_it2_cellmath__63__W1[9]), .CK(clk));
DFFQXL inst_cellmath__17_0_10__I100 (.Q(inst_cellmath__17[10]), .D(inst_it2_cellmath__63__W1[10]), .CK(clk));
DFFQXL inst_cellmath__17_0_11__I101 (.Q(inst_cellmath__17[11]), .D(inst_it2_cellmath__63__W1[11]), .CK(clk));
DFFQXL inst_cellmath__17_0_12__I102 (.Q(inst_cellmath__17[12]), .D(inst_it2_cellmath__63__W1[12]), .CK(clk));
DFFQXL inst_cellmath__17_0_13__I103 (.Q(inst_cellmath__17[13]), .D(inst_it2_cellmath__63__W1[13]), .CK(clk));
DFFQXL inst_cellmath__17_0_14__I104 (.Q(inst_cellmath__17[14]), .D(inst_it2_cellmath__63__W1[14]), .CK(clk));
DFFQXL inst_cellmath__17_0_15__I105 (.Q(inst_cellmath__17[15]), .D(inst_it2_cellmath__63__W1[15]), .CK(clk));
DFFQXL inst_cellmath__17_0_16__I106 (.Q(inst_cellmath__17[16]), .D(inst_it2_cellmath__63__W1[16]), .CK(clk));
DFFQXL inst_cellmath__17_0_17__I107 (.Q(inst_cellmath__17[17]), .D(inst_it2_cellmath__63__W1[17]), .CK(clk));
DFFQXL inst_cellmath__17_0_18__I108 (.Q(inst_cellmath__17[18]), .D(inst_it2_cellmath__63__W1[18]), .CK(clk));
DFFQXL inst_cellmath__17_0_19__I109 (.Q(inst_cellmath__17[19]), .D(inst_it2_cellmath__63__W1[19]), .CK(clk));
DFFQXL inst_cellmath__17_0_20__I110 (.Q(inst_cellmath__17[20]), .D(inst_it2_cellmath__63__W1[20]), .CK(clk));
DFFQXL inst_cellmath__17_0_21__I111 (.Q(inst_cellmath__17[21]), .D(inst_it2_cellmath__63__W1[21]), .CK(clk));
DFFQXL inst_cellmath__17_0_22__I112 (.Q(inst_cellmath__17[22]), .D(inst_it2_cellmath__63__W1[22]), .CK(clk));
DFFQXL inst_cellmath__17_0_23__I113 (.Q(inst_cellmath__17[23]), .D(inst_it2_cellmath__63__W1[23]), .CK(clk));
DFFQXL inst_cellmath__17_0_24__I114 (.Q(inst_cellmath__17[24]), .D(inst_it2_cellmath__63__W1[24]), .CK(clk));
DFFQXL inst_cellmath__17_0_25__I115 (.Q(inst_cellmath__17[25]), .D(inst_it2_cellmath__63__W1[25]), .CK(clk));
ADDHX1 inst_cellmath__23_0_I1788 (.CO(N12290), .S(inst_cellmath__23[0]), .A(inst_cellmath__17[21]), .B(inst_cellmath__16[21]));
ADDFX1 inst_cellmath__23_0_I1789 (.CO(N12286), .S(inst_cellmath__23[1]), .A(inst_cellmath__16[22]), .B(inst_cellmath__17[22]), .CI(N12290));
ADDFX1 inst_cellmath__23_0_I1790 (.CO(N12297), .S(inst_cellmath__23[2]), .A(inst_cellmath__16[23]), .B(inst_cellmath__17[23]), .CI(N12286));
ADDFX1 inst_cellmath__23_0_I1791 (.CO(N12283), .S(inst_cellmath__23[3]), .A(inst_cellmath__16[24]), .B(inst_cellmath__17[24]), .CI(N12297));
ADDFX1 inst_cellmath__23_0_I1792 (.CO(N12294), .S(inst_cellmath__23[4]), .A(inst_cellmath__16[25]), .B(inst_cellmath__17[25]), .CI(N12283));
EDFFHQX1 inst_cellmath__8_0_0__I117 (.Q(inst_cellmath__8[0]), .D(a_man[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_1__I118 (.Q(inst_cellmath__8[1]), .D(a_man[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_2__I119 (.Q(inst_cellmath__8[2]), .D(a_man[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_3__I120 (.Q(inst_cellmath__8[3]), .D(a_man[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_4__I121 (.Q(inst_cellmath__8[4]), .D(a_man[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_5__I122 (.Q(inst_cellmath__8[5]), .D(a_man[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_6__I123 (.Q(inst_cellmath__8[6]), .D(a_man[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_7__I124 (.Q(inst_cellmath__8[7]), .D(a_man[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_8__I125 (.Q(inst_cellmath__8[8]), .D(a_man[8]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_9__I126 (.Q(inst_cellmath__8[9]), .D(a_man[9]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_10__I127 (.Q(inst_cellmath__8[10]), .D(a_man[10]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_11__I128 (.Q(inst_cellmath__8[11]), .D(a_man[11]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_12__I129 (.Q(inst_cellmath__8[12]), .D(a_man[12]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_13__I130 (.Q(inst_cellmath__8[13]), .D(a_man[13]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_14__I131 (.Q(inst_cellmath__8[14]), .D(a_man[14]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_15__I132 (.Q(inst_cellmath__8[15]), .D(a_man[15]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_16__I133 (.Q(inst_cellmath__8[16]), .D(a_man[16]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_17__I134 (.Q(inst_cellmath__8[17]), .D(a_man[17]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_18__I135 (.Q(inst_cellmath__8[18]), .D(a_man[18]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_19__I136 (.Q(inst_cellmath__8[19]), .D(a_man[19]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_20__I137 (.Q(inst_cellmath__8[20]), .D(a_man[20]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_21__I138 (.Q(inst_cellmath__8[21]), .D(a_man[21]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_22__I139 (.Q(inst_cellmath__8[22]), .D(a_man[22]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_23__I140 (.Q(inst_cellmath__8[23]), .D(a_exp[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_24__I141 (.Q(inst_cellmath__8[24]), .D(a_exp[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_25__I142 (.Q(inst_cellmath__8[25]), .D(a_exp[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_26__I143 (.Q(inst_cellmath__8[26]), .D(a_exp[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_27__I144 (.Q(inst_cellmath__8[27]), .D(a_exp[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_28__I145 (.Q(inst_cellmath__8[28]), .D(a_exp[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_29__I146 (.Q(inst_cellmath__8[29]), .D(a_exp[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_30__I147 (.Q(inst_cellmath__8[30]), .D(a_exp[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_31__I148 (.Q(inst_cellmath__8[31]), .D(a_sign), .E(accept), .CK(clk));
INVXL cynw_cm_float_div_ieee_I149 (.Y(N1386), .A(inst_cellmath__9[20]));
INVXL cynw_cm_float_div_ieee_I150 (.Y(N1387), .A(inst_it2_lookup1_cellmath__53[0]));
INVXL cynw_cm_float_div_ieee_I151 (.Y(N1388), .A(inst_it2_lookup1_cellmath__53[1]));
NAND2XL inst_cellmath__22_0_I1793 (.Y(N12322), .A(inst_cellmath__8[20]), .B(N1386));
NOR2XL inst_cellmath__22_0_I1794 (.Y(N12326), .A(inst_cellmath__8[21]), .B(N1387));
NAND2XL inst_cellmath__22_0_I1795 (.Y(N12313), .A(inst_cellmath__8[21]), .B(N1387));
NOR2XL inst_cellmath__22_0_I1796 (.Y(N12315), .A(inst_cellmath__8[22]), .B(N1388));
NAND2XL inst_cellmath__22_0_I1797 (.Y(N12318), .A(inst_cellmath__8[22]), .B(N1388));
AO21XL inst_cellmath__22_0_I1798 (.Y(N12314), .A0(N12313), .A1(N12322), .B0(N12326));
AO21XL inst_cellmath__22_0_I1799 (.Y(inst_cellmath__22[4]), .A0(N12318), .A1(N12314), .B0(N12315));
NAND2BXL inst_cellmath__22_0_I1800 (.Y(N12310), .AN(N12326), .B(N12313));
NAND2BXL inst_cellmath__22_0_I1801 (.Y(N12323), .AN(N12315), .B(N12318));
XOR2XL inst_cellmath__22_0_I1802 (.Y(inst_cellmath__22[0]), .A(inst_cellmath__8[20]), .B(N1386));
XOR2XL inst_cellmath__22_0_I1803 (.Y(inst_cellmath__22[1]), .A(N12322), .B(N12310));
XOR2XL inst_cellmath__22_0_I1804 (.Y(inst_cellmath__22[2]), .A(N12314), .B(N12323));
MX2XL inst_cellmath__24_0_I1805 (.Y(inst_lookup0_cellmath__27[2]), .A(inst_cellmath__23[0]), .B(inst_cellmath__22[0]), .S0(inst_cellmath__11));
MX2XL inst_cellmath__24_0_I1806 (.Y(inst_lookup0_cellmath__27[3]), .A(inst_cellmath__23[1]), .B(inst_cellmath__22[1]), .S0(inst_cellmath__11));
MX2XL inst_cellmath__24_0_I1807 (.Y(inst_lookup0_cellmath__27[4]), .A(inst_cellmath__23[2]), .B(inst_cellmath__22[2]), .S0(inst_cellmath__11));
MX2XL inst_cellmath__24_0_I1808 (.Y(inst_lookup0_cellmath__27[5]), .A(inst_cellmath__23[3]), .B(inst_cellmath__22[4]), .S0(inst_cellmath__11));
MX2XL inst_cellmath__24_0_I1809 (.Y(inst_lookup0_cellmath__27[6]), .A(inst_cellmath__23[4]), .B(inst_cellmath__22[4]), .S0(inst_cellmath__11));
INVXL inst_lookup0_cellmath__29_0_I1812 (.Y(N12397), .A(inst_lookup0_cellmath__27[2]));
INVXL inst_lookup0_cellmath__29_0_I1813 (.Y(N12386), .A(inst_lookup0_cellmath__27[3]));
NOR2XL inst_lookup0_cellmath__29_0_I1814 (.Y(N12381), .A(N12386), .B(N12397));
NOR2XL inst_lookup0_cellmath__29_0_I1815 (.Y(N12418), .A(N12397), .B(N1388));
NAND2XL inst_lookup0_cellmath__29_0_I1816 (.Y(N12379), .A(N1387), .B(N1388));
AOI22XL inst_lookup0_cellmath__29_0_I1817 (.Y(N12366), .A0(N12397), .A1(inst_it2_lookup1_cellmath__53[1]), .B0(N12379), .B1(inst_lookup0_cellmath__27[2]));
AOI22XL inst_lookup0_cellmath__29_0_I1818 (.Y(N12421), .A0(N12386), .A1(N12366), .B0(N12418), .B1(inst_lookup0_cellmath__27[3]));
NAND2XL inst_lookup0_cellmath__29_0_I1819 (.Y(N12365), .A(inst_it2_lookup1_cellmath__53[1]), .B(inst_lookup0_cellmath__27[2]));
NOR2XL inst_lookup0_cellmath__29_0_I1820 (.Y(N12373), .A(N12386), .B(N12365));
INVXL inst_lookup0_cellmath__29_0_I1821 (.Y(N12363), .A(inst_lookup0_cellmath__27[4]));
AOI22XL inst_lookup0_cellmath__29_0_I1822 (.Y(N12394), .A0(N12363), .A1(N12421), .B0(N12381), .B1(inst_lookup0_cellmath__27[4]));
NAND2XL inst_lookup0_cellmath__29_0_I1823 (.Y(N12385), .A(N12381), .B(inst_lookup0_cellmath__27[4]));
NOR2XL inst_lookup0_cellmath__29_0_I1824 (.Y(N12404), .A(N1387), .B(N1388));
NOR2XL inst_lookup0_cellmath__29_0_I1825 (.Y(N12407), .A(inst_it2_lookup1_cellmath__53[0]), .B(inst_it2_lookup1_cellmath__53[1]));
NAND2XL inst_lookup0_cellmath__29_0_I1826 (.Y(N12401), .A(N12397), .B(N12407));
NOR2XL inst_lookup0_cellmath__29_0_I1827 (.Y(N12411), .A(inst_lookup0_cellmath__27[3]), .B(N12401));
AOI22XL inst_lookup0_cellmath__29_0_I1828 (.Y(N12408), .A0(N12397), .A1(N1388), .B0(N12407), .B1(inst_lookup0_cellmath__27[2]));
NAND2XL inst_lookup0_cellmath__29_0_I1829 (.Y(N12368), .A(inst_it2_lookup1_cellmath__53[1]), .B(inst_it2_lookup1_cellmath__53[0]));
AOI22XL inst_lookup0_cellmath__29_0_I1830 (.Y(N12376), .A0(N12397), .A1(N12368), .B0(N1388), .B1(inst_lookup0_cellmath__27[2]));
AOI22XL inst_lookup0_cellmath__29_0_I1831 (.Y(N12396), .A0(N12386), .A1(N12376), .B0(N12408), .B1(inst_lookup0_cellmath__27[3]));
NAND4BXL inst_lookup0_cellmath__29_0_I1832 (.Y(N12419), .AN(N12386), .B(inst_lookup0_cellmath__27[2]), .C(inst_lookup0_cellmath__27[4]), .D(N12404));
AOI22XL inst_lookup0_cellmath__29_0_I1833 (.Y(N12403), .A0(N12363), .A1(N12396), .B0(N12411), .B1(inst_lookup0_cellmath__27[4]));
INVXL inst_lookup0_cellmath__29_0_I1834 (.Y(N12409), .A(inst_lookup0_cellmath__27[5]));
AOI22XL inst_lookup0_cellmath__29_0_I1835 (.Y(N12362), .A0(N12409), .A1(N12419), .B0(N12394), .B1(inst_lookup0_cellmath__27[5]));
NOR2XL inst_lookup0_cellmath__29_0_I1836 (.Y(N12369), .A(inst_lookup0_cellmath__27[4]), .B(N12373));
NOR2XL inst_lookup0_cellmath__29_0_I1837 (.Y(N12380), .A(N12369), .B(N12409));
AOI22XL inst_lookup0_cellmath__29_0_I1838 (.Y(N12417), .A0(N12409), .A1(N12403), .B0(N12385), .B1(inst_lookup0_cellmath__27[5]));
NAND4BXL inst_lookup0_cellmath__29_0_I1839 (.Y(N12364), .AN(inst_lookup0_cellmath__27[3]), .B(N12404), .C(N12363), .D(N12397));
AOI22XL inst_lookup0_cellmath__29_0_I1840 (.Y(N12377), .A0(N1387), .A1(N1388), .B0(inst_it2_lookup1_cellmath__53[1]), .B1(inst_it2_lookup1_cellmath__53[0]));
AOI22XL inst_lookup0_cellmath__29_0_I1841 (.Y(N12395), .A0(N12397), .A1(N1388), .B0(N12377), .B1(inst_lookup0_cellmath__27[2]));
AOI22XL inst_lookup0_cellmath__29_0_I1842 (.Y(N12410), .A0(N12397), .A1(inst_it2_lookup1_cellmath__53[1]), .B0(N12404), .B1(inst_lookup0_cellmath__27[2]));
AOI22XL inst_lookup0_cellmath__29_0_I1843 (.Y(N12400), .A0(N12386), .A1(N12395), .B0(N1388), .B1(inst_lookup0_cellmath__27[3]));
NOR2XL inst_lookup0_cellmath__29_0_I1844 (.Y(N12414), .A(inst_lookup0_cellmath__27[3]), .B(N12410));
NAND2XL inst_lookup0_cellmath__29_0_I1845 (.Y(N12375), .A(N12407), .B(inst_lookup0_cellmath__27[2]));
NOR2XL inst_lookup0_cellmath__29_0_I1846 (.Y(N12405), .A(N12397), .B(N12379));
NOR2XL inst_lookup0_cellmath__29_0_I1847 (.Y(N12387), .A(N12397), .B(inst_it2_lookup1_cellmath__53[1]));
AOI22XL inst_lookup0_cellmath__29_0_I1848 (.Y(N12371), .A0(N12386), .A1(N12387), .B0(N12375), .B1(inst_lookup0_cellmath__27[3]));
NAND2XL inst_lookup0_cellmath__29_0_I1849 (.Y(N12384), .A(N12405), .B(inst_lookup0_cellmath__27[3]));
AOI22XL inst_lookup0_cellmath__29_0_I1850 (.Y(N12378), .A0(N12363), .A1(N12371), .B0(N12400), .B1(inst_lookup0_cellmath__27[4]));
AOI22XL inst_lookup0_cellmath__29_0_I1851 (.Y(N12392), .A0(N12363), .A1(N12384), .B0(N12414), .B1(inst_lookup0_cellmath__27[4]));
AOI22XL inst_lookup0_cellmath__29_0_I1852 (.Y(N12383), .A0(N12409), .A1(N12378), .B0(N12364), .B1(inst_lookup0_cellmath__27[5]));
NOR2XL inst_lookup0_cellmath__29_0_I1853 (.Y(N12399), .A(inst_lookup0_cellmath__27[5]), .B(N12392));
INVXL inst_lookup0_cellmath__29_0_I1854 (.Y(N12389), .A(inst_lookup0_cellmath__27[6]));
AOI22XL inst_lookup0_cellmath__29_0_I1855 (.Y(inst_cellmath__42[0]), .A0(inst_lookup0_cellmath__27[6]), .A1(N12362), .B0(N12389), .B1(N12383));
AOI22XL inst_lookup0_cellmath__29_0_I1856 (.Y(inst_lookup0_cellmath__29[1]), .A0(N12389), .A1(N12399), .B0(N12380), .B1(inst_lookup0_cellmath__27[6]));
NOR2XL inst_lookup0_cellmath__29_0_I1857 (.Y(inst_lookup0_cellmath__29[2]), .A(N12389), .B(N12417));
INVXL inst_cellmath__30__31__I1858 (.Y(inst_cellmath__43[0]), .A(inst_cellmath__42[0]));
INVXL inst_cellmath__30__31__I1859 (.Y(N2068), .A(inst_cellmath__43[0]));
AND2XL inst_cellmath__30__31__I1860 (.Y(N2045), .A(N2068), .B(inst_cellmath__9[0]));
AND2XL inst_cellmath__30__31__I1861 (.Y(N2046), .A(N2068), .B(inst_cellmath__9[1]));
AND2XL inst_cellmath__30__31__I1862 (.Y(N2047), .A(N2068), .B(inst_cellmath__9[2]));
AND2XL inst_cellmath__30__31__I1863 (.Y(N2048), .A(N2068), .B(inst_cellmath__9[3]));
AND2XL inst_cellmath__30__31__I1864 (.Y(N2049), .A(N2068), .B(inst_cellmath__9[4]));
AND2XL inst_cellmath__30__31__I1865 (.Y(N2050), .A(N2068), .B(inst_cellmath__9[5]));
AND2XL inst_cellmath__30__31__I1866 (.Y(N2051), .A(N2068), .B(inst_cellmath__9[6]));
AND2XL inst_cellmath__30__31__I1867 (.Y(N2052), .A(N2068), .B(inst_cellmath__9[7]));
AND2XL inst_cellmath__30__31__I1868 (.Y(N2053), .A(N2068), .B(inst_cellmath__9[8]));
AND2XL inst_cellmath__30__31__I1869 (.Y(N2054), .A(N2068), .B(inst_cellmath__9[9]));
AND2XL inst_cellmath__30__31__I1870 (.Y(N2055), .A(N2068), .B(inst_cellmath__9[10]));
AND2XL inst_cellmath__30__31__I1871 (.Y(N2056), .A(N2068), .B(inst_cellmath__9[11]));
AND2XL inst_cellmath__30__31__I1872 (.Y(N2057), .A(N2068), .B(inst_cellmath__9[12]));
AND2XL inst_cellmath__30__31__I1873 (.Y(N2058), .A(N2068), .B(inst_cellmath__9[13]));
AND2XL inst_cellmath__30__31__I1874 (.Y(N2059), .A(N2068), .B(inst_cellmath__9[14]));
AND2XL inst_cellmath__30__31__I1875 (.Y(N2060), .A(N2068), .B(inst_cellmath__9[15]));
AND2XL inst_cellmath__30__31__I1876 (.Y(N2061), .A(N2068), .B(inst_cellmath__9[16]));
AND2XL inst_cellmath__30__31__I1877 (.Y(N2062), .A(N2068), .B(inst_cellmath__9[17]));
AND2XL inst_cellmath__30__31__I1878 (.Y(N2063), .A(N2068), .B(inst_cellmath__9[18]));
AND2XL inst_cellmath__30__31__I1879 (.Y(N2064), .A(N2068), .B(inst_cellmath__9[19]));
AND2XL inst_cellmath__30__31__I1880 (.Y(N2065), .A(N2068), .B(inst_cellmath__9[20]));
AND2XL inst_cellmath__30__31__I1881 (.Y(N2066), .A(N2068), .B(inst_it2_lookup1_cellmath__53[0]));
AND2XL inst_cellmath__30__31__I1882 (.Y(N2067), .A(N2068), .B(inst_it2_lookup1_cellmath__53[1]));
INVXL inst_cellmath__31__35__I1883 (.Y(N12573), .A(inst_lookup0_cellmath__29[1]));
INVXL inst_cellmath__31__35__I1884 (.Y(N2173), .A(N12573));
NAND2XL inst_cellmath__31__35__I1885 (.Y(N2150), .A(N2173), .B(inst_cellmath__9[0]));
NAND2XL inst_cellmath__31__35__I1886 (.Y(N2151), .A(N2173), .B(inst_cellmath__9[1]));
NAND2XL inst_cellmath__31__35__I1887 (.Y(N2152), .A(N2173), .B(inst_cellmath__9[2]));
NAND2XL inst_cellmath__31__35__I1888 (.Y(N2153), .A(N2173), .B(inst_cellmath__9[3]));
NAND2XL inst_cellmath__31__35__I1889 (.Y(N2154), .A(N2173), .B(inst_cellmath__9[4]));
NAND2XL inst_cellmath__31__35__I1890 (.Y(N2155), .A(N2173), .B(inst_cellmath__9[5]));
NAND2XL inst_cellmath__31__35__I1891 (.Y(N2156), .A(N2173), .B(inst_cellmath__9[6]));
NAND2XL inst_cellmath__31__35__I1892 (.Y(N2157), .A(N2173), .B(inst_cellmath__9[7]));
NAND2XL inst_cellmath__31__35__I1893 (.Y(N2158), .A(N2173), .B(inst_cellmath__9[8]));
NAND2XL inst_cellmath__31__35__I1894 (.Y(N2159), .A(N2173), .B(inst_cellmath__9[9]));
NAND2XL inst_cellmath__31__35__I1895 (.Y(N2160), .A(N2173), .B(inst_cellmath__9[10]));
NAND2XL inst_cellmath__31__35__I1896 (.Y(N2161), .A(N2173), .B(inst_cellmath__9[11]));
NAND2XL inst_cellmath__31__35__I1897 (.Y(N2162), .A(N2173), .B(inst_cellmath__9[12]));
NAND2XL inst_cellmath__31__35__I1898 (.Y(N2163), .A(N2173), .B(inst_cellmath__9[13]));
NAND2XL inst_cellmath__31__35__I1899 (.Y(N2164), .A(N2173), .B(inst_cellmath__9[14]));
NAND2XL inst_cellmath__31__35__I1900 (.Y(N2165), .A(N2173), .B(inst_cellmath__9[15]));
NAND2XL inst_cellmath__31__35__I1901 (.Y(N2166), .A(N2173), .B(inst_cellmath__9[16]));
NAND2XL inst_cellmath__31__35__I1902 (.Y(N2167), .A(N2173), .B(inst_cellmath__9[17]));
NAND2XL inst_cellmath__31__35__I1903 (.Y(N2168), .A(N2173), .B(inst_cellmath__9[18]));
NAND2XL inst_cellmath__31__35__I1904 (.Y(N2169), .A(N2173), .B(inst_cellmath__9[19]));
NAND2XL inst_cellmath__31__35__I1905 (.Y(N2170), .A(N2173), .B(inst_cellmath__9[20]));
NAND2XL inst_cellmath__31__35__I1906 (.Y(N2171), .A(N2173), .B(inst_it2_lookup1_cellmath__53[0]));
NAND2XL inst_cellmath__31__35__I1907 (.Y(N2172), .A(N2173), .B(inst_it2_lookup1_cellmath__53[1]));
INVX1 inst_cellmath__20_0_I1908 (.Y(N12658), .A(inst_cellmath__11));
INVX1 inst_cellmath__20_0_I1909 (.Y(inst_cellmath__38__W0[2]), .A(N12658));
MX2XL inst_cellmath__20_0_I1911 (.Y(inst_cellmath__34[3]), .A(inst_cellmath__16[1]), .B(inst_cellmath__8[0]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1912 (.Y(inst_cellmath__34[4]), .A(inst_cellmath__16[2]), .B(inst_cellmath__8[1]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1913 (.Y(inst_cellmath__34[5]), .A(inst_cellmath__16[3]), .B(inst_cellmath__8[2]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1914 (.Y(inst_cellmath__34[6]), .A(inst_cellmath__16[4]), .B(inst_cellmath__8[3]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1915 (.Y(inst_cellmath__34[7]), .A(inst_cellmath__16[5]), .B(inst_cellmath__8[4]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1916 (.Y(inst_cellmath__34[8]), .A(inst_cellmath__16[6]), .B(inst_cellmath__8[5]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1917 (.Y(inst_cellmath__34[9]), .A(inst_cellmath__16[7]), .B(inst_cellmath__8[6]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1918 (.Y(inst_cellmath__34[10]), .A(inst_cellmath__16[8]), .B(inst_cellmath__8[7]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1919 (.Y(inst_cellmath__34[11]), .A(inst_cellmath__16[9]), .B(inst_cellmath__8[8]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1920 (.Y(inst_cellmath__34[12]), .A(inst_cellmath__16[10]), .B(inst_cellmath__8[9]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1921 (.Y(inst_cellmath__34[13]), .A(inst_cellmath__16[11]), .B(inst_cellmath__8[10]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1922 (.Y(inst_cellmath__34[14]), .A(inst_cellmath__16[12]), .B(inst_cellmath__8[11]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1923 (.Y(inst_cellmath__34[15]), .A(inst_cellmath__16[13]), .B(inst_cellmath__8[12]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1924 (.Y(inst_cellmath__34[16]), .A(inst_cellmath__16[14]), .B(inst_cellmath__8[13]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1925 (.Y(inst_cellmath__34[17]), .A(inst_cellmath__16[15]), .B(inst_cellmath__8[14]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1926 (.Y(inst_cellmath__34[18]), .A(inst_cellmath__16[16]), .B(inst_cellmath__8[15]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1927 (.Y(inst_cellmath__34[19]), .A(inst_cellmath__16[17]), .B(inst_cellmath__8[16]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1928 (.Y(inst_cellmath__34[20]), .A(inst_cellmath__16[18]), .B(inst_cellmath__8[17]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1929 (.Y(inst_cellmath__34[21]), .A(inst_cellmath__16[19]), .B(inst_cellmath__8[18]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1930 (.Y(inst_cellmath__34[22]), .A(inst_cellmath__16[20]), .B(inst_cellmath__8[19]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1931 (.Y(inst_cellmath__34[23]), .A(inst_cellmath__16[21]), .B(inst_cellmath__8[20]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1932 (.Y(inst_cellmath__34[24]), .A(inst_cellmath__16[22]), .B(inst_cellmath__8[21]), .S0(inst_cellmath__38__W0[2]));
MX2XL inst_cellmath__20_0_I1933 (.Y(inst_cellmath__34[25]), .A(inst_cellmath__16[23]), .B(inst_cellmath__8[22]), .S0(inst_cellmath__38__W0[2]));
INVXL cynw_cm_float_div_ieee_I158 (.Y(inst_it2_cellmath__60[4]), .A(inst_lookup0_cellmath__29[2]));
INVXL inst_cellmath__21_0_I1934 (.Y(N12797), .A(inst_cellmath__17[1]));
INVXL inst_cellmath__21_0_I1935 (.Y(N12723), .A(inst_cellmath__17[2]));
INVXL inst_cellmath__21_0_I1936 (.Y(N12744), .A(inst_cellmath__17[3]));
INVXL inst_cellmath__21_0_I1937 (.Y(N12764), .A(inst_cellmath__17[4]));
INVXL inst_cellmath__21_0_I1938 (.Y(N12785), .A(inst_cellmath__17[5]));
INVXL inst_cellmath__21_0_I1939 (.Y(N12806), .A(inst_cellmath__17[6]));
INVXL inst_cellmath__21_0_I1940 (.Y(N12732), .A(inst_cellmath__17[7]));
INVXL inst_cellmath__21_0_I1941 (.Y(N12754), .A(inst_cellmath__17[8]));
INVXL inst_cellmath__21_0_I1942 (.Y(N12774), .A(inst_cellmath__17[9]));
INVXL inst_cellmath__21_0_I1943 (.Y(N12794), .A(inst_cellmath__17[10]));
INVXL inst_cellmath__21_0_I1944 (.Y(N12720), .A(inst_cellmath__17[11]));
INVXL inst_cellmath__21_0_I1945 (.Y(N12740), .A(inst_cellmath__17[12]));
INVXL inst_cellmath__21_0_I1946 (.Y(N12761), .A(inst_cellmath__17[13]));
INVXL inst_cellmath__21_0_I1947 (.Y(N12782), .A(inst_cellmath__17[14]));
INVXL inst_cellmath__21_0_I1948 (.Y(N12803), .A(inst_cellmath__17[15]));
INVXL inst_cellmath__21_0_I1949 (.Y(N12729), .A(inst_cellmath__17[16]));
INVXL inst_cellmath__21_0_I1950 (.Y(N12751), .A(inst_cellmath__17[17]));
INVXL inst_cellmath__21_0_I1951 (.Y(N12771), .A(inst_cellmath__17[18]));
INVXL inst_cellmath__21_0_I1952 (.Y(N12791), .A(inst_cellmath__17[19]));
INVXL inst_cellmath__21_0_I1953 (.Y(N12813), .A(inst_cellmath__17[20]));
INVXL inst_cellmath__21_0_I1954 (.Y(N12738), .A(inst_cellmath__17[21]));
AOI22XL inst_cellmath__21_0_I1957 (.Y(inst_cellmath__35[3]), .A0(N12658), .A1(N12797), .B0(inst_cellmath__9[0]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1958 (.Y(inst_cellmath__35[4]), .A0(N12658), .A1(N12723), .B0(inst_cellmath__9[1]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1959 (.Y(inst_cellmath__35[5]), .A0(N12658), .A1(N12744), .B0(inst_cellmath__9[2]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1960 (.Y(inst_cellmath__35[6]), .A0(N12658), .A1(N12764), .B0(inst_cellmath__9[3]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1961 (.Y(inst_cellmath__35[7]), .A0(N12658), .A1(N12785), .B0(inst_cellmath__9[4]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1962 (.Y(inst_cellmath__35[8]), .A0(N12658), .A1(N12806), .B0(inst_cellmath__9[5]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1963 (.Y(inst_cellmath__35[9]), .A0(N12658), .A1(N12732), .B0(inst_cellmath__9[6]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1964 (.Y(inst_cellmath__35[10]), .A0(N12658), .A1(N12754), .B0(inst_cellmath__9[7]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1965 (.Y(inst_cellmath__35[11]), .A0(N12658), .A1(N12774), .B0(inst_cellmath__9[8]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1966 (.Y(inst_cellmath__35[12]), .A0(N12658), .A1(N12794), .B0(inst_cellmath__9[9]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1967 (.Y(inst_cellmath__35[13]), .A0(N12658), .A1(N12720), .B0(inst_cellmath__9[10]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1968 (.Y(inst_cellmath__35[14]), .A0(N12658), .A1(N12740), .B0(inst_cellmath__9[11]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1969 (.Y(inst_cellmath__35[15]), .A0(N12658), .A1(N12761), .B0(inst_cellmath__9[12]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1970 (.Y(inst_cellmath__35[16]), .A0(N12658), .A1(N12782), .B0(inst_cellmath__9[13]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1971 (.Y(inst_cellmath__35[17]), .A0(N12658), .A1(N12803), .B0(inst_cellmath__9[14]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1972 (.Y(inst_cellmath__35[18]), .A0(N12658), .A1(N12729), .B0(inst_cellmath__9[15]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1973 (.Y(inst_cellmath__35[19]), .A0(N12658), .A1(N12751), .B0(inst_cellmath__9[16]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1974 (.Y(inst_cellmath__35[20]), .A0(N12658), .A1(N12771), .B0(inst_cellmath__9[17]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1975 (.Y(inst_cellmath__35[21]), .A0(N12658), .A1(N12791), .B0(inst_cellmath__9[18]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1976 (.Y(inst_cellmath__35[22]), .A0(N12658), .A1(N12813), .B0(inst_cellmath__9[19]), .B1(inst_cellmath__11));
AOI22XL inst_cellmath__21_0_I1977 (.Y(inst_cellmath__35[23]), .A0(N12658), .A1(N12738), .B0(inst_cellmath__9[20]), .B1(inst_cellmath__11));
INVXL inst_cellmath__21_0_I1978 (.Y(N12811), .A(inst_cellmath__17[22]));
AOI22XL inst_cellmath__21_0_I1979 (.Y(inst_cellmath__35[24]), .A0(N12658), .A1(N12811), .B0(inst_it2_lookup1_cellmath__53[0]), .B1(inst_cellmath__11));
INVXL inst_cellmath__21_0_I1980 (.Y(N12736), .A(inst_cellmath__17[23]));
AOI22XL inst_cellmath__21_0_I1981 (.Y(inst_cellmath__35[25]), .A0(N12658), .A1(N12736), .B0(inst_it2_lookup1_cellmath__53[1]), .B1(inst_cellmath__11));
INVX1 cynw_cm_float_div_ieee_I1983 (.Y(N12870), .A(inst_it2_cellmath__60[4]));
XNOR2X1 cynw_cm_float_div_ieee_I1984 (.Y(inst_it2_cellmath__61[3]), .A(N2045), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1985 (.Y(inst_cellmath__38__W1[2]), .A(N2046), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1986 (.Y(inst_cellmath__30[3]), .A(N2047), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1987 (.Y(inst_cellmath__30[4]), .A(N2048), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1988 (.Y(inst_cellmath__30[5]), .A(N2049), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1989 (.Y(inst_cellmath__30[6]), .A(N2050), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1990 (.Y(inst_cellmath__30[7]), .A(N2051), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1991 (.Y(inst_cellmath__30[8]), .A(N2052), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1992 (.Y(inst_cellmath__30[9]), .A(N2053), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1993 (.Y(inst_cellmath__30[10]), .A(N2054), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1994 (.Y(inst_cellmath__30[11]), .A(N2055), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1995 (.Y(inst_cellmath__30[12]), .A(N2056), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1996 (.Y(inst_cellmath__30[13]), .A(N2057), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1997 (.Y(inst_cellmath__30[14]), .A(N2058), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1998 (.Y(inst_cellmath__30[15]), .A(N2059), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I1999 (.Y(inst_cellmath__30[16]), .A(N2060), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2000 (.Y(inst_cellmath__30[17]), .A(N2061), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2001 (.Y(inst_cellmath__30[18]), .A(N2062), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2002 (.Y(inst_cellmath__30[19]), .A(N2063), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2003 (.Y(inst_cellmath__30[20]), .A(N2064), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2004 (.Y(inst_cellmath__30[21]), .A(N2065), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2005 (.Y(inst_cellmath__30[22]), .A(N2066), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2006 (.Y(inst_cellmath__30[23]), .A(N2067), .B(N12870));
XNOR2X1 cynw_cm_float_div_ieee_I2007 (.Y(inst_cellmath__30[24]), .A(N2068), .B(N12870));
ADDFX1 inst_fa_1033_10_I2009 (.CO(inst_cellmath__38__W0[3]), .S(inst_cellmath__38__W1[3]), .A(inst_cellmath__35[3]), .B(inst_cellmath__34[3]), .CI(inst_cellmath__30[3]));
ADDFX1 inst_fa_1033_10_I2010 (.CO(inst_cellmath__38__W0[4]), .S(inst_cellmath__38__W1[4]), .A(inst_cellmath__35[4]), .B(inst_cellmath__34[4]), .CI(inst_cellmath__30[4]));
ADDFX1 inst_fa_1033_10_I2011 (.CO(inst_cellmath__38__W0[5]), .S(inst_cellmath__38__W1[5]), .A(inst_cellmath__35[5]), .B(inst_cellmath__34[5]), .CI(inst_cellmath__30[5]));
ADDFX1 inst_fa_1033_10_I2012 (.CO(inst_cellmath__38__W0[6]), .S(inst_cellmath__38__W1[6]), .A(inst_cellmath__35[6]), .B(inst_cellmath__34[6]), .CI(inst_cellmath__30[6]));
ADDFX1 inst_fa_1033_10_I2013 (.CO(inst_cellmath__38__W0[7]), .S(inst_cellmath__38__W1[7]), .A(inst_cellmath__35[7]), .B(inst_cellmath__34[7]), .CI(inst_cellmath__30[7]));
ADDFX1 inst_fa_1033_10_I2014 (.CO(inst_cellmath__38__W0[8]), .S(inst_cellmath__38__W1[8]), .A(inst_cellmath__35[8]), .B(inst_cellmath__34[8]), .CI(inst_cellmath__30[8]));
ADDFX1 inst_fa_1033_10_I2015 (.CO(inst_cellmath__38__W0[9]), .S(inst_cellmath__38__W1[9]), .A(inst_cellmath__35[9]), .B(inst_cellmath__34[9]), .CI(inst_cellmath__30[9]));
ADDFX1 inst_fa_1033_10_I2016 (.CO(inst_cellmath__38__W0[10]), .S(inst_cellmath__38__W1[10]), .A(inst_cellmath__35[10]), .B(inst_cellmath__34[10]), .CI(inst_cellmath__30[10]));
ADDFX1 inst_fa_1033_10_I2017 (.CO(inst_cellmath__38__W0[11]), .S(inst_cellmath__38__W1[11]), .A(inst_cellmath__35[11]), .B(inst_cellmath__34[11]), .CI(inst_cellmath__30[11]));
ADDFX1 inst_fa_1033_10_I2018 (.CO(inst_cellmath__38__W0[12]), .S(inst_cellmath__38__W1[12]), .A(inst_cellmath__35[12]), .B(inst_cellmath__34[12]), .CI(inst_cellmath__30[12]));
ADDFX1 inst_fa_1033_10_I2019 (.CO(inst_cellmath__38__W0[13]), .S(inst_cellmath__38__W1[13]), .A(inst_cellmath__35[13]), .B(inst_cellmath__34[13]), .CI(inst_cellmath__30[13]));
ADDFX1 inst_fa_1033_10_I2020 (.CO(inst_cellmath__38__W0[14]), .S(inst_cellmath__38__W1[14]), .A(inst_cellmath__35[14]), .B(inst_cellmath__34[14]), .CI(inst_cellmath__30[14]));
ADDFX1 inst_fa_1033_10_I2021 (.CO(inst_cellmath__38__W0[15]), .S(inst_cellmath__38__W1[15]), .A(inst_cellmath__35[15]), .B(inst_cellmath__34[15]), .CI(inst_cellmath__30[15]));
ADDFX1 inst_fa_1033_10_I2022 (.CO(inst_cellmath__38__W0[16]), .S(inst_cellmath__38__W1[16]), .A(inst_cellmath__35[16]), .B(inst_cellmath__34[16]), .CI(inst_cellmath__30[16]));
ADDFX1 inst_fa_1033_10_I2023 (.CO(inst_cellmath__38__W0[17]), .S(inst_cellmath__38__W1[17]), .A(inst_cellmath__35[17]), .B(inst_cellmath__34[17]), .CI(inst_cellmath__30[17]));
ADDFX1 inst_fa_1033_10_I2024 (.CO(inst_cellmath__38__W0[18]), .S(inst_cellmath__38__W1[18]), .A(inst_cellmath__35[18]), .B(inst_cellmath__34[18]), .CI(inst_cellmath__30[18]));
ADDFX1 inst_fa_1033_10_I2025 (.CO(inst_cellmath__38__W0[19]), .S(inst_cellmath__38__W1[19]), .A(inst_cellmath__35[19]), .B(inst_cellmath__34[19]), .CI(inst_cellmath__30[19]));
ADDFX1 inst_fa_1033_10_I2026 (.CO(inst_cellmath__38__W0[20]), .S(inst_cellmath__38__W1[20]), .A(inst_cellmath__35[20]), .B(inst_cellmath__34[20]), .CI(inst_cellmath__30[20]));
ADDFX1 inst_fa_1033_10_I2027 (.CO(inst_cellmath__38__W0[21]), .S(inst_cellmath__38__W1[21]), .A(inst_cellmath__35[21]), .B(inst_cellmath__34[21]), .CI(inst_cellmath__30[21]));
ADDFX1 inst_fa_1033_10_I2028 (.CO(inst_cellmath__38__W0[22]), .S(inst_cellmath__38__W1[22]), .A(inst_cellmath__35[22]), .B(inst_cellmath__34[22]), .CI(inst_cellmath__30[22]));
ADDFX1 inst_fa_1033_10_I2029 (.CO(inst_cellmath__38__W0[23]), .S(inst_cellmath__38__W1[23]), .A(inst_cellmath__35[23]), .B(inst_cellmath__34[23]), .CI(inst_cellmath__30[23]));
ADDFX1 inst_fa_1033_10_I2030 (.CO(inst_cellmath__38__W0[24]), .S(inst_cellmath__38__W1[24]), .A(inst_cellmath__35[24]), .B(inst_cellmath__34[24]), .CI(inst_cellmath__30[24]));
ADDFX1 inst_fa_1033_10_I2031 (.CO(N12983), .S(inst_cellmath__38__W1[25]), .A(inst_cellmath__35[25]), .B(inst_cellmath__34[25]), .CI(inst_it2_cellmath__60[4]));
INVXL cynw_cm_float_div_ieee_I2034 (.Y(inst_cellmath__31[1]), .A(N12870));
MXI2XL cynw_cm_float_div_ieee_I2035 (.Y(inst_cellmath__31[2]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2150));
MXI2XL cynw_cm_float_div_ieee_I2036 (.Y(inst_cellmath__31[3]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2151));
MXI2XL cynw_cm_float_div_ieee_I2037 (.Y(inst_cellmath__31[4]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2152));
MXI2XL cynw_cm_float_div_ieee_I2038 (.Y(inst_cellmath__31[5]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2153));
MXI2XL cynw_cm_float_div_ieee_I2039 (.Y(inst_cellmath__31[6]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2154));
MXI2XL cynw_cm_float_div_ieee_I2040 (.Y(inst_cellmath__31[7]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2155));
MXI2XL cynw_cm_float_div_ieee_I2041 (.Y(inst_cellmath__31[8]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2156));
MXI2XL cynw_cm_float_div_ieee_I2042 (.Y(inst_cellmath__31[9]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2157));
MXI2XL cynw_cm_float_div_ieee_I2043 (.Y(inst_cellmath__31[10]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2158));
MXI2XL cynw_cm_float_div_ieee_I2044 (.Y(inst_cellmath__31[11]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2159));
MXI2XL cynw_cm_float_div_ieee_I2045 (.Y(inst_cellmath__31[12]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2160));
MXI2XL cynw_cm_float_div_ieee_I2046 (.Y(inst_cellmath__31[13]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2161));
MXI2XL cynw_cm_float_div_ieee_I2047 (.Y(inst_cellmath__31[14]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2162));
MXI2XL cynw_cm_float_div_ieee_I2048 (.Y(inst_cellmath__31[15]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2163));
MXI2XL cynw_cm_float_div_ieee_I2049 (.Y(inst_cellmath__31[16]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2164));
MXI2XL cynw_cm_float_div_ieee_I2050 (.Y(inst_cellmath__31[17]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2165));
MXI2XL cynw_cm_float_div_ieee_I2051 (.Y(inst_cellmath__31[18]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2166));
MXI2XL cynw_cm_float_div_ieee_I2052 (.Y(inst_cellmath__31[19]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2167));
MXI2XL cynw_cm_float_div_ieee_I2053 (.Y(inst_cellmath__31[20]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2168));
MXI2XL cynw_cm_float_div_ieee_I2054 (.Y(inst_cellmath__31[21]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2169));
MXI2XL cynw_cm_float_div_ieee_I2055 (.Y(inst_cellmath__31[22]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2170));
MXI2XL cynw_cm_float_div_ieee_I2056 (.Y(inst_cellmath__31[23]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2171));
MXI2XL cynw_cm_float_div_ieee_I2057 (.Y(inst_cellmath__31[24]), .A(inst_cellmath__31[1]), .B(N12870), .S0(N2172));
MXI2XL cynw_cm_float_div_ieee_I2058 (.Y(inst_cellmath__31[25]), .A(N12870), .B(inst_cellmath__31[1]), .S0(N2173));
INVXL buf1_A_I9199 (.Y(N28016), .A(inst_it2_cellmath__60[4]));
INVXL buf1_A_I9200 (.Y(inst_it2_cellmath__60[3]), .A(N28016));
ADDHX1 inst_fa_1052_10_I2061 (.CO(inst_it2_cellmath__60[5]), .S(inst_it2_cellmath__61[4]), .A(inst_cellmath__38__W1[2]), .B(inst_cellmath__31[2]));
ADDFX1 inst_fa_1052_10_I2062 (.CO(inst_it2_cellmath__60[6]), .S(inst_it2_cellmath__61[5]), .A(inst_cellmath__38__W0[2]), .B(inst_cellmath__38__W1[3]), .CI(inst_cellmath__31[3]));
ADDFX1 inst_fa_1052_10_I2063 (.CO(inst_it2_cellmath__60[7]), .S(inst_it2_cellmath__61[6]), .A(inst_cellmath__38__W0[3]), .B(inst_cellmath__38__W1[4]), .CI(inst_cellmath__31[4]));
ADDFX1 inst_fa_1052_10_I2064 (.CO(inst_it2_cellmath__60[8]), .S(inst_it2_cellmath__61[7]), .A(inst_cellmath__38__W0[4]), .B(inst_cellmath__38__W1[5]), .CI(inst_cellmath__31[5]));
ADDFX1 inst_fa_1052_10_I2065 (.CO(inst_it2_cellmath__60[9]), .S(inst_it2_cellmath__61[8]), .A(inst_cellmath__38__W0[5]), .B(inst_cellmath__38__W1[6]), .CI(inst_cellmath__31[6]));
ADDFX1 inst_fa_1052_10_I2066 (.CO(inst_it2_cellmath__60[10]), .S(inst_it2_cellmath__61[9]), .A(inst_cellmath__38__W0[6]), .B(inst_cellmath__38__W1[7]), .CI(inst_cellmath__31[7]));
ADDFX1 inst_fa_1052_10_I2067 (.CO(inst_it2_cellmath__60[11]), .S(inst_it2_cellmath__61[10]), .A(inst_cellmath__38__W0[7]), .B(inst_cellmath__38__W1[8]), .CI(inst_cellmath__31[8]));
ADDFX1 inst_fa_1052_10_I2068 (.CO(inst_it2_cellmath__60[12]), .S(inst_it2_cellmath__61[11]), .A(inst_cellmath__38__W0[8]), .B(inst_cellmath__38__W1[9]), .CI(inst_cellmath__31[9]));
ADDFX1 inst_fa_1052_10_I2069 (.CO(inst_it2_cellmath__60[13]), .S(inst_it2_cellmath__61[12]), .A(inst_cellmath__38__W0[9]), .B(inst_cellmath__38__W1[10]), .CI(inst_cellmath__31[10]));
ADDFX1 inst_fa_1052_10_I2070 (.CO(inst_it2_cellmath__60[14]), .S(inst_it2_cellmath__61[13]), .A(inst_cellmath__38__W0[10]), .B(inst_cellmath__38__W1[11]), .CI(inst_cellmath__31[11]));
ADDFX1 inst_fa_1052_10_I2071 (.CO(inst_it2_cellmath__60[15]), .S(inst_it2_cellmath__61[14]), .A(inst_cellmath__38__W0[11]), .B(inst_cellmath__38__W1[12]), .CI(inst_cellmath__31[12]));
ADDFX1 inst_fa_1052_10_I2072 (.CO(inst_it2_cellmath__60[16]), .S(inst_it2_cellmath__61[15]), .A(inst_cellmath__38__W0[12]), .B(inst_cellmath__38__W1[13]), .CI(inst_cellmath__31[13]));
ADDFX1 inst_fa_1052_10_I2073 (.CO(inst_it2_cellmath__60[17]), .S(inst_it2_cellmath__61[16]), .A(inst_cellmath__38__W0[13]), .B(inst_cellmath__38__W1[14]), .CI(inst_cellmath__31[14]));
ADDFX1 inst_fa_1052_10_I2074 (.CO(inst_it2_cellmath__60[18]), .S(inst_it2_cellmath__61[17]), .A(inst_cellmath__38__W0[14]), .B(inst_cellmath__38__W1[15]), .CI(inst_cellmath__31[15]));
ADDFX1 inst_fa_1052_10_I2075 (.CO(inst_it2_cellmath__60[19]), .S(inst_it2_cellmath__61[18]), .A(inst_cellmath__38__W0[15]), .B(inst_cellmath__38__W1[16]), .CI(inst_cellmath__31[16]));
ADDFX1 inst_fa_1052_10_I2076 (.CO(inst_it2_cellmath__60[20]), .S(inst_it2_cellmath__61[19]), .A(inst_cellmath__38__W0[16]), .B(inst_cellmath__38__W1[17]), .CI(inst_cellmath__31[17]));
ADDFX1 inst_fa_1052_10_I2077 (.CO(inst_it2_cellmath__60[21]), .S(inst_it2_cellmath__61[20]), .A(inst_cellmath__38__W0[17]), .B(inst_cellmath__38__W1[18]), .CI(inst_cellmath__31[18]));
ADDFX1 inst_fa_1052_10_I2078 (.CO(inst_it2_cellmath__60[22]), .S(inst_it2_cellmath__61[21]), .A(inst_cellmath__38__W0[18]), .B(inst_cellmath__38__W1[19]), .CI(inst_cellmath__31[19]));
ADDFX1 inst_fa_1052_10_I2079 (.CO(inst_it2_cellmath__60[23]), .S(inst_it2_cellmath__61[22]), .A(inst_cellmath__38__W0[19]), .B(inst_cellmath__38__W1[20]), .CI(inst_cellmath__31[20]));
ADDFX1 inst_fa_1052_10_I2080 (.CO(inst_it2_cellmath__60[24]), .S(inst_it2_cellmath__61[23]), .A(inst_cellmath__38__W0[20]), .B(inst_cellmath__38__W1[21]), .CI(inst_cellmath__31[21]));
ADDFX1 inst_fa_1052_10_I2081 (.CO(inst_it2_cellmath__60[25]), .S(inst_it2_cellmath__61[24]), .A(inst_cellmath__38__W0[21]), .B(inst_cellmath__38__W1[22]), .CI(inst_cellmath__31[22]));
ADDFX1 inst_fa_1052_10_I2082 (.CO(inst_cellmath__39__W0[23]), .S(inst_it2_cellmath__61[25]), .A(inst_cellmath__38__W0[22]), .B(inst_cellmath__38__W1[23]), .CI(inst_cellmath__31[23]));
ADDFX1 inst_fa_1052_10_I2083 (.CO(inst_cellmath__39__W0[24]), .S(inst_cellmath__39__W1[24]), .A(inst_cellmath__38__W0[23]), .B(inst_cellmath__38__W1[24]), .CI(inst_cellmath__31[24]));
ADDFX1 inst_fa_1052_10_I2084 (.CO(N13206), .S(inst_cellmath__39__W1[25]), .A(inst_cellmath__38__W0[24]), .B(inst_cellmath__38__W1[25]), .CI(inst_cellmath__31[25]));
ADDHX1 inst_it2_cellmath__51_0_I2085 (.CO(N13380), .S(inst_it2_lookup1_cellmath__53[2]), .A(inst_it2_cellmath__60[23]), .B(inst_it2_cellmath__61[23]));
ADDFX1 inst_it2_cellmath__51_0_I2086 (.CO(N13376), .S(inst_it2_lookup1_cellmath__53[3]), .A(inst_it2_cellmath__61[24]), .B(inst_it2_cellmath__60[24]), .CI(N13380));
ADDFX1 inst_it2_cellmath__51_0_I2087 (.CO(N13387), .S(inst_it2_lookup1_cellmath__53[4]), .A(inst_it2_cellmath__61[25]), .B(inst_it2_cellmath__60[25]), .CI(N13376));
ADDFX1 inst_it2_cellmath__51_0_I2088 (.CO(N13373), .S(inst_it2_lookup1_cellmath__53[5]), .A(inst_cellmath__39__W1[24]), .B(inst_cellmath__39__W0[23]), .CI(N13387));
ADDFX1 inst_it2_cellmath__51_0_I2089 (.CO(N13384), .S(inst_it2_lookup1_cellmath__53[6]), .A(inst_cellmath__39__W0[24]), .B(inst_cellmath__39__W1[25]), .CI(N13373));
INVXL inst_it2_lookup1_cellmath__55_0_I2092 (.Y(N13436), .A(inst_it2_lookup1_cellmath__53[2]));
INVXL inst_it2_lookup1_cellmath__55_0_I2093 (.Y(N13425), .A(inst_it2_lookup1_cellmath__53[3]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2094 (.Y(N13420), .A(N13425), .B(N13436));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2095 (.Y(N13457), .A(N13436), .B(N1388));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2097 (.Y(N13405), .A0(N13436), .A1(inst_it2_lookup1_cellmath__53[1]), .B0(N12379), .B1(inst_it2_lookup1_cellmath__53[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2098 (.Y(N13460), .A0(N13425), .A1(N13405), .B0(N13457), .B1(inst_it2_lookup1_cellmath__53[3]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I2099 (.Y(N13404), .A(inst_it2_lookup1_cellmath__53[1]), .B(inst_it2_lookup1_cellmath__53[2]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2100 (.Y(N13412), .A(N13425), .B(N13404));
INVXL inst_it2_lookup1_cellmath__55_0_I2101 (.Y(N13402), .A(inst_it2_lookup1_cellmath__53[4]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2102 (.Y(N13433), .A0(N13402), .A1(N13460), .B0(N13420), .B1(inst_it2_lookup1_cellmath__53[4]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I2103 (.Y(N13424), .A(N13420), .B(inst_it2_lookup1_cellmath__53[4]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I2106 (.Y(N13440), .A(N13436), .B(N12407));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2107 (.Y(N13450), .A(inst_it2_lookup1_cellmath__53[3]), .B(N13440));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2108 (.Y(N13447), .A0(N13436), .A1(N1388), .B0(N12407), .B1(inst_it2_lookup1_cellmath__53[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2110 (.Y(N13415), .A0(N13436), .A1(N12368), .B0(N1388), .B1(inst_it2_lookup1_cellmath__53[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2111 (.Y(N13435), .A0(N13425), .A1(N13415), .B0(N13447), .B1(inst_it2_lookup1_cellmath__53[3]));
NAND4BXL inst_it2_lookup1_cellmath__55_0_I2112 (.Y(N13458), .AN(N13425), .B(N12404), .C(inst_it2_lookup1_cellmath__53[4]), .D(inst_it2_lookup1_cellmath__53[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2113 (.Y(N13442), .A0(N13402), .A1(N13435), .B0(N13450), .B1(inst_it2_lookup1_cellmath__53[4]));
INVXL inst_it2_lookup1_cellmath__55_0_I2114 (.Y(N13448), .A(inst_it2_lookup1_cellmath__53[5]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2115 (.Y(N13401), .A0(N13448), .A1(N13458), .B0(N13433), .B1(inst_it2_lookup1_cellmath__53[5]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2116 (.Y(N13408), .A(inst_it2_lookup1_cellmath__53[4]), .B(N13412));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2117 (.Y(N13419), .A(N13408), .B(N13448));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2118 (.Y(N13456), .A0(N13448), .A1(N13442), .B0(N13424), .B1(inst_it2_lookup1_cellmath__53[5]));
NAND4BXL inst_it2_lookup1_cellmath__55_0_I2119 (.Y(N13403), .AN(inst_it2_lookup1_cellmath__53[3]), .B(N12404), .C(N13402), .D(N13436));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2121 (.Y(N13434), .A0(N13436), .A1(N1388), .B0(N12377), .B1(inst_it2_lookup1_cellmath__53[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2122 (.Y(N13449), .A0(N13436), .A1(inst_it2_lookup1_cellmath__53[1]), .B0(N12404), .B1(inst_it2_lookup1_cellmath__53[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2123 (.Y(N13439), .A0(N13425), .A1(N13434), .B0(N1388), .B1(inst_it2_lookup1_cellmath__53[3]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2124 (.Y(N13453), .A(inst_it2_lookup1_cellmath__53[3]), .B(N13449));
NAND2XL inst_it2_lookup1_cellmath__55_0_I2125 (.Y(N13414), .A(N12407), .B(inst_it2_lookup1_cellmath__53[2]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2126 (.Y(N13444), .A(N13436), .B(N12379));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2127 (.Y(N13426), .A(N13436), .B(inst_it2_lookup1_cellmath__53[1]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2128 (.Y(N13410), .A0(N13425), .A1(N13426), .B0(N13414), .B1(inst_it2_lookup1_cellmath__53[3]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I2129 (.Y(N13423), .A(N13444), .B(inst_it2_lookup1_cellmath__53[3]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2130 (.Y(N13417), .A0(N13402), .A1(N13410), .B0(N13439), .B1(inst_it2_lookup1_cellmath__53[4]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2131 (.Y(N13431), .A0(N13402), .A1(N13423), .B0(N13453), .B1(inst_it2_lookup1_cellmath__53[4]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2132 (.Y(N13422), .A0(N13448), .A1(N13417), .B0(N13403), .B1(inst_it2_lookup1_cellmath__53[5]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2133 (.Y(N13438), .A(inst_it2_lookup1_cellmath__53[5]), .B(N13431));
INVXL inst_it2_lookup1_cellmath__55_0_I2134 (.Y(N13428), .A(inst_it2_lookup1_cellmath__53[6]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2135 (.Y(inst_cellmath__40[0]), .A0(inst_it2_lookup1_cellmath__53[6]), .A1(N13401), .B0(N13428), .B1(N13422));
AOI22XL inst_it2_lookup1_cellmath__55_0_I2136 (.Y(inst_it2_lookup1_cellmath__55[1]), .A0(N13428), .A1(N13438), .B0(N13419), .B1(inst_it2_lookup1_cellmath__53[6]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I2137 (.Y(inst_it2_lookup1_cellmath__55[2]), .A(N13428), .B(N13456));
INVXL inst_it2_cellmath__56__57__I2138 (.Y(inst_cellmath__41[0]), .A(inst_cellmath__40[0]));
INVXL inst_it2_cellmath__56__57__I2139 (.Y(N2224), .A(inst_cellmath__41[0]));
AND2XL inst_it2_cellmath__56__57__I2140 (.Y(N2201), .A(N2224), .B(inst_cellmath__9[0]));
AND2XL inst_it2_cellmath__56__57__I2141 (.Y(N2202), .A(N2224), .B(inst_cellmath__9[1]));
AND2XL inst_it2_cellmath__56__57__I2142 (.Y(N2203), .A(N2224), .B(inst_cellmath__9[2]));
AND2XL inst_it2_cellmath__56__57__I2143 (.Y(N2204), .A(N2224), .B(inst_cellmath__9[3]));
AND2XL inst_it2_cellmath__56__57__I2144 (.Y(N2205), .A(N2224), .B(inst_cellmath__9[4]));
AND2XL inst_it2_cellmath__56__57__I2145 (.Y(N2206), .A(N2224), .B(inst_cellmath__9[5]));
AND2XL inst_it2_cellmath__56__57__I2146 (.Y(N2207), .A(N2224), .B(inst_cellmath__9[6]));
AND2XL inst_it2_cellmath__56__57__I2147 (.Y(N2208), .A(N2224), .B(inst_cellmath__9[7]));
AND2XL inst_it2_cellmath__56__57__I2148 (.Y(N2209), .A(N2224), .B(inst_cellmath__9[8]));
AND2XL inst_it2_cellmath__56__57__I2149 (.Y(N2210), .A(N2224), .B(inst_cellmath__9[9]));
AND2XL inst_it2_cellmath__56__57__I2150 (.Y(N2211), .A(N2224), .B(inst_cellmath__9[10]));
AND2XL inst_it2_cellmath__56__57__I2151 (.Y(N2212), .A(N2224), .B(inst_cellmath__9[11]));
AND2XL inst_it2_cellmath__56__57__I2152 (.Y(N2213), .A(N2224), .B(inst_cellmath__9[12]));
AND2XL inst_it2_cellmath__56__57__I2153 (.Y(N2214), .A(N2224), .B(inst_cellmath__9[13]));
AND2XL inst_it2_cellmath__56__57__I2154 (.Y(N2215), .A(N2224), .B(inst_cellmath__9[14]));
AND2XL inst_it2_cellmath__56__57__I2155 (.Y(N2216), .A(N2224), .B(inst_cellmath__9[15]));
AND2XL inst_it2_cellmath__56__57__I2156 (.Y(N2217), .A(N2224), .B(inst_cellmath__9[16]));
AND2XL inst_it2_cellmath__56__57__I2157 (.Y(N2218), .A(N2224), .B(inst_cellmath__9[17]));
AND2XL inst_it2_cellmath__56__57__I2158 (.Y(N2219), .A(N2224), .B(inst_cellmath__9[18]));
AND2XL inst_it2_cellmath__56__57__I2159 (.Y(N2220), .A(N2224), .B(inst_cellmath__9[19]));
AND2XL inst_it2_cellmath__56__57__I2160 (.Y(N2221), .A(N2224), .B(inst_cellmath__9[20]));
AND2XL inst_it2_cellmath__56__57__I2161 (.Y(N2222), .A(N2224), .B(inst_it2_lookup1_cellmath__53[0]));
AND2XL inst_it2_cellmath__56__57__I2162 (.Y(N2223), .A(N2224), .B(inst_it2_lookup1_cellmath__53[1]));
INVXL inst_it2_cellmath__57__61__I2163 (.Y(N13614), .A(inst_it2_lookup1_cellmath__55[1]));
INVXL inst_it2_cellmath__57__61__I2164 (.Y(N2277), .A(N13614));
NAND2XL inst_it2_cellmath__57__61__I2165 (.Y(N2254), .A(N2277), .B(inst_cellmath__9[0]));
NAND2XL inst_it2_cellmath__57__61__I2166 (.Y(N2255), .A(N2277), .B(inst_cellmath__9[1]));
NAND2XL inst_it2_cellmath__57__61__I2167 (.Y(N2256), .A(N2277), .B(inst_cellmath__9[2]));
NAND2XL inst_it2_cellmath__57__61__I2168 (.Y(N2257), .A(N2277), .B(inst_cellmath__9[3]));
NAND2XL inst_it2_cellmath__57__61__I2169 (.Y(N2258), .A(N2277), .B(inst_cellmath__9[4]));
NAND2XL inst_it2_cellmath__57__61__I2170 (.Y(N2259), .A(N2277), .B(inst_cellmath__9[5]));
NAND2XL inst_it2_cellmath__57__61__I2171 (.Y(N2260), .A(N2277), .B(inst_cellmath__9[6]));
NAND2XL inst_it2_cellmath__57__61__I2172 (.Y(N2261), .A(N2277), .B(inst_cellmath__9[7]));
NAND2XL inst_it2_cellmath__57__61__I2173 (.Y(N2262), .A(N2277), .B(inst_cellmath__9[8]));
NAND2XL inst_it2_cellmath__57__61__I2174 (.Y(N2263), .A(N2277), .B(inst_cellmath__9[9]));
NAND2XL inst_it2_cellmath__57__61__I2175 (.Y(N2264), .A(N2277), .B(inst_cellmath__9[10]));
NAND2XL inst_it2_cellmath__57__61__I2176 (.Y(N2265), .A(N2277), .B(inst_cellmath__9[11]));
NAND2XL inst_it2_cellmath__57__61__I2177 (.Y(N2266), .A(N2277), .B(inst_cellmath__9[12]));
NAND2XL inst_it2_cellmath__57__61__I2178 (.Y(N2267), .A(N2277), .B(inst_cellmath__9[13]));
NAND2XL inst_it2_cellmath__57__61__I2179 (.Y(N2268), .A(N2277), .B(inst_cellmath__9[14]));
NAND2XL inst_it2_cellmath__57__61__I2180 (.Y(N2269), .A(N2277), .B(inst_cellmath__9[15]));
NAND2XL inst_it2_cellmath__57__61__I2181 (.Y(N2270), .A(N2277), .B(inst_cellmath__9[16]));
NAND2XL inst_it2_cellmath__57__61__I2182 (.Y(N2271), .A(N2277), .B(inst_cellmath__9[17]));
NAND2XL inst_it2_cellmath__57__61__I2183 (.Y(N2272), .A(N2277), .B(inst_cellmath__9[18]));
NAND2XL inst_it2_cellmath__57__61__I2184 (.Y(N2273), .A(N2277), .B(inst_cellmath__9[19]));
NAND2XL inst_it2_cellmath__57__61__I2185 (.Y(N2274), .A(N2277), .B(inst_cellmath__9[20]));
NAND2XL inst_it2_cellmath__57__61__I2186 (.Y(N2275), .A(N2277), .B(inst_it2_lookup1_cellmath__53[0]));
NAND2XL inst_it2_cellmath__57__61__I2187 (.Y(N2276), .A(N2277), .B(inst_it2_lookup1_cellmath__53[1]));
DFFQXL inst_cellmath__112_0_0__I168 (.Q(inst_cellmath__112[0]), .D(N1751), .CK(clk));
DFFQXL inst_cellmath__112_0_1__I169 (.Q(inst_cellmath__112[1]), .D(N1752), .CK(clk));
DFFQXL inst_cellmath__112_0_2__I170 (.Q(inst_cellmath__112[2]), .D(N1753), .CK(clk));
DFFQXL inst_cellmath__112_0_3__I171 (.Q(inst_cellmath__112[3]), .D(N1754), .CK(clk));
DFFQXL inst_cellmath__112_0_4__I172 (.Q(inst_cellmath__112[4]), .D(N1755), .CK(clk));
DFFQXL inst_cellmath__112_0_5__I173 (.Q(inst_cellmath__112[5]), .D(N1756), .CK(clk));
DFFQXL inst_cellmath__112_0_6__I174 (.Q(inst_cellmath__112[6]), .D(N1757), .CK(clk));
DFFQXL inst_cellmath__112_0_7__I175 (.Q(inst_cellmath__112[7]), .D(N1758), .CK(clk));
DFFQXL inst_cellmath__112_0_8__I176 (.Q(inst_cellmath__112[8]), .D(N1759), .CK(clk));
DFFQXL inst_cellmath__112_0_9__I177 (.Q(inst_cellmath__112[9]), .D(N1760), .CK(clk));
DFFQXL inst_cellmath__112_0_10__I178 (.Q(inst_cellmath__112[10]), .D(N1761), .CK(clk));
DFFQXL inst_cellmath__112_0_11__I179 (.Q(inst_cellmath__112[11]), .D(N1762), .CK(clk));
DFFQXL inst_cellmath__112_0_12__I180 (.Q(inst_cellmath__112[12]), .D(N1763), .CK(clk));
DFFQXL inst_cellmath__112_0_13__I181 (.Q(inst_cellmath__112[13]), .D(N1764), .CK(clk));
DFFQXL inst_cellmath__112_0_14__I182 (.Q(inst_cellmath__112[14]), .D(N1765), .CK(clk));
DFFQXL inst_cellmath__112_0_15__I183 (.Q(inst_cellmath__112[15]), .D(N1766), .CK(clk));
DFFQXL inst_cellmath__112_0_16__I184 (.Q(inst_cellmath__112[16]), .D(N1767), .CK(clk));
DFFQXL inst_cellmath__112_0_17__I185 (.Q(inst_cellmath__112[17]), .D(N1768), .CK(clk));
DFFQXL inst_cellmath__112_0_18__I186 (.Q(inst_cellmath__112[18]), .D(N1769), .CK(clk));
DFFQXL inst_cellmath__112_0_19__I187 (.Q(inst_cellmath__112[19]), .D(N1770), .CK(clk));
DFFQXL inst_cellmath__112_0_20__I188 (.Q(inst_cellmath__112[20]), .D(N1771), .CK(clk));
DFFQXL inst_cellmath__112_0_21__I189 (.Q(inst_cellmath__112[21]), .D(N1772), .CK(clk));
ADDHX1 inst_cellmath__120_0_I2189 (.CO(N13719), .S(inst_cellmath__120[1]), .A(inst_cellmath__16[1]), .B(inst_cellmath__17[1]));
ADDFX1 inst_cellmath__120_0_I2190 (.CO(N13661), .S(inst_cellmath__120[2]), .A(inst_cellmath__17[2]), .B(inst_cellmath__16[2]), .CI(N13719));
ADDFX1 inst_cellmath__120_0_I2191 (.CO(N13705), .S(inst_cellmath__120[3]), .A(inst_cellmath__17[3]), .B(inst_cellmath__16[3]), .CI(N13661));
ADDFX1 inst_cellmath__120_0_I2192 (.CO(N13753), .S(inst_cellmath__120[4]), .A(inst_cellmath__17[4]), .B(inst_cellmath__16[4]), .CI(N13705));
ADDFX1 inst_cellmath__120_0_I2193 (.CO(N13692), .S(inst_cellmath__120[5]), .A(inst_cellmath__17[5]), .B(inst_cellmath__16[5]), .CI(N13753));
ADDFX1 inst_cellmath__120_0_I2194 (.CO(N13738), .S(inst_cellmath__120[6]), .A(inst_cellmath__17[6]), .B(inst_cellmath__16[6]), .CI(N13692));
ADDFX1 inst_cellmath__120_0_I2195 (.CO(N13680), .S(inst_cellmath__120[7]), .A(inst_cellmath__17[7]), .B(inst_cellmath__16[7]), .CI(N13738));
ADDFX1 inst_cellmath__120_0_I2196 (.CO(N13725), .S(inst_cellmath__120[8]), .A(inst_cellmath__17[8]), .B(inst_cellmath__16[8]), .CI(N13680));
ADDFX1 inst_cellmath__120_0_I2197 (.CO(N13667), .S(inst_cellmath__120[9]), .A(inst_cellmath__17[9]), .B(inst_cellmath__16[9]), .CI(N13725));
ADDFX1 inst_cellmath__120_0_I2198 (.CO(N13712), .S(inst_cellmath__120[10]), .A(inst_cellmath__17[10]), .B(inst_cellmath__16[10]), .CI(N13667));
ADDFX1 inst_cellmath__120_0_I2199 (.CO(N13758), .S(inst_cellmath__120[11]), .A(inst_cellmath__17[11]), .B(inst_cellmath__16[11]), .CI(N13712));
ADDFX1 inst_cellmath__120_0_I2200 (.CO(N13697), .S(inst_cellmath__120[12]), .A(inst_cellmath__17[12]), .B(inst_cellmath__16[12]), .CI(N13758));
ADDFX1 inst_cellmath__120_0_I2201 (.CO(N13745), .S(inst_cellmath__120[13]), .A(inst_cellmath__17[13]), .B(inst_cellmath__16[13]), .CI(N13697));
ADDFX1 inst_cellmath__120_0_I2202 (.CO(N13685), .S(inst_cellmath__120[14]), .A(inst_cellmath__17[14]), .B(inst_cellmath__16[14]), .CI(N13745));
ADDFX1 inst_cellmath__120_0_I2203 (.CO(N13730), .S(inst_cellmath__120[15]), .A(inst_cellmath__17[15]), .B(inst_cellmath__16[15]), .CI(N13685));
ADDFX1 inst_cellmath__120_0_I2204 (.CO(N13673), .S(inst_cellmath__120[16]), .A(inst_cellmath__17[16]), .B(inst_cellmath__16[16]), .CI(N13730));
ADDFX1 inst_cellmath__120_0_I2205 (.CO(N13716), .S(inst_cellmath__120[17]), .A(inst_cellmath__17[17]), .B(inst_cellmath__16[17]), .CI(N13673));
ADDFX1 inst_cellmath__120_0_I2206 (.CO(N13658), .S(inst_cellmath__120[18]), .A(inst_cellmath__17[18]), .B(inst_cellmath__16[18]), .CI(N13716));
ADDFX1 inst_cellmath__120_0_I2207 (.CO(N13704), .S(inst_cellmath__120[19]), .A(inst_cellmath__17[19]), .B(inst_cellmath__16[19]), .CI(N13658));
ADDFX1 inst_cellmath__120_0_I2208 (.CO(N13750), .S(inst_cellmath__120[20]), .A(inst_cellmath__17[20]), .B(inst_cellmath__16[20]), .CI(N13704));
ADDFX1 inst_cellmath__120_0_I2209 (.CO(N13689), .S(inst_cellmath__120[21]), .A(inst_cellmath__16[21]), .B(inst_cellmath__17[21]), .CI(N13750));
ADDFX1 inst_cellmath__120_0_I2210 (.CO(N13737), .S(inst_cellmath__120[22]), .A(inst_cellmath__16[22]), .B(inst_cellmath__17[22]), .CI(N13689));
ADDFX1 inst_cellmath__120_0_I2211 (.CO(N13677), .S(inst_cellmath__120[23]), .A(inst_cellmath__16[23]), .B(inst_cellmath__17[23]), .CI(N13737));
ADDFX1 inst_cellmath__120_0_I2212 (.CO(N13722), .S(inst_cellmath__120[24]), .A(inst_cellmath__16[24]), .B(inst_cellmath__17[24]), .CI(N13677));
ADDFX1 inst_cellmath__120_0_I2213 (.CO(N13665), .S(inst_cellmath__120[25]), .A(inst_cellmath__16[25]), .B(inst_cellmath__17[25]), .CI(N13722));
DFFQXL inst_cellmath__44_0_0__I191 (.Q(inst_cellmath__44[0]), .D(inst_cellmath__40[0]), .CK(clk));
DFFQXL inst_cellmath__44_0_1__I192 (.Q(inst_cellmath__44[1]), .D(inst_cellmath__40[1]), .CK(clk));
DFFQXL inst_cellmath__44_0_2__I193 (.Q(inst_cellmath__44[2]), .D(inst_cellmath__40[2]), .CK(clk));
DFFQXL inst_cellmath__44_0_3__I194 (.Q(inst_cellmath__44[3]), .D(inst_cellmath__40[3]), .CK(clk));
DFFQXL inst_cellmath__44_0_4__I195 (.Q(inst_cellmath__44[4]), .D(inst_cellmath__40[4]), .CK(clk));
DFFQXL inst_cellmath__44_0_5__I196 (.Q(inst_cellmath__44[5]), .D(inst_cellmath__40[5]), .CK(clk));
DFFQXL inst_cellmath__44_0_6__I197 (.Q(inst_cellmath__44[6]), .D(inst_cellmath__40[6]), .CK(clk));
DFFQXL inst_cellmath__44_0_7__I198 (.Q(inst_cellmath__44[7]), .D(inst_cellmath__40[7]), .CK(clk));
DFFQXL inst_cellmath__44_0_8__I199 (.Q(inst_cellmath__44[8]), .D(inst_cellmath__40[8]), .CK(clk));
DFFQXL inst_cellmath__44_0_9__I200 (.Q(inst_cellmath__44[9]), .D(inst_cellmath__40[9]), .CK(clk));
DFFQXL inst_cellmath__44_0_10__I201 (.Q(inst_cellmath__44[10]), .D(inst_cellmath__40[10]), .CK(clk));
DFFQXL inst_cellmath__44_0_11__I202 (.Q(inst_cellmath__44[11]), .D(inst_cellmath__40[11]), .CK(clk));
DFFQXL inst_cellmath__44_0_12__I203 (.Q(inst_cellmath__44[12]), .D(inst_cellmath__40[12]), .CK(clk));
DFFQXL inst_cellmath__44_0_13__I204 (.Q(inst_cellmath__44[13]), .D(inst_cellmath__40[13]), .CK(clk));
DFFQXL inst_cellmath__44_0_14__I205 (.Q(inst_cellmath__44[14]), .D(inst_cellmath__40[14]), .CK(clk));
DFFQXL inst_cellmath__44_0_15__I206 (.Q(inst_cellmath__44[15]), .D(inst_cellmath__40[15]), .CK(clk));
DFFQXL inst_cellmath__44_0_16__I207 (.Q(inst_cellmath__44[16]), .D(inst_cellmath__40[16]), .CK(clk));
DFFQXL inst_cellmath__44_0_17__I208 (.Q(inst_cellmath__44[17]), .D(inst_cellmath__40[17]), .CK(clk));
DFFQXL inst_cellmath__44_0_18__I209 (.Q(inst_cellmath__44[18]), .D(inst_cellmath__40[18]), .CK(clk));
DFFQXL inst_cellmath__44_0_19__I210 (.Q(inst_cellmath__44[19]), .D(inst_cellmath__40[19]), .CK(clk));
DFFQXL inst_cellmath__44_0_20__I211 (.Q(inst_cellmath__44[20]), .D(inst_cellmath__40[20]), .CK(clk));
DFFQXL inst_cellmath__44_0_21__I212 (.Q(inst_cellmath__44[21]), .D(inst_cellmath__40[21]), .CK(clk));
DFFQXL inst_cellmath__44_0_22__I213 (.Q(inst_cellmath__44[22]), .D(inst_cellmath__40[22]), .CK(clk));
DFFQXL inst_cellmath__44_0_23__I214 (.Q(inst_cellmath__44[23]), .D(inst_cellmath__40[23]), .CK(clk));
DFFQXL inst_cellmath__44_0_24__I215 (.Q(inst_cellmath__44[24]), .D(inst_cellmath__40[24]), .CK(clk));
DFFQXL inst_cellmath__44_0_25__I216 (.Q(inst_cellmath__44[25]), .D(inst_cellmath__40[25]), .CK(clk));
DFFQXL inst_cellmath__44_0_26__I217 (.Q(inst_cellmath__44[26]), .D(inst_cellmath__40[26]), .CK(clk));
DFFQXL inst_cellmath__44_0_27__I218 (.Q(inst_cellmath__44[27]), .D(inst_cellmath__40[27]), .CK(clk));
DFFQXL inst_cellmath__44_0_28__I219 (.Q(inst_cellmath__44[28]), .D(inst_cellmath__40[28]), .CK(clk));
DFFQXL inst_cellmath__45_0_0__I220 (.Q(inst_cellmath__45[0]), .D(inst_cellmath__41[0]), .CK(clk));
DFFQXL inst_cellmath__45_0_1__I221 (.Q(inst_cellmath__45[1]), .D(inst_cellmath__41[1]), .CK(clk));
DFFQXL inst_cellmath__45_0_2__I222 (.Q(inst_cellmath__45[2]), .D(inst_cellmath__41[2]), .CK(clk));
DFFQXL inst_cellmath__45_0_3__I223 (.Q(inst_cellmath__45[3]), .D(inst_cellmath__41[3]), .CK(clk));
DFFQXL inst_cellmath__45_0_4__I224 (.Q(inst_cellmath__45[4]), .D(inst_cellmath__41[4]), .CK(clk));
DFFQXL inst_cellmath__45_0_5__I225 (.Q(inst_cellmath__45[5]), .D(inst_cellmath__41[5]), .CK(clk));
DFFQXL inst_cellmath__45_0_6__I226 (.Q(inst_cellmath__45[6]), .D(inst_cellmath__41[6]), .CK(clk));
DFFQXL inst_cellmath__45_0_7__I227 (.Q(inst_cellmath__45[7]), .D(inst_cellmath__41[7]), .CK(clk));
DFFQXL inst_cellmath__45_0_8__I228 (.Q(inst_cellmath__45[8]), .D(inst_cellmath__41[8]), .CK(clk));
DFFQXL inst_cellmath__45_0_9__I229 (.Q(inst_cellmath__45[9]), .D(inst_cellmath__41[9]), .CK(clk));
DFFQXL inst_cellmath__45_0_10__I230 (.Q(inst_cellmath__45[10]), .D(inst_cellmath__41[10]), .CK(clk));
DFFQXL inst_cellmath__45_0_11__I231 (.Q(inst_cellmath__45[11]), .D(inst_cellmath__41[11]), .CK(clk));
DFFQXL inst_cellmath__45_0_12__I232 (.Q(inst_cellmath__45[12]), .D(inst_cellmath__41[12]), .CK(clk));
DFFQXL inst_cellmath__45_0_13__I233 (.Q(inst_cellmath__45[13]), .D(inst_cellmath__41[13]), .CK(clk));
DFFQXL inst_cellmath__45_0_14__I234 (.Q(inst_cellmath__45[14]), .D(inst_cellmath__41[14]), .CK(clk));
DFFQXL inst_cellmath__45_0_15__I235 (.Q(inst_cellmath__45[15]), .D(inst_cellmath__41[15]), .CK(clk));
DFFQXL inst_cellmath__45_0_16__I236 (.Q(inst_cellmath__45[16]), .D(inst_cellmath__41[16]), .CK(clk));
DFFQXL inst_cellmath__45_0_17__I237 (.Q(inst_cellmath__45[17]), .D(inst_cellmath__41[17]), .CK(clk));
DFFQXL inst_cellmath__45_0_18__I238 (.Q(inst_cellmath__45[18]), .D(inst_cellmath__41[18]), .CK(clk));
DFFQXL inst_cellmath__45_0_19__I239 (.Q(inst_cellmath__45[19]), .D(inst_cellmath__41[19]), .CK(clk));
DFFQXL inst_cellmath__45_0_20__I240 (.Q(inst_cellmath__45[20]), .D(inst_cellmath__41[20]), .CK(clk));
DFFQXL inst_cellmath__45_0_21__I241 (.Q(inst_cellmath__45[21]), .D(inst_cellmath__41[21]), .CK(clk));
DFFQXL inst_cellmath__45_0_22__I242 (.Q(inst_cellmath__45[22]), .D(inst_cellmath__41[22]), .CK(clk));
DFFQXL inst_cellmath__45_0_23__I243 (.Q(inst_cellmath__45[23]), .D(inst_cellmath__41[23]), .CK(clk));
DFFQXL inst_cellmath__45_0_24__I244 (.Q(inst_cellmath__45[24]), .D(inst_cellmath__41[24]), .CK(clk));
DFFQXL inst_cellmath__45_0_25__I245 (.Q(inst_cellmath__45[25]), .D(inst_cellmath__41[25]), .CK(clk));
DFFQXL inst_cellmath__45_0_26__I246 (.Q(inst_cellmath__45[26]), .D(inst_cellmath__41[26]), .CK(clk));
DFFQXL inst_cellmath__45_0_27__I247 (.Q(inst_cellmath__45[27]), .D(inst_cellmath__41[27]), .CK(clk));
DFFQXL inst_cellmath__45_0_28__I248 (.Q(inst_cellmath__45[28]), .D(inst_cellmath__41[28]), .CK(clk));
MX2XL inst_cellmath__124_0_I2214 (.Y(inst_cellmath__124[0]), .A(inst_cellmath__44[0]), .B(inst_cellmath__45[0]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2215 (.Y(inst_cellmath__124[1]), .A(inst_cellmath__44[1]), .B(inst_cellmath__45[1]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2216 (.Y(inst_cellmath__124[2]), .A(inst_cellmath__44[2]), .B(inst_cellmath__45[2]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2217 (.Y(inst_cellmath__124[3]), .A(inst_cellmath__44[3]), .B(inst_cellmath__45[3]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2218 (.Y(inst_cellmath__124[4]), .A(inst_cellmath__44[4]), .B(inst_cellmath__45[4]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2219 (.Y(inst_cellmath__124[5]), .A(inst_cellmath__44[5]), .B(inst_cellmath__45[5]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2220 (.Y(inst_cellmath__124[6]), .A(inst_cellmath__44[6]), .B(inst_cellmath__45[6]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2221 (.Y(inst_cellmath__124[7]), .A(inst_cellmath__44[7]), .B(inst_cellmath__45[7]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2222 (.Y(inst_cellmath__124[8]), .A(inst_cellmath__44[8]), .B(inst_cellmath__45[8]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2223 (.Y(inst_cellmath__124[9]), .A(inst_cellmath__44[9]), .B(inst_cellmath__45[9]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2224 (.Y(inst_cellmath__124[10]), .A(inst_cellmath__44[10]), .B(inst_cellmath__45[10]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2225 (.Y(inst_cellmath__124[11]), .A(inst_cellmath__44[11]), .B(inst_cellmath__45[11]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2226 (.Y(inst_cellmath__124[12]), .A(inst_cellmath__44[12]), .B(inst_cellmath__45[12]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2227 (.Y(inst_cellmath__124[13]), .A(inst_cellmath__44[13]), .B(inst_cellmath__45[13]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2228 (.Y(inst_cellmath__124[14]), .A(inst_cellmath__44[14]), .B(inst_cellmath__45[14]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2229 (.Y(inst_cellmath__124[15]), .A(inst_cellmath__44[15]), .B(inst_cellmath__45[15]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2230 (.Y(inst_cellmath__124[16]), .A(inst_cellmath__44[16]), .B(inst_cellmath__45[16]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2231 (.Y(inst_cellmath__124[17]), .A(inst_cellmath__44[17]), .B(inst_cellmath__45[17]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2232 (.Y(inst_cellmath__124[18]), .A(inst_cellmath__44[18]), .B(inst_cellmath__45[18]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2233 (.Y(inst_cellmath__124[19]), .A(inst_cellmath__44[19]), .B(inst_cellmath__45[19]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2234 (.Y(inst_cellmath__124[20]), .A(inst_cellmath__44[20]), .B(inst_cellmath__45[20]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2235 (.Y(inst_cellmath__124[21]), .A(inst_cellmath__44[21]), .B(inst_cellmath__45[21]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2236 (.Y(inst_cellmath__124[22]), .A(inst_cellmath__44[22]), .B(inst_cellmath__45[22]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2237 (.Y(inst_cellmath__124[23]), .A(inst_cellmath__44[23]), .B(inst_cellmath__45[23]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2238 (.Y(inst_cellmath__124[24]), .A(inst_cellmath__44[24]), .B(inst_cellmath__45[24]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2239 (.Y(inst_cellmath__124[25]), .A(inst_cellmath__44[25]), .B(inst_cellmath__45[25]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2240 (.Y(inst_cellmath__124[26]), .A(inst_cellmath__44[26]), .B(inst_cellmath__45[26]), .S0(inst_cellmath__120[25]));
MX2XL inst_cellmath__124_0_I2241 (.Y(inst_cellmath__124[27]), .A(inst_cellmath__44[27]), .B(inst_cellmath__45[27]), .S0(inst_cellmath__120[25]));
MXI2XL cynw_cm_float_div_ieee_I4146 (.Y(inst_cellmath__122), .A(inst_cellmath__44[28]), .B(inst_cellmath__45[28]), .S0(inst_cellmath__120[25]));
INVXL inst_cellmath__125_0_I2243 (.Y(N13935), .A(inst_cellmath__122));
INVXL inst_cellmath__125_0_I2244 (.Y(N13952), .A(N13935));
MX2XL inst_cellmath__125_0_I2245 (.Y(inst_cellmath__125[0]), .A(inst_cellmath__124[5]), .B(inst_cellmath__124[4]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2246 (.Y(inst_cellmath__125[1]), .A(inst_cellmath__124[6]), .B(inst_cellmath__124[5]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2247 (.Y(inst_cellmath__125[2]), .A(inst_cellmath__124[7]), .B(inst_cellmath__124[6]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2248 (.Y(inst_cellmath__125[3]), .A(inst_cellmath__124[8]), .B(inst_cellmath__124[7]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2249 (.Y(inst_cellmath__125[4]), .A(inst_cellmath__124[9]), .B(inst_cellmath__124[8]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2250 (.Y(inst_cellmath__125[5]), .A(inst_cellmath__124[10]), .B(inst_cellmath__124[9]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2251 (.Y(inst_cellmath__125[6]), .A(inst_cellmath__124[11]), .B(inst_cellmath__124[10]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2252 (.Y(inst_cellmath__125[7]), .A(inst_cellmath__124[12]), .B(inst_cellmath__124[11]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2253 (.Y(inst_cellmath__125[8]), .A(inst_cellmath__124[13]), .B(inst_cellmath__124[12]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2254 (.Y(inst_cellmath__125[9]), .A(inst_cellmath__124[14]), .B(inst_cellmath__124[13]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2255 (.Y(inst_cellmath__125[10]), .A(inst_cellmath__124[15]), .B(inst_cellmath__124[14]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2256 (.Y(inst_cellmath__125[11]), .A(inst_cellmath__124[16]), .B(inst_cellmath__124[15]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2257 (.Y(inst_cellmath__125[12]), .A(inst_cellmath__124[17]), .B(inst_cellmath__124[16]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2258 (.Y(inst_cellmath__125[13]), .A(inst_cellmath__124[18]), .B(inst_cellmath__124[17]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2259 (.Y(inst_cellmath__125[14]), .A(inst_cellmath__124[19]), .B(inst_cellmath__124[18]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2260 (.Y(inst_cellmath__125[15]), .A(inst_cellmath__124[20]), .B(inst_cellmath__124[19]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2261 (.Y(inst_cellmath__125[16]), .A(inst_cellmath__124[21]), .B(inst_cellmath__124[20]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2262 (.Y(inst_cellmath__125[17]), .A(inst_cellmath__124[22]), .B(inst_cellmath__124[21]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2263 (.Y(inst_cellmath__125[18]), .A(inst_cellmath__124[23]), .B(inst_cellmath__124[22]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2264 (.Y(inst_cellmath__125[19]), .A(inst_cellmath__124[24]), .B(inst_cellmath__124[23]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2265 (.Y(inst_cellmath__125[20]), .A(inst_cellmath__124[25]), .B(inst_cellmath__124[24]), .S0(N13952));
MX2XL inst_cellmath__125_0_I2266 (.Y(inst_cellmath__125[21]), .A(inst_cellmath__124[26]), .B(inst_cellmath__124[25]), .S0(N13952));
MXI2XL inst_cellmath__125_0_I2267 (.Y(inst_cellmath__125[22]), .A(inst_cellmath__124[27]), .B(inst_cellmath__124[26]), .S0(N13952));
MX2XL cynw_cm_float_div_ieee_I2268 (.Y(inst_cellmath__126), .A(inst_cellmath__124[4]), .B(inst_cellmath__124[3]), .S0(inst_cellmath__122));
ADDHX1 inst_cellmath__129_0_I2269 (.CO(N14058), .S(inst_cellmath__129[0]), .A(inst_cellmath__126), .B(inst_cellmath__125[0]));
ADDHX1 inst_cellmath__129_0_I2270 (.CO(N14047), .S(inst_cellmath__129[1]), .A(inst_cellmath__125[1]), .B(N14058));
ADDHX1 inst_cellmath__129_0_I2271 (.CO(N14038), .S(inst_cellmath__129[2]), .A(inst_cellmath__125[2]), .B(N14047));
ADDHX1 inst_cellmath__129_0_I2272 (.CO(N14030), .S(inst_cellmath__129[3]), .A(inst_cellmath__125[3]), .B(N14038));
ADDHX1 inst_cellmath__129_0_I2273 (.CO(N14020), .S(inst_cellmath__129[4]), .A(inst_cellmath__125[4]), .B(N14030));
ADDHX1 inst_cellmath__129_0_I2274 (.CO(N14012), .S(inst_cellmath__129[5]), .A(inst_cellmath__125[5]), .B(N14020));
ADDHX1 inst_cellmath__129_0_I2275 (.CO(N14072), .S(inst_cellmath__129[6]), .A(inst_cellmath__125[6]), .B(N14012));
ADDHX1 inst_cellmath__129_0_I2276 (.CO(N14063), .S(inst_cellmath__129[7]), .A(inst_cellmath__125[7]), .B(N14072));
ADDHX1 inst_cellmath__129_0_I2277 (.CO(N14055), .S(inst_cellmath__129[8]), .A(inst_cellmath__125[8]), .B(N14063));
ADDHX1 inst_cellmath__129_0_I2278 (.CO(N14045), .S(inst_cellmath__129[9]), .A(inst_cellmath__125[9]), .B(N14055));
ADDHX1 inst_cellmath__129_0_I2279 (.CO(N14035), .S(inst_cellmath__129[10]), .A(inst_cellmath__125[10]), .B(N14045));
ADDHX1 inst_cellmath__129_0_I2280 (.CO(N14027), .S(inst_cellmath__129[11]), .A(inst_cellmath__125[11]), .B(N14035));
ADDHX1 inst_cellmath__129_0_I2281 (.CO(N14018), .S(inst_cellmath__129[12]), .A(inst_cellmath__125[12]), .B(N14027));
ADDHX1 inst_cellmath__129_0_I2282 (.CO(N14010), .S(inst_cellmath__129[13]), .A(inst_cellmath__125[13]), .B(N14018));
ADDHX1 inst_cellmath__129_0_I2283 (.CO(N14070), .S(inst_cellmath__129[14]), .A(inst_cellmath__125[14]), .B(N14010));
ADDHX1 inst_cellmath__129_0_I2284 (.CO(N14061), .S(inst_cellmath__129[15]), .A(inst_cellmath__125[15]), .B(N14070));
ADDHX1 inst_cellmath__129_0_I2285 (.CO(N14053), .S(inst_cellmath__129[16]), .A(inst_cellmath__125[16]), .B(N14061));
ADDHX1 inst_cellmath__129_0_I2286 (.CO(N14043), .S(inst_cellmath__129[17]), .A(inst_cellmath__125[17]), .B(N14053));
ADDHX1 inst_cellmath__129_0_I2287 (.CO(N14033), .S(inst_cellmath__129[18]), .A(inst_cellmath__125[18]), .B(N14043));
ADDHX1 inst_cellmath__129_0_I2288 (.CO(N14025), .S(inst_cellmath__129[19]), .A(inst_cellmath__125[19]), .B(N14033));
ADDHX1 inst_cellmath__129_0_I2289 (.CO(N14016), .S(inst_cellmath__129[20]), .A(inst_cellmath__125[20]), .B(N14025));
ADDHX1 inst_cellmath__129_0_I2290 (.CO(N14077), .S(inst_cellmath__129[21]), .A(inst_cellmath__125[21]), .B(N14016));
XNOR2X1 inst_cellmath__129_0_I2291 (.Y(inst_cellmath__129[22]), .A(inst_cellmath__125[22]), .B(N14077));
OR4X1 cynw_cm_float_div_ieee_I9187 (.Y(N1682), .A(inst_cellmath__124[2]), .B(inst_cellmath__124[1]), .C(inst_cellmath__124[3]), .D(inst_cellmath__124[0]));
OR3XL cynw_cm_float_div_ieee_I2295 (.Y(N1681), .A(inst_cellmath__124[0]), .B(inst_cellmath__124[1]), .C(inst_cellmath__124[2]));
MX2XL cynw_cm_float_div_ieee_I2296 (.Y(inst_cellmath__127), .A(N1682), .B(N1681), .S0(inst_cellmath__122));
NOR3XL inst_cellmath__130__105__I2297 (.Y(N14181), .A(inst_cellmath__120[1]), .B(inst_cellmath__120[2]), .C(inst_cellmath__120[6]));
NOR3XL inst_cellmath__130__105__I2298 (.Y(N14169), .A(inst_cellmath__120[5]), .B(inst_cellmath__120[11]), .C(inst_cellmath__120[15]));
NOR3BXL inst_cellmath__130__105__I2299 (.Y(N14179), .AN(N14181), .B(inst_cellmath__120[14]), .C(inst_cellmath__120[12]));
NOR3XL inst_cellmath__130__105__I2300 (.Y(N14153), .A(inst_cellmath__120[10]), .B(inst_cellmath__120[8]), .C(inst_cellmath__120[9]));
NOR3XL inst_cellmath__130__105__I2301 (.Y(N14173), .A(inst_cellmath__120[13]), .B(inst_cellmath__120[16]), .C(inst_cellmath__120[19]));
NOR2XL inst_cellmath__130__105__I2302 (.Y(N14185), .A(inst_cellmath__120[20]), .B(inst_cellmath__120[18]));
NOR4X1 inst_cellmath__130__105__I2303 (.Y(N14149), .A(inst_cellmath__120[4]), .B(inst_cellmath__120[3]), .C(inst_cellmath__120[7]), .D(inst_cellmath__120[17]));
NOR2XL inst_cellmath__130__105__I2304 (.Y(N14158), .A(inst_cellmath__120[22]), .B(inst_cellmath__120[24]));
NAND2XL inst_cellmath__130__105__I2306 (.Y(N14177), .A(N14179), .B(N14169));
NAND4XL inst_cellmath__130__105__I2309 (.Y(N14146), .A(N14153), .B(N14185), .C(N14149), .D(N14158));
NOR4BX1 inst_cellmath__130__105__I9188 (.Y(N14165), .AN(N14173), .B(inst_cellmath__120[21]), .C(N14146), .D(inst_cellmath__120[23]));
NOR2XL inst_cellmath__130__105__I2308 (.Y(N14182), .A(inst_cellmath__120[25]), .B(N14177));
NAND3BXL inst_cellmath__130__105__I2311 (.Y(N14160), .AN(inst_cellmath__127), .B(N14182), .C(N14165));
OA21X1 cynw_cm_float_div_ieee_I4147 (.Y(N1922), .A0(N14160), .A1(inst_cellmath__125[0]), .B0(inst_cellmath__129[0]));
INVXL cynw_cm_float_div_ieee_I259 (.Y(N1322), .A(accept));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_0__I260 (.q(inst_cellmath__13[0]), .r(N1322), .d(inst_cellmath__12[0]), .clk(clk));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_1__I261 (.q(inst_cellmath__13[1]), .r(N1322), .d(inst_cellmath__12[1]), .clk(clk));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_2__I262 (.q(inst_cellmath__13[2]), .r(N1322), .d(inst_cellmath__12[2]), .clk(clk));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_3__I263 (.q(inst_cellmath__13[3]), .r(N1322), .d(inst_cellmath__12[3]), .clk(clk));
ADDHX1 inst_cellmath__12__18__I2315 (.CO(N14214), .S(N1324), .A(inst_cellmath__13[1]), .B(inst_cellmath__13[0]));
ADDHX1 inst_cellmath__12__18__I2316 (.CO(N14213), .S(N1325), .A(inst_cellmath__13[2]), .B(N14214));
XOR2XL inst_cellmath__12__18__I2317 (.Y(N1326), .A(inst_cellmath__13[3]), .B(N14213));
AND4XL cynw_cm_float_div_ieee_I9189 (.Y(N1327), .A(inst_cellmath__13[3]), .B(inst_cellmath__13[0]), .C(inst_cellmath__13[1]), .D(inst_cellmath__13[2]));
NAND2BXL inst_cellmath__12_0_I4148 (.Y(inst_cellmath__12[0]), .AN(N1327), .B(inst_cellmath__13[0]));
OR2XL inst_cellmath__12_0_I2322 (.Y(inst_cellmath__12[1]), .A(N1327), .B(N1324));
OR2XL inst_cellmath__12_0_I2323 (.Y(inst_cellmath__12[2]), .A(N1327), .B(N1325));
OR2XL inst_cellmath__12_0_I2324 (.Y(inst_cellmath__12[3]), .A(N1327), .B(N1326));
NAND2BXL inst_cellmath__46_0_I2326 (.Y(inst_cellmath__46[0]), .AN(inst_cellmath__44[0]), .B(N12658));
AND2XL inst_cellmath__46_0_I2327 (.Y(inst_cellmath__46[1]), .A(N12658), .B(inst_cellmath__44[1]));
AND2XL inst_cellmath__46_0_I2328 (.Y(inst_cellmath__46[2]), .A(N12658), .B(inst_cellmath__44[2]));
AND2XL inst_cellmath__46_0_I2329 (.Y(inst_cellmath__46[3]), .A(N12658), .B(inst_cellmath__44[3]));
AND2XL inst_cellmath__46_0_I2330 (.Y(inst_cellmath__46[4]), .A(N12658), .B(inst_cellmath__44[4]));
AND2XL inst_cellmath__46_0_I2331 (.Y(inst_cellmath__46[5]), .A(N12658), .B(inst_cellmath__44[5]));
AND2XL inst_cellmath__46_0_I2332 (.Y(inst_cellmath__46[6]), .A(N12658), .B(inst_cellmath__44[6]));
AND2XL inst_cellmath__46_0_I2333 (.Y(inst_cellmath__46[7]), .A(N12658), .B(inst_cellmath__44[7]));
AND2XL inst_cellmath__46_0_I2334 (.Y(inst_cellmath__46[8]), .A(N12658), .B(inst_cellmath__44[8]));
AND2XL inst_cellmath__46_0_I2335 (.Y(inst_cellmath__46[9]), .A(N12658), .B(inst_cellmath__44[9]));
AND2XL inst_cellmath__46_0_I2336 (.Y(inst_cellmath__46[10]), .A(N12658), .B(inst_cellmath__44[10]));
AND2XL inst_cellmath__46_0_I2337 (.Y(inst_cellmath__46[11]), .A(N12658), .B(inst_cellmath__44[11]));
AND2XL inst_cellmath__46_0_I2338 (.Y(inst_cellmath__46[12]), .A(N12658), .B(inst_cellmath__44[12]));
AND2XL inst_cellmath__46_0_I2339 (.Y(inst_cellmath__46[13]), .A(N12658), .B(inst_cellmath__44[13]));
AND2XL inst_cellmath__46_0_I2340 (.Y(inst_cellmath__46[14]), .A(N12658), .B(inst_cellmath__44[14]));
AND2XL inst_cellmath__46_0_I2341 (.Y(inst_cellmath__46[15]), .A(N12658), .B(inst_cellmath__44[15]));
AND2XL inst_cellmath__46_0_I2342 (.Y(inst_cellmath__46[16]), .A(N12658), .B(inst_cellmath__44[16]));
AND2XL inst_cellmath__46_0_I2343 (.Y(inst_cellmath__46[17]), .A(N12658), .B(inst_cellmath__44[17]));
AND2XL inst_cellmath__46_0_I2344 (.Y(inst_cellmath__46[18]), .A(N12658), .B(inst_cellmath__44[18]));
AND2XL inst_cellmath__46_0_I2345 (.Y(inst_cellmath__46[19]), .A(N12658), .B(inst_cellmath__44[19]));
AND2XL inst_cellmath__46_0_I2346 (.Y(inst_cellmath__46[20]), .A(N12658), .B(inst_cellmath__44[20]));
AND2XL inst_cellmath__46_0_I2347 (.Y(inst_cellmath__46[21]), .A(N12658), .B(inst_cellmath__44[21]));
AND2XL inst_cellmath__46_0_I2348 (.Y(inst_cellmath__46[22]), .A(N12658), .B(inst_cellmath__44[22]));
AND2XL inst_cellmath__46_0_I2349 (.Y(inst_cellmath__46[23]), .A(N12658), .B(inst_cellmath__44[23]));
AND2XL inst_cellmath__46_0_I2350 (.Y(inst_cellmath__46[24]), .A(N12658), .B(inst_cellmath__44[24]));
NOR2BX1 inst_cellmath__47_0_I2353 (.Y(inst_cellmath__47[0]), .AN(inst_cellmath__45[0]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2354 (.Y(inst_cellmath__47[1]), .AN(inst_cellmath__45[1]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2355 (.Y(inst_cellmath__47[2]), .AN(inst_cellmath__45[2]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2356 (.Y(inst_cellmath__47[3]), .AN(inst_cellmath__45[3]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2357 (.Y(inst_cellmath__47[4]), .AN(inst_cellmath__45[4]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2358 (.Y(inst_cellmath__47[5]), .AN(inst_cellmath__45[5]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2359 (.Y(inst_cellmath__47[6]), .AN(inst_cellmath__45[6]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2360 (.Y(inst_cellmath__47[7]), .AN(inst_cellmath__45[7]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2361 (.Y(inst_cellmath__47[8]), .AN(inst_cellmath__45[8]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2362 (.Y(inst_cellmath__47[9]), .AN(inst_cellmath__45[9]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2363 (.Y(inst_cellmath__47[10]), .AN(inst_cellmath__45[10]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2364 (.Y(inst_cellmath__47[11]), .AN(inst_cellmath__45[11]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2365 (.Y(inst_cellmath__47[12]), .AN(inst_cellmath__45[12]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2366 (.Y(inst_cellmath__47[13]), .AN(inst_cellmath__45[13]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2367 (.Y(inst_cellmath__47[14]), .AN(inst_cellmath__45[14]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2368 (.Y(inst_cellmath__47[15]), .AN(inst_cellmath__45[15]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2369 (.Y(inst_cellmath__47[16]), .AN(inst_cellmath__45[16]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2370 (.Y(inst_cellmath__47[17]), .AN(inst_cellmath__45[17]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2371 (.Y(inst_cellmath__47[18]), .AN(inst_cellmath__45[18]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2372 (.Y(inst_cellmath__47[19]), .AN(inst_cellmath__45[19]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2373 (.Y(inst_cellmath__47[20]), .AN(inst_cellmath__45[20]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2374 (.Y(inst_cellmath__47[21]), .AN(inst_cellmath__45[21]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2375 (.Y(inst_cellmath__47[22]), .AN(inst_cellmath__45[22]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2376 (.Y(inst_cellmath__47[23]), .AN(inst_cellmath__45[23]), .B(inst_cellmath__38__W0[2]));
NOR2BX1 inst_cellmath__47_0_I2377 (.Y(inst_cellmath__47[24]), .AN(inst_cellmath__45[24]), .B(inst_cellmath__38__W0[2]));
NAND2XL cynw_cm_float_div_ieee_I2378 (.Y(N1417), .A(inst_lookup0_cellmath__29[1]), .B(inst_cellmath__42[0]));
MX2XL cynw_cm_float_div_ieee_I2379 (.Y(inst_cellmath__42[1]), .A(inst_lookup0_cellmath__29[1]), .B(N1417), .S0(inst_lookup0_cellmath__29[2]));
MX2XL cynw_cm_float_div_ieee_I2381 (.Y(inst_cellmath__42[2]), .A(inst_cellmath__47[0]), .B(inst_cellmath__46[0]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2382 (.Y(inst_cellmath__42[3]), .A(inst_cellmath__47[1]), .B(inst_cellmath__46[1]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2383 (.Y(inst_cellmath__42[4]), .A(inst_cellmath__47[2]), .B(inst_cellmath__46[2]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2384 (.Y(inst_cellmath__42[5]), .A(inst_cellmath__47[3]), .B(inst_cellmath__46[3]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2385 (.Y(inst_cellmath__42[6]), .A(inst_cellmath__47[4]), .B(inst_cellmath__46[4]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2386 (.Y(inst_cellmath__42[7]), .A(inst_cellmath__47[5]), .B(inst_cellmath__46[5]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2387 (.Y(inst_cellmath__42[8]), .A(inst_cellmath__47[6]), .B(inst_cellmath__46[6]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2388 (.Y(inst_cellmath__42[9]), .A(inst_cellmath__47[7]), .B(inst_cellmath__46[7]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2389 (.Y(inst_cellmath__42[10]), .A(inst_cellmath__47[8]), .B(inst_cellmath__46[8]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2390 (.Y(inst_cellmath__42[11]), .A(inst_cellmath__47[9]), .B(inst_cellmath__46[9]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2391 (.Y(inst_cellmath__42[12]), .A(inst_cellmath__47[10]), .B(inst_cellmath__46[10]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2392 (.Y(inst_cellmath__42[13]), .A(inst_cellmath__47[11]), .B(inst_cellmath__46[11]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2393 (.Y(inst_cellmath__42[14]), .A(inst_cellmath__47[12]), .B(inst_cellmath__46[12]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2394 (.Y(inst_cellmath__42[15]), .A(inst_cellmath__47[13]), .B(inst_cellmath__46[13]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2395 (.Y(inst_cellmath__42[16]), .A(inst_cellmath__47[14]), .B(inst_cellmath__46[14]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2396 (.Y(inst_cellmath__42[17]), .A(inst_cellmath__47[15]), .B(inst_cellmath__46[15]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2397 (.Y(inst_cellmath__42[18]), .A(inst_cellmath__47[16]), .B(inst_cellmath__46[16]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2398 (.Y(inst_cellmath__42[19]), .A(inst_cellmath__47[17]), .B(inst_cellmath__46[17]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2399 (.Y(inst_cellmath__42[20]), .A(inst_cellmath__47[18]), .B(inst_cellmath__46[18]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2400 (.Y(inst_cellmath__42[21]), .A(inst_cellmath__47[19]), .B(inst_cellmath__46[19]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2401 (.Y(inst_cellmath__42[22]), .A(inst_cellmath__47[20]), .B(inst_cellmath__46[20]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2402 (.Y(inst_cellmath__42[23]), .A(inst_cellmath__47[21]), .B(inst_cellmath__46[21]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2403 (.Y(inst_cellmath__42[24]), .A(inst_cellmath__47[22]), .B(inst_cellmath__46[22]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2404 (.Y(inst_cellmath__42[25]), .A(inst_cellmath__47[23]), .B(inst_cellmath__46[23]), .S0(inst_it2_cellmath__60[3]));
MX2XL cynw_cm_float_div_ieee_I2405 (.Y(inst_cellmath__42[26]), .A(inst_cellmath__47[24]), .B(inst_cellmath__46[24]), .S0(inst_it2_cellmath__60[3]));
XOR2XL cynw_cm_float_div_ieee_I2407 (.Y(inst_cellmath__43[1]), .A(inst_cellmath__42[1]), .B(inst_cellmath__43[0]));
OA21X1 inst_cellmath__43_0_I4150 (.Y(N14594), .A0(inst_cellmath__42[0]), .A1(inst_cellmath__42[1]), .B0(inst_it2_cellmath__60[4]));
MX2XL inst_cellmath__43_0_I2412 (.Y(inst_cellmath__43[2]), .A(inst_cellmath__47[0]), .B(inst_cellmath__46[0]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2413 (.Y(inst_cellmath__43[3]), .A(inst_cellmath__47[1]), .B(inst_cellmath__46[1]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2414 (.Y(inst_cellmath__43[4]), .A(inst_cellmath__47[2]), .B(inst_cellmath__46[2]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2415 (.Y(inst_cellmath__43[5]), .A(inst_cellmath__47[3]), .B(inst_cellmath__46[3]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2416 (.Y(inst_cellmath__43[6]), .A(inst_cellmath__47[4]), .B(inst_cellmath__46[4]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2417 (.Y(inst_cellmath__43[7]), .A(inst_cellmath__47[5]), .B(inst_cellmath__46[5]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2418 (.Y(inst_cellmath__43[8]), .A(inst_cellmath__47[6]), .B(inst_cellmath__46[6]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2419 (.Y(inst_cellmath__43[9]), .A(inst_cellmath__47[7]), .B(inst_cellmath__46[7]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2420 (.Y(inst_cellmath__43[10]), .A(inst_cellmath__47[8]), .B(inst_cellmath__46[8]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2421 (.Y(inst_cellmath__43[11]), .A(inst_cellmath__47[9]), .B(inst_cellmath__46[9]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2422 (.Y(inst_cellmath__43[12]), .A(inst_cellmath__47[10]), .B(inst_cellmath__46[10]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2423 (.Y(inst_cellmath__43[13]), .A(inst_cellmath__47[11]), .B(inst_cellmath__46[11]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2424 (.Y(inst_cellmath__43[14]), .A(inst_cellmath__47[12]), .B(inst_cellmath__46[12]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2425 (.Y(inst_cellmath__43[15]), .A(inst_cellmath__47[13]), .B(inst_cellmath__46[13]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2426 (.Y(inst_cellmath__43[16]), .A(inst_cellmath__47[14]), .B(inst_cellmath__46[14]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2427 (.Y(inst_cellmath__43[17]), .A(inst_cellmath__47[15]), .B(inst_cellmath__46[15]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2428 (.Y(inst_cellmath__43[18]), .A(inst_cellmath__47[16]), .B(inst_cellmath__46[16]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2429 (.Y(inst_cellmath__43[19]), .A(inst_cellmath__47[17]), .B(inst_cellmath__46[17]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2430 (.Y(inst_cellmath__43[20]), .A(inst_cellmath__47[18]), .B(inst_cellmath__46[18]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2431 (.Y(inst_cellmath__43[21]), .A(inst_cellmath__47[19]), .B(inst_cellmath__46[19]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2432 (.Y(inst_cellmath__43[22]), .A(inst_cellmath__47[20]), .B(inst_cellmath__46[20]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2433 (.Y(inst_cellmath__43[23]), .A(inst_cellmath__47[21]), .B(inst_cellmath__46[21]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2434 (.Y(inst_cellmath__43[24]), .A(inst_cellmath__47[22]), .B(inst_cellmath__46[22]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2435 (.Y(inst_cellmath__43[25]), .A(inst_cellmath__47[23]), .B(inst_cellmath__46[23]), .S0(N14594));
MX2XL inst_cellmath__43_0_I2436 (.Y(inst_cellmath__43[26]), .A(inst_cellmath__47[24]), .B(inst_cellmath__46[24]), .S0(N14594));
INVXL inst_it2_cellmath__56_2mx_I2437 (.Y(inst_cellmath__14[2]), .A(inst_it2_lookup1_cellmath__55[2]));
INVX1 inst_it2_cellmath__56_2mx_I2438 (.Y(N14648), .A(inst_cellmath__14[2]));
XNOR2X1 inst_it2_cellmath__56_2mx_I2439 (.Y(inst_it2_cellmath__63__W1[1]), .A(N2201), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2440 (.Y(inst_it2_cellmath__56[2]), .A(N2202), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2441 (.Y(inst_it2_cellmath__56[3]), .A(N2203), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2442 (.Y(inst_it2_cellmath__56[4]), .A(N2204), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2443 (.Y(inst_it2_cellmath__56[5]), .A(N2205), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2444 (.Y(inst_it2_cellmath__56[6]), .A(N2206), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2445 (.Y(inst_it2_cellmath__56[7]), .A(N2207), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2446 (.Y(inst_it2_cellmath__56[8]), .A(N2208), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2447 (.Y(inst_it2_cellmath__56[9]), .A(N2209), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2448 (.Y(inst_it2_cellmath__56[10]), .A(N2210), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2449 (.Y(inst_it2_cellmath__56[11]), .A(N2211), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2450 (.Y(inst_it2_cellmath__56[12]), .A(N2212), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2451 (.Y(inst_it2_cellmath__56[13]), .A(N2213), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2452 (.Y(inst_it2_cellmath__56[14]), .A(N2214), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2453 (.Y(inst_it2_cellmath__56[15]), .A(N2215), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2454 (.Y(inst_it2_cellmath__56[16]), .A(N2216), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2455 (.Y(inst_it2_cellmath__56[17]), .A(N2217), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2456 (.Y(inst_it2_cellmath__56[18]), .A(N2218), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2457 (.Y(inst_it2_cellmath__56[19]), .A(N2219), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2458 (.Y(inst_it2_cellmath__56[20]), .A(N2220), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2459 (.Y(inst_it2_cellmath__56[21]), .A(N2221), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2460 (.Y(inst_it2_cellmath__56[22]), .A(N2222), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2461 (.Y(inst_it2_cellmath__56[23]), .A(N2223), .B(N14648));
XNOR2X1 inst_it2_cellmath__56_2mx_I2462 (.Y(inst_it2_cellmath__56[24]), .A(N2224), .B(N14648));
INVXL cynw_cm_float_div_ieee_I2465 (.Y(inst_it2_cellmath__57[1]), .A(N14648));
MXI2XL cynw_cm_float_div_ieee_I2466 (.Y(inst_it2_cellmath__57[2]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2254));
MXI2XL cynw_cm_float_div_ieee_I2467 (.Y(inst_it2_cellmath__57[3]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2255));
MXI2XL cynw_cm_float_div_ieee_I2468 (.Y(inst_it2_cellmath__57[4]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2256));
MXI2XL cynw_cm_float_div_ieee_I2469 (.Y(inst_it2_cellmath__57[5]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2257));
MXI2XL cynw_cm_float_div_ieee_I2470 (.Y(inst_it2_cellmath__57[6]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2258));
MXI2XL cynw_cm_float_div_ieee_I2471 (.Y(inst_it2_cellmath__57[7]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2259));
MXI2XL cynw_cm_float_div_ieee_I2472 (.Y(inst_it2_cellmath__57[8]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2260));
MXI2XL cynw_cm_float_div_ieee_I2473 (.Y(inst_it2_cellmath__57[9]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2261));
MXI2XL cynw_cm_float_div_ieee_I2474 (.Y(inst_it2_cellmath__57[10]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2262));
MXI2XL cynw_cm_float_div_ieee_I2475 (.Y(inst_it2_cellmath__57[11]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2263));
MXI2XL cynw_cm_float_div_ieee_I2476 (.Y(inst_it2_cellmath__57[12]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2264));
MXI2XL cynw_cm_float_div_ieee_I2477 (.Y(inst_it2_cellmath__57[13]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2265));
MXI2XL cynw_cm_float_div_ieee_I2478 (.Y(inst_it2_cellmath__57[14]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2266));
MXI2XL cynw_cm_float_div_ieee_I2479 (.Y(inst_it2_cellmath__57[15]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2267));
MXI2XL cynw_cm_float_div_ieee_I2480 (.Y(inst_it2_cellmath__57[16]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2268));
MXI2XL cynw_cm_float_div_ieee_I2481 (.Y(inst_it2_cellmath__57[17]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2269));
MXI2XL cynw_cm_float_div_ieee_I2482 (.Y(inst_it2_cellmath__57[18]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2270));
MXI2XL cynw_cm_float_div_ieee_I2483 (.Y(inst_it2_cellmath__57[19]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2271));
MXI2XL cynw_cm_float_div_ieee_I2484 (.Y(inst_it2_cellmath__57[20]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2272));
MXI2XL cynw_cm_float_div_ieee_I2485 (.Y(inst_it2_cellmath__57[21]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2273));
MXI2XL cynw_cm_float_div_ieee_I2486 (.Y(inst_it2_cellmath__57[22]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2274));
MXI2XL cynw_cm_float_div_ieee_I2487 (.Y(inst_it2_cellmath__57[23]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2275));
MXI2XL cynw_cm_float_div_ieee_I2488 (.Y(inst_it2_cellmath__57[24]), .A(inst_it2_cellmath__57[1]), .B(N14648), .S0(N2276));
MXI2XL cynw_cm_float_div_ieee_I2489 (.Y(inst_it2_cellmath__57[25]), .A(N14648), .B(inst_it2_cellmath__57[1]), .S0(N2277));
ADDFX1 inst_fa_1820_10_I2491 (.CO(inst_it2_cellmath__62__W0[3]), .S(inst_it2_cellmath__62__W1[3]), .A(inst_it2_cellmath__61[3]), .B(inst_it2_cellmath__60[3]), .CI(inst_it2_cellmath__56[3]));
ADDFX1 inst_fa_1820_10_I2492 (.CO(inst_it2_cellmath__62__W0[4]), .S(inst_it2_cellmath__62__W1[4]), .A(inst_it2_cellmath__61[4]), .B(inst_it2_cellmath__60[4]), .CI(inst_it2_cellmath__56[4]));
ADDFX1 inst_fa_1820_10_I2493 (.CO(inst_it2_cellmath__62__W0[5]), .S(inst_it2_cellmath__62__W1[5]), .A(inst_it2_cellmath__61[5]), .B(inst_it2_cellmath__60[5]), .CI(inst_it2_cellmath__56[5]));
ADDFX1 inst_fa_1820_10_I2494 (.CO(inst_it2_cellmath__62__W0[6]), .S(inst_it2_cellmath__62__W1[6]), .A(inst_it2_cellmath__61[6]), .B(inst_it2_cellmath__60[6]), .CI(inst_it2_cellmath__56[6]));
ADDFX1 inst_fa_1820_10_I2495 (.CO(inst_it2_cellmath__62__W0[7]), .S(inst_it2_cellmath__62__W1[7]), .A(inst_it2_cellmath__61[7]), .B(inst_it2_cellmath__60[7]), .CI(inst_it2_cellmath__56[7]));
ADDFX1 inst_fa_1820_10_I2496 (.CO(inst_it2_cellmath__62__W0[8]), .S(inst_it2_cellmath__62__W1[8]), .A(inst_it2_cellmath__61[8]), .B(inst_it2_cellmath__60[8]), .CI(inst_it2_cellmath__56[8]));
ADDFX1 inst_fa_1820_10_I2497 (.CO(inst_it2_cellmath__62__W0[9]), .S(inst_it2_cellmath__62__W1[9]), .A(inst_it2_cellmath__61[9]), .B(inst_it2_cellmath__60[9]), .CI(inst_it2_cellmath__56[9]));
ADDFX1 inst_fa_1820_10_I2498 (.CO(inst_it2_cellmath__62__W0[10]), .S(inst_it2_cellmath__62__W1[10]), .A(inst_it2_cellmath__61[10]), .B(inst_it2_cellmath__60[10]), .CI(inst_it2_cellmath__56[10]));
ADDFX1 inst_fa_1820_10_I2499 (.CO(inst_it2_cellmath__62__W0[11]), .S(inst_it2_cellmath__62__W1[11]), .A(inst_it2_cellmath__61[11]), .B(inst_it2_cellmath__60[11]), .CI(inst_it2_cellmath__56[11]));
ADDFX1 inst_fa_1820_10_I2500 (.CO(inst_it2_cellmath__62__W0[12]), .S(inst_it2_cellmath__62__W1[12]), .A(inst_it2_cellmath__61[12]), .B(inst_it2_cellmath__60[12]), .CI(inst_it2_cellmath__56[12]));
ADDFX1 inst_fa_1820_10_I2501 (.CO(inst_it2_cellmath__62__W0[13]), .S(inst_it2_cellmath__62__W1[13]), .A(inst_it2_cellmath__61[13]), .B(inst_it2_cellmath__60[13]), .CI(inst_it2_cellmath__56[13]));
ADDFX1 inst_fa_1820_10_I2502 (.CO(inst_it2_cellmath__62__W0[14]), .S(inst_it2_cellmath__62__W1[14]), .A(inst_it2_cellmath__61[14]), .B(inst_it2_cellmath__60[14]), .CI(inst_it2_cellmath__56[14]));
ADDFX1 inst_fa_1820_10_I2503 (.CO(inst_it2_cellmath__62__W0[15]), .S(inst_it2_cellmath__62__W1[15]), .A(inst_it2_cellmath__61[15]), .B(inst_it2_cellmath__60[15]), .CI(inst_it2_cellmath__56[15]));
ADDFX1 inst_fa_1820_10_I2504 (.CO(inst_it2_cellmath__62__W0[16]), .S(inst_it2_cellmath__62__W1[16]), .A(inst_it2_cellmath__61[16]), .B(inst_it2_cellmath__60[16]), .CI(inst_it2_cellmath__56[16]));
ADDFX1 inst_fa_1820_10_I2505 (.CO(inst_it2_cellmath__62__W0[17]), .S(inst_it2_cellmath__62__W1[17]), .A(inst_it2_cellmath__61[17]), .B(inst_it2_cellmath__60[17]), .CI(inst_it2_cellmath__56[17]));
ADDFX1 inst_fa_1820_10_I2506 (.CO(inst_it2_cellmath__62__W0[18]), .S(inst_it2_cellmath__62__W1[18]), .A(inst_it2_cellmath__61[18]), .B(inst_it2_cellmath__60[18]), .CI(inst_it2_cellmath__56[18]));
ADDFX1 inst_fa_1820_10_I2507 (.CO(inst_it2_cellmath__62__W0[19]), .S(inst_it2_cellmath__62__W1[19]), .A(inst_it2_cellmath__61[19]), .B(inst_it2_cellmath__60[19]), .CI(inst_it2_cellmath__56[19]));
ADDFX1 inst_fa_1820_10_I2508 (.CO(inst_it2_cellmath__62__W0[20]), .S(inst_it2_cellmath__62__W1[20]), .A(inst_it2_cellmath__61[20]), .B(inst_it2_cellmath__60[20]), .CI(inst_it2_cellmath__56[20]));
ADDFX1 inst_fa_1820_10_I2509 (.CO(inst_it2_cellmath__62__W0[21]), .S(inst_it2_cellmath__62__W1[21]), .A(inst_it2_cellmath__61[21]), .B(inst_it2_cellmath__60[21]), .CI(inst_it2_cellmath__56[21]));
ADDFX1 inst_fa_1820_10_I2510 (.CO(inst_it2_cellmath__62__W0[22]), .S(inst_it2_cellmath__62__W1[22]), .A(inst_it2_cellmath__61[22]), .B(inst_it2_cellmath__60[22]), .CI(inst_it2_cellmath__56[22]));
ADDFX1 inst_fa_1820_10_I2511 (.CO(inst_it2_cellmath__62__W0[23]), .S(inst_it2_cellmath__62__W1[23]), .A(inst_it2_cellmath__61[23]), .B(inst_it2_cellmath__60[23]), .CI(inst_it2_cellmath__56[23]));
ADDFX1 inst_fa_1820_10_I2512 (.CO(inst_it2_cellmath__62__W0[24]), .S(inst_it2_cellmath__62__W1[24]), .A(inst_it2_cellmath__61[24]), .B(inst_it2_cellmath__60[24]), .CI(inst_it2_cellmath__56[24]));
XOR3XL inst_fa_1820_10_I2513 (.Y(inst_it2_cellmath__62__W1[25]), .A(inst_it2_cellmath__60[25]), .B(inst_it2_cellmath__61[25]), .C(inst_cellmath__14[2]));
INVXL buf1_A_I9201 (.Y(N28021), .A(inst_cellmath__14[2]));
INVXL buf1_A_I9202 (.Y(inst_cellmath__14[1]), .A(N28021));
ADDHX1 inst_fa_1839_10_I2516 (.CO(inst_cellmath__14[3]), .S(inst_it2_cellmath__63__W1[2]), .A(inst_it2_cellmath__56[2]), .B(inst_it2_cellmath__57[2]));
ADDHX1 inst_fa_1839_10_I2517 (.CO(inst_cellmath__14[4]), .S(inst_it2_cellmath__63__W1[3]), .A(inst_it2_cellmath__62__W1[3]), .B(inst_it2_cellmath__57[3]));
ADDFX1 inst_fa_1839_10_I2518 (.CO(inst_cellmath__14[5]), .S(inst_it2_cellmath__63__W1[4]), .A(inst_it2_cellmath__62__W0[3]), .B(inst_it2_cellmath__62__W1[4]), .CI(inst_it2_cellmath__57[4]));
ADDFX1 inst_fa_1839_10_I2519 (.CO(inst_cellmath__14[6]), .S(inst_it2_cellmath__63__W1[5]), .A(inst_it2_cellmath__62__W0[4]), .B(inst_it2_cellmath__62__W1[5]), .CI(inst_it2_cellmath__57[5]));
ADDFX1 inst_fa_1839_10_I2520 (.CO(inst_cellmath__14[7]), .S(inst_it2_cellmath__63__W1[6]), .A(inst_it2_cellmath__62__W0[5]), .B(inst_it2_cellmath__62__W1[6]), .CI(inst_it2_cellmath__57[6]));
ADDFX1 inst_fa_1839_10_I2521 (.CO(inst_cellmath__14[8]), .S(inst_it2_cellmath__63__W1[7]), .A(inst_it2_cellmath__62__W0[6]), .B(inst_it2_cellmath__62__W1[7]), .CI(inst_it2_cellmath__57[7]));
ADDFX1 inst_fa_1839_10_I2522 (.CO(inst_cellmath__14[9]), .S(inst_it2_cellmath__63__W1[8]), .A(inst_it2_cellmath__62__W0[7]), .B(inst_it2_cellmath__62__W1[8]), .CI(inst_it2_cellmath__57[8]));
ADDFX1 inst_fa_1839_10_I2523 (.CO(inst_cellmath__14[10]), .S(inst_it2_cellmath__63__W1[9]), .A(inst_it2_cellmath__62__W0[8]), .B(inst_it2_cellmath__62__W1[9]), .CI(inst_it2_cellmath__57[9]));
ADDFX1 inst_fa_1839_10_I2524 (.CO(inst_cellmath__14[11]), .S(inst_it2_cellmath__63__W1[10]), .A(inst_it2_cellmath__62__W0[9]), .B(inst_it2_cellmath__62__W1[10]), .CI(inst_it2_cellmath__57[10]));
ADDFX1 inst_fa_1839_10_I2525 (.CO(inst_cellmath__14[12]), .S(inst_it2_cellmath__63__W1[11]), .A(inst_it2_cellmath__62__W0[10]), .B(inst_it2_cellmath__62__W1[11]), .CI(inst_it2_cellmath__57[11]));
ADDFX1 inst_fa_1839_10_I2526 (.CO(inst_cellmath__14[13]), .S(inst_it2_cellmath__63__W1[12]), .A(inst_it2_cellmath__62__W0[11]), .B(inst_it2_cellmath__62__W1[12]), .CI(inst_it2_cellmath__57[12]));
ADDFX1 inst_fa_1839_10_I2527 (.CO(inst_cellmath__14[14]), .S(inst_it2_cellmath__63__W1[13]), .A(inst_it2_cellmath__62__W0[12]), .B(inst_it2_cellmath__62__W1[13]), .CI(inst_it2_cellmath__57[13]));
ADDFX1 inst_fa_1839_10_I2528 (.CO(inst_cellmath__14[15]), .S(inst_it2_cellmath__63__W1[14]), .A(inst_it2_cellmath__62__W0[13]), .B(inst_it2_cellmath__62__W1[14]), .CI(inst_it2_cellmath__57[14]));
ADDFX1 inst_fa_1839_10_I2529 (.CO(inst_cellmath__14[16]), .S(inst_it2_cellmath__63__W1[15]), .A(inst_it2_cellmath__62__W0[14]), .B(inst_it2_cellmath__62__W1[15]), .CI(inst_it2_cellmath__57[15]));
ADDFX1 inst_fa_1839_10_I2530 (.CO(inst_cellmath__14[17]), .S(inst_it2_cellmath__63__W1[16]), .A(inst_it2_cellmath__62__W0[15]), .B(inst_it2_cellmath__62__W1[16]), .CI(inst_it2_cellmath__57[16]));
ADDFX1 inst_fa_1839_10_I2531 (.CO(inst_cellmath__14[18]), .S(inst_it2_cellmath__63__W1[17]), .A(inst_it2_cellmath__62__W0[16]), .B(inst_it2_cellmath__62__W1[17]), .CI(inst_it2_cellmath__57[17]));
ADDFX1 inst_fa_1839_10_I2532 (.CO(inst_cellmath__14[19]), .S(inst_it2_cellmath__63__W1[18]), .A(inst_it2_cellmath__62__W0[17]), .B(inst_it2_cellmath__62__W1[18]), .CI(inst_it2_cellmath__57[18]));
ADDFX1 inst_fa_1839_10_I2533 (.CO(inst_cellmath__14[20]), .S(inst_it2_cellmath__63__W1[19]), .A(inst_it2_cellmath__62__W0[18]), .B(inst_it2_cellmath__62__W1[19]), .CI(inst_it2_cellmath__57[19]));
ADDFX1 inst_fa_1839_10_I2534 (.CO(inst_cellmath__14[21]), .S(inst_it2_cellmath__63__W1[20]), .A(inst_it2_cellmath__62__W0[19]), .B(inst_it2_cellmath__62__W1[20]), .CI(inst_it2_cellmath__57[20]));
ADDFX1 inst_fa_1839_10_I2535 (.CO(inst_cellmath__14[22]), .S(inst_it2_cellmath__63__W1[21]), .A(inst_it2_cellmath__62__W0[20]), .B(inst_it2_cellmath__62__W1[21]), .CI(inst_it2_cellmath__57[21]));
ADDFX1 inst_fa_1839_10_I2536 (.CO(inst_cellmath__14[23]), .S(inst_it2_cellmath__63__W1[22]), .A(inst_it2_cellmath__62__W0[21]), .B(inst_it2_cellmath__62__W1[22]), .CI(inst_it2_cellmath__57[22]));
ADDFX1 inst_fa_1839_10_I2537 (.CO(inst_cellmath__14[24]), .S(inst_it2_cellmath__63__W1[23]), .A(inst_it2_cellmath__62__W0[22]), .B(inst_it2_cellmath__62__W1[23]), .CI(inst_it2_cellmath__57[23]));
ADDFX1 inst_fa_1839_10_I2538 (.CO(inst_cellmath__14[25]), .S(inst_it2_cellmath__63__W1[24]), .A(inst_it2_cellmath__62__W0[23]), .B(inst_it2_cellmath__62__W1[24]), .CI(inst_it2_cellmath__57[24]));
ADDFX1 inst_fa_1839_10_I2539 (.CO(N14981), .S(inst_it2_cellmath__63__W1[25]), .A(inst_it2_cellmath__62__W0[24]), .B(inst_it2_cellmath__62__W1[25]), .CI(inst_it2_cellmath__57[25]));
NAND2XL cynw_cm_float_div_ieee_I2540 (.Y(N1555), .A(inst_it2_lookup1_cellmath__55[1]), .B(inst_cellmath__40[0]));
MX2XL cynw_cm_float_div_ieee_I2541 (.Y(inst_cellmath__40[1]), .A(inst_it2_lookup1_cellmath__55[1]), .B(N1555), .S0(inst_it2_lookup1_cellmath__55[2]));
MX2XL cynw_cm_float_div_ieee_I2543 (.Y(inst_cellmath__40[2]), .A(inst_cellmath__43[0]), .B(inst_cellmath__42[0]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2544 (.Y(inst_cellmath__40[3]), .A(inst_cellmath__43[1]), .B(inst_cellmath__42[1]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2545 (.Y(inst_cellmath__40[4]), .A(inst_cellmath__43[2]), .B(inst_cellmath__42[2]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2546 (.Y(inst_cellmath__40[5]), .A(inst_cellmath__43[3]), .B(inst_cellmath__42[3]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2547 (.Y(inst_cellmath__40[6]), .A(inst_cellmath__43[4]), .B(inst_cellmath__42[4]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2548 (.Y(inst_cellmath__40[7]), .A(inst_cellmath__43[5]), .B(inst_cellmath__42[5]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2549 (.Y(inst_cellmath__40[8]), .A(inst_cellmath__43[6]), .B(inst_cellmath__42[6]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2550 (.Y(inst_cellmath__40[9]), .A(inst_cellmath__43[7]), .B(inst_cellmath__42[7]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2551 (.Y(inst_cellmath__40[10]), .A(inst_cellmath__43[8]), .B(inst_cellmath__42[8]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2552 (.Y(inst_cellmath__40[11]), .A(inst_cellmath__43[9]), .B(inst_cellmath__42[9]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2553 (.Y(inst_cellmath__40[12]), .A(inst_cellmath__43[10]), .B(inst_cellmath__42[10]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2554 (.Y(inst_cellmath__40[13]), .A(inst_cellmath__43[11]), .B(inst_cellmath__42[11]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2555 (.Y(inst_cellmath__40[14]), .A(inst_cellmath__43[12]), .B(inst_cellmath__42[12]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2556 (.Y(inst_cellmath__40[15]), .A(inst_cellmath__43[13]), .B(inst_cellmath__42[13]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2557 (.Y(inst_cellmath__40[16]), .A(inst_cellmath__43[14]), .B(inst_cellmath__42[14]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2558 (.Y(inst_cellmath__40[17]), .A(inst_cellmath__43[15]), .B(inst_cellmath__42[15]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2559 (.Y(inst_cellmath__40[18]), .A(inst_cellmath__43[16]), .B(inst_cellmath__42[16]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2560 (.Y(inst_cellmath__40[19]), .A(inst_cellmath__43[17]), .B(inst_cellmath__42[17]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2561 (.Y(inst_cellmath__40[20]), .A(inst_cellmath__43[18]), .B(inst_cellmath__42[18]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2562 (.Y(inst_cellmath__40[21]), .A(inst_cellmath__43[19]), .B(inst_cellmath__42[19]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2563 (.Y(inst_cellmath__40[22]), .A(inst_cellmath__43[20]), .B(inst_cellmath__42[20]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2564 (.Y(inst_cellmath__40[23]), .A(inst_cellmath__43[21]), .B(inst_cellmath__42[21]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2565 (.Y(inst_cellmath__40[24]), .A(inst_cellmath__43[22]), .B(inst_cellmath__42[22]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2566 (.Y(inst_cellmath__40[25]), .A(inst_cellmath__43[23]), .B(inst_cellmath__42[23]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2567 (.Y(inst_cellmath__40[26]), .A(inst_cellmath__43[24]), .B(inst_cellmath__42[24]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2568 (.Y(inst_cellmath__40[27]), .A(inst_cellmath__43[25]), .B(inst_cellmath__42[25]), .S0(inst_cellmath__14[1]));
MX2XL cynw_cm_float_div_ieee_I2569 (.Y(inst_cellmath__40[28]), .A(inst_cellmath__43[26]), .B(inst_cellmath__42[26]), .S0(inst_cellmath__14[1]));
XOR2XL cynw_cm_float_div_ieee_I2571 (.Y(inst_cellmath__41[1]), .A(inst_cellmath__40[1]), .B(inst_cellmath__41[0]));
OA21X1 inst_cellmath__41_0_I4152 (.Y(N15334), .A0(inst_cellmath__40[0]), .A1(inst_cellmath__40[1]), .B0(inst_cellmath__14[2]));
MX2XL inst_cellmath__41_0_I2576 (.Y(inst_cellmath__41[2]), .A(inst_cellmath__43[0]), .B(inst_cellmath__42[0]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2577 (.Y(inst_cellmath__41[3]), .A(inst_cellmath__43[1]), .B(inst_cellmath__42[1]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2578 (.Y(inst_cellmath__41[4]), .A(inst_cellmath__43[2]), .B(inst_cellmath__42[2]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2579 (.Y(inst_cellmath__41[5]), .A(inst_cellmath__43[3]), .B(inst_cellmath__42[3]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2580 (.Y(inst_cellmath__41[6]), .A(inst_cellmath__43[4]), .B(inst_cellmath__42[4]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2581 (.Y(inst_cellmath__41[7]), .A(inst_cellmath__43[5]), .B(inst_cellmath__42[5]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2582 (.Y(inst_cellmath__41[8]), .A(inst_cellmath__43[6]), .B(inst_cellmath__42[6]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2583 (.Y(inst_cellmath__41[9]), .A(inst_cellmath__43[7]), .B(inst_cellmath__42[7]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2584 (.Y(inst_cellmath__41[10]), .A(inst_cellmath__43[8]), .B(inst_cellmath__42[8]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2585 (.Y(inst_cellmath__41[11]), .A(inst_cellmath__43[9]), .B(inst_cellmath__42[9]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2586 (.Y(inst_cellmath__41[12]), .A(inst_cellmath__43[10]), .B(inst_cellmath__42[10]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2587 (.Y(inst_cellmath__41[13]), .A(inst_cellmath__43[11]), .B(inst_cellmath__42[11]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2588 (.Y(inst_cellmath__41[14]), .A(inst_cellmath__43[12]), .B(inst_cellmath__42[12]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2589 (.Y(inst_cellmath__41[15]), .A(inst_cellmath__43[13]), .B(inst_cellmath__42[13]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2590 (.Y(inst_cellmath__41[16]), .A(inst_cellmath__43[14]), .B(inst_cellmath__42[14]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2591 (.Y(inst_cellmath__41[17]), .A(inst_cellmath__43[15]), .B(inst_cellmath__42[15]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2592 (.Y(inst_cellmath__41[18]), .A(inst_cellmath__43[16]), .B(inst_cellmath__42[16]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2593 (.Y(inst_cellmath__41[19]), .A(inst_cellmath__43[17]), .B(inst_cellmath__42[17]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2594 (.Y(inst_cellmath__41[20]), .A(inst_cellmath__43[18]), .B(inst_cellmath__42[18]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2595 (.Y(inst_cellmath__41[21]), .A(inst_cellmath__43[19]), .B(inst_cellmath__42[19]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2596 (.Y(inst_cellmath__41[22]), .A(inst_cellmath__43[20]), .B(inst_cellmath__42[20]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2597 (.Y(inst_cellmath__41[23]), .A(inst_cellmath__43[21]), .B(inst_cellmath__42[21]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2598 (.Y(inst_cellmath__41[24]), .A(inst_cellmath__43[22]), .B(inst_cellmath__42[22]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2599 (.Y(inst_cellmath__41[25]), .A(inst_cellmath__43[23]), .B(inst_cellmath__42[23]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2600 (.Y(inst_cellmath__41[26]), .A(inst_cellmath__43[24]), .B(inst_cellmath__42[24]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2601 (.Y(inst_cellmath__41[27]), .A(inst_cellmath__43[25]), .B(inst_cellmath__42[25]), .S0(N15334));
MX2XL inst_cellmath__41_0_I2602 (.Y(inst_cellmath__41[28]), .A(inst_cellmath__43[26]), .B(inst_cellmath__42[26]), .S0(N15334));
INVXL inst_cellmath__67_0_I2603 (.Y(N15444), .A(inst_cellmath__9[23]));
INVXL inst_cellmath__67_0_I2604 (.Y(N15413), .A(inst_cellmath__9[24]));
INVXL inst_cellmath__67_0_I2605 (.Y(N15436), .A(inst_cellmath__9[25]));
INVXL inst_cellmath__67_0_I2606 (.Y(N15406), .A(inst_cellmath__9[26]));
INVXL inst_cellmath__67_0_I2607 (.Y(N15431), .A(inst_cellmath__9[27]));
INVXL inst_cellmath__67_0_I2608 (.Y(N15401), .A(inst_cellmath__9[28]));
INVXL inst_cellmath__67_0_I2609 (.Y(N15423), .A(inst_cellmath__9[29]));
INVXL inst_cellmath__67_0_I2610 (.Y(N15432), .A(inst_cellmath__8[24]));
XNOR2X1 inst_cellmath__67_0_I2611 (.Y(N15424), .A(inst_cellmath__8[24]), .B(N15436));
OR2XL inst_cellmath__67_0_I2612 (.Y(N15435), .A(inst_cellmath__8[24]), .B(N15436));
XNOR2X1 inst_cellmath__67_0_I2613 (.Y(N15417), .A(inst_cellmath__8[26]), .B(N15406));
OR2XL inst_cellmath__67_0_I2614 (.Y(N15430), .A(inst_cellmath__8[26]), .B(N15406));
XNOR2X1 inst_cellmath__67_0_I2615 (.Y(N15411), .A(inst_cellmath__8[27]), .B(N15431));
OR2XL inst_cellmath__67_0_I2616 (.Y(N15421), .A(inst_cellmath__8[27]), .B(N15431));
XNOR2X1 inst_cellmath__67_0_I2617 (.Y(N15403), .A(inst_cellmath__8[28]), .B(N15401));
OR2XL inst_cellmath__67_0_I2618 (.Y(N15415), .A(inst_cellmath__8[28]), .B(N15401));
XNOR2X1 inst_cellmath__67_0_I2619 (.Y(N15398), .A(inst_cellmath__8[29]), .B(N15423));
OR2XL inst_cellmath__67_0_I2620 (.Y(N15409), .A(inst_cellmath__8[29]), .B(N15423));
XNOR2X1 inst_cellmath__67_0_I2621 (.Y(N15443), .A(inst_cellmath__8[30]), .B(inst_cellmath__9[30]));
XNOR2X1 inst_cellmath__67_0_I2622 (.Y(inst_cellmath__67[0]), .A(N15444), .B(inst_cellmath__8[23]));
OR2XL inst_cellmath__67_0_I2623 (.Y(N15426), .A(N15444), .B(inst_cellmath__8[23]));
ADDFX1 inst_cellmath__67_0_I2624 (.CO(N15418), .S(inst_cellmath__67[1]), .A(N15432), .B(N15413), .CI(N15426));
ADDFX1 inst_cellmath__67_0_I2625 (.CO(N15440), .S(inst_cellmath__67[2]), .A(N15424), .B(inst_cellmath__8[25]), .CI(N15418));
ADDFX1 inst_cellmath__67_0_I2626 (.CO(N15412), .S(inst_cellmath__67[3]), .A(N15417), .B(N15435), .CI(N15440));
ADDFX1 inst_cellmath__67_0_I2627 (.CO(N15434), .S(inst_cellmath__67[4]), .A(N15411), .B(N15430), .CI(N15412));
ADDFX1 inst_cellmath__67_0_I2628 (.CO(N15404), .S(inst_cellmath__67[5]), .A(N15403), .B(N15421), .CI(N15434));
ADDFX1 inst_cellmath__67_0_I2629 (.CO(N15429), .S(inst_cellmath__67[6]), .A(N15398), .B(N15415), .CI(N15404));
ADDFX1 inst_cellmath__67_0_I2630 (.CO(N15400), .S(inst_cellmath__67[7]), .A(N15443), .B(N15409), .CI(N15429));
INVXL inst_cellmath__68_0_I2638 (.Y(N15503), .A(inst_cellmath__9[30]));
INVXL inst_cellmath__68_0_I2639 (.Y(N15497), .A(inst_cellmath__8[30]));
ADDHX1 inst_cellmath__68_0_I2640 (.CO(N15504), .S(inst_cellmath__68[0]), .A(inst_cellmath__8[23]), .B(N15444));
ADDFX1 inst_cellmath__68_0_I2641 (.CO(N15495), .S(inst_cellmath__68[1]), .A(N15413), .B(inst_cellmath__8[24]), .CI(N15504));
ADDFX1 inst_cellmath__68_0_I2642 (.CO(N15518), .S(inst_cellmath__68[2]), .A(N15436), .B(inst_cellmath__8[25]), .CI(N15495));
ADDFX1 inst_cellmath__68_0_I2643 (.CO(N15491), .S(inst_cellmath__68[3]), .A(N15406), .B(inst_cellmath__8[26]), .CI(N15518));
ADDFX1 inst_cellmath__68_0_I2644 (.CO(N15511), .S(inst_cellmath__68[4]), .A(N15431), .B(inst_cellmath__8[27]), .CI(N15491));
ADDFX1 inst_cellmath__68_0_I2645 (.CO(N15486), .S(inst_cellmath__68[5]), .A(N15401), .B(inst_cellmath__8[28]), .CI(N15511));
ADDFX1 inst_cellmath__68_0_I2646 (.CO(N15506), .S(inst_cellmath__68[6]), .A(N15423), .B(inst_cellmath__8[29]), .CI(N15486));
ADDFX1 inst_cellmath__68_0_I2647 (.CO(N15523), .S(inst_cellmath__68[7]), .A(N15503), .B(N15497), .CI(N15506));
XNOR2X1 inst_cellmath__68_0_I2648 (.Y(inst_cellmath__68[8]), .A(inst_cellmath__8[30]), .B(N15523));
NOR2XL inst_cellmath__68_0_I2649 (.Y(inst_cellmath__68[9]), .A(inst_cellmath__8[30]), .B(N15523));
AND2XL inst_cellmath__69__82__I2650 (.Y(N15554), .A(inst_cellmath__68[0]), .B(inst_cellmath__68[1]));
NAND3XL inst_cellmath__69__82__I2651 (.Y(N15560), .A(inst_cellmath__68[3]), .B(inst_cellmath__68[4]), .C(inst_cellmath__68[7]));
NAND4XL inst_cellmath__69__82__I2652 (.Y(N15552), .A(inst_cellmath__68[2]), .B(N15554), .C(inst_cellmath__68[6]), .D(inst_cellmath__68[5]));
NOR2XL inst_cellmath__69__82__I2653 (.Y(N1675), .A(N15560), .B(N15552));
NOR2XL andori2bb1_A_I4163 (.Y(N18408), .A(inst_cellmath__68[8]), .B(N1675));
NOR2XL andori2bb1_A_I4164 (.Y(inst_cellmath__69), .A(N18408), .B(inst_cellmath__68[9]));
NOR2XL inst_cellmath__70__83__I2656 (.Y(N15585), .A(inst_cellmath__68[0]), .B(inst_cellmath__68[1]));
NOR2XL inst_cellmath__70__83__I2657 (.Y(N15589), .A(inst_cellmath__68[2]), .B(inst_cellmath__68[3]));
NOR2XL inst_cellmath__70__83__I2658 (.Y(N15582), .A(inst_cellmath__68[6]), .B(inst_cellmath__68[7]));
INVXL inst_cellmath__70__83__I2659 (.Y(N15583), .A(inst_cellmath__68[8]));
NOR4BBX1 inst_cellmath__70__83__I4159 (.Y(N15579), .AN(N15583), .BN(N15585), .C(inst_cellmath__68[4]), .D(inst_cellmath__68[5]));
NAND3XL inst_cellmath__70__83__I2663 (.Y(N1677), .A(N15589), .B(N15582), .C(N15579));
NAND2BXL cynw_cm_float_div_ieee_I2664 (.Y(inst_cellmath__70), .AN(inst_cellmath__68[9]), .B(N1677));
NAND3BXL inst_cellmath__71_0_I2665 (.Y(N15608), .AN(inst_cellmath__68[9]), .B(inst_cellmath__68[0]), .C(inst_cellmath__68[1]));
AND4XL inst_cellmath__71_0_I9190 (.Y(N15618), .A(inst_cellmath__68[2]), .B(inst_cellmath__68[3]), .C(inst_cellmath__68[4]), .D(inst_cellmath__68[6]));
NAND3BXL inst_cellmath__71_0_I2669 (.Y(N15605), .AN(inst_cellmath__68[8]), .B(inst_cellmath__68[7]), .C(N15618));
NOR3BXL inst_cellmath__71_0_I2670 (.Y(inst_cellmath__71), .AN(inst_cellmath__68[5]), .B(N15608), .C(N15605));
NOR2XL inst_cellmath__72_0_I2672 (.Y(N15631), .A(inst_cellmath__68[4]), .B(inst_cellmath__68[6]));
INVXL inst_cellmath__72_0_I2673 (.Y(N15640), .A(inst_cellmath__68[7]));
NAND4XL inst_cellmath__72_0_I2675 (.Y(N15636), .A(N15640), .B(N15583), .C(N15589), .D(N15631));
NOR4BX1 inst_cellmath__72_0_I2676 (.Y(inst_cellmath__72), .AN(inst_cellmath__68[0]), .B(inst_cellmath__68[1]), .C(inst_cellmath__68[5]), .D(N15636));
NOR2BX1 cynw_cm_float_div_ieee_I2677 (.Y(inst_cellmath__73), .AN(inst_cellmath__69), .B(inst_cellmath__71));
OR2XL cynw_cm_float_div_ieee_I2678 (.Y(inst_cellmath__74), .A(inst_cellmath__72), .B(inst_cellmath__70));
NAND2XL inst_cellmath__75_0_I2679 (.Y(N15660), .A(inst_cellmath__8[30]), .B(inst_cellmath__8[24]));
NAND2XL inst_cellmath__75_0_I2680 (.Y(N15663), .A(inst_cellmath__8[29]), .B(inst_cellmath__8[25]));
NAND2XL inst_cellmath__75_0_I2681 (.Y(N15666), .A(inst_cellmath__8[27]), .B(inst_cellmath__8[28]));
NAND2XL inst_cellmath__75_0_I2682 (.Y(N15656), .A(inst_cellmath__8[26]), .B(inst_cellmath__8[23]));
NOR4X1 inst_cellmath__75_0_I2683 (.Y(inst_cellmath__75), .A(N15663), .B(N15660), .C(N15666), .D(N15656));
NAND2XL inst_cellmath__76_0_I2684 (.Y(N15679), .A(inst_cellmath__9[25]), .B(inst_cellmath__9[27]));
AND4XL inst_cellmath__76_0_I9191 (.Y(N15681), .A(inst_cellmath__9[26]), .B(inst_cellmath__9[24]), .C(inst_cellmath__9[29]), .D(inst_cellmath__9[30]));
NAND3XL hyperpropagate_4_1_A_I4165 (.Y(N18417), .A(inst_cellmath__9[28]), .B(inst_cellmath__9[23]), .C(N15681));
NOR2XL hyperpropagate_4_1_A_I4166 (.Y(inst_cellmath__76), .A(N15679), .B(N18417));
NOR2XL inst_cellmath__77_0_I2691 (.Y(N15722), .A(inst_cellmath__8[1]), .B(inst_cellmath__8[2]));
NOR2XL inst_cellmath__77_0_I2692 (.Y(N15732), .A(inst_cellmath__8[18]), .B(inst_cellmath__8[16]));
NOR2XL inst_cellmath__77_0_I2693 (.Y(N15699), .A(inst_cellmath__8[14]), .B(inst_cellmath__8[12]));
NOR2XL inst_cellmath__77_0_I2696 (.Y(N15726), .A(inst_cellmath__8[19]), .B(inst_cellmath__8[17]));
NOR2XL inst_cellmath__77_0_I2697 (.Y(N15736), .A(inst_cellmath__8[15]), .B(inst_cellmath__8[13]));
NOR2XL inst_cellmath__77_0_I2698 (.Y(N15702), .A(inst_cellmath__8[11]), .B(inst_cellmath__8[9]));
NOR2XL inst_cellmath__77_0_I2699 (.Y(N15711), .A(inst_cellmath__8[7]), .B(inst_cellmath__8[5]));
NOR2XL inst_cellmath__77_0_I2700 (.Y(N15720), .A(inst_cellmath__8[3]), .B(inst_cellmath__8[0]));
NOR2XL inst_cellmath__77_0_I2701 (.Y(N15730), .A(inst_cellmath__8[22]), .B(inst_cellmath__8[21]));
OR4X1 inst_cellmath__77_0_I9192 (.Y(N15724), .A(inst_cellmath__8[4]), .B(inst_cellmath__8[8]), .C(inst_cellmath__8[6]), .D(inst_cellmath__8[10]));
AND4XL inst_cellmath__77_0_I2703 (.Y(N15728), .A(N15736), .B(N15711), .C(N15702), .D(N15726));
NAND3XL inst_cellmath__77_0_I2704 (.Y(N15710), .A(N15722), .B(N15720), .C(N15730));
NAND3XL inst_cellmath__77_0_I2706 (.Y(N15733), .A(N15732), .B(N15699), .C(N15728));
OR4X1 inst_cellmath__77_0_I9193 (.Y(inst_cellmath__77), .A(inst_cellmath__8[20]), .B(N15710), .C(N15724), .D(N15733));
NOR2XL inst_cellmath__78_0_I2709 (.Y(N15782), .A(inst_cellmath__9[1]), .B(inst_cellmath__9[2]));
NOR2XL inst_cellmath__78_0_I2710 (.Y(N15792), .A(inst_cellmath__9[18]), .B(inst_cellmath__9[16]));
NOR2XL inst_cellmath__78_0_I2711 (.Y(N15758), .A(inst_cellmath__9[14]), .B(inst_cellmath__9[12]));
NOR2XL inst_cellmath__78_0_I2714 (.Y(N15786), .A(inst_cellmath__9[19]), .B(inst_cellmath__9[17]));
NOR2XL inst_cellmath__78_0_I2715 (.Y(N15795), .A(inst_cellmath__9[15]), .B(inst_cellmath__9[13]));
NOR2XL inst_cellmath__78_0_I2716 (.Y(N15762), .A(inst_cellmath__9[11]), .B(inst_cellmath__9[9]));
NOR2XL inst_cellmath__78_0_I2717 (.Y(N15770), .A(inst_cellmath__9[7]), .B(inst_cellmath__9[5]));
NOR2XL inst_cellmath__78_0_I2718 (.Y(N15779), .A(inst_cellmath__9[3]), .B(inst_cellmath__9[0]));
NOR2XL inst_cellmath__78_0_I2719 (.Y(N15790), .A(inst_cellmath__9[20]), .B(inst_it2_lookup1_cellmath__53[1]));
OR4X1 inst_cellmath__78_0_I9194 (.Y(N15784), .A(inst_cellmath__9[4]), .B(inst_cellmath__9[8]), .C(inst_cellmath__9[6]), .D(inst_cellmath__9[10]));
AND4XL inst_cellmath__78_0_I2721 (.Y(N15788), .A(N15795), .B(N15770), .C(N15762), .D(N15786));
NAND3XL inst_cellmath__78_0_I2722 (.Y(N15759), .A(N15779), .B(N15782), .C(N15790));
NAND3XL inst_cellmath__78_0_I2724 (.Y(N15780), .A(N15792), .B(N15758), .C(N15788));
OR4X1 inst_cellmath__78_0_I9195 (.Y(inst_cellmath__78), .A(inst_it2_lookup1_cellmath__53[0]), .B(N15759), .C(N15784), .D(N15780));
AND2XL cynw_cm_float_div_ieee_I2727 (.Y(inst_cellmath__79), .A(inst_cellmath__75), .B(inst_cellmath__77));
AND2XL cynw_cm_float_div_ieee_I2728 (.Y(inst_cellmath__80), .A(inst_cellmath__76), .B(inst_cellmath__78));
NOR2BX1 cynw_cm_float_div_ieee_I2729 (.Y(inst_cellmath__83), .AN(inst_cellmath__75), .B(inst_cellmath__77));
NOR2BX1 cynw_cm_float_div_ieee_I2730 (.Y(inst_cellmath__84), .AN(inst_cellmath__76), .B(inst_cellmath__78));
NOR2XL inst_cellmath__85__85__I2731 (.Y(N15834), .A(inst_cellmath__8[30]), .B(inst_cellmath__8[24]));
NOR2XL inst_cellmath__85__85__I2732 (.Y(N15837), .A(inst_cellmath__8[29]), .B(inst_cellmath__8[25]));
NOR2XL inst_cellmath__85__85__I2733 (.Y(N15840), .A(inst_cellmath__8[27]), .B(inst_cellmath__8[28]));
NOR2XL inst_cellmath__85__85__I2734 (.Y(N15830), .A(inst_cellmath__8[26]), .B(inst_cellmath__8[23]));
AND4XL inst_cellmath__85__85__I2735 (.Y(inst_cellmath__85), .A(N15834), .B(N15837), .C(N15840), .D(N15830));
NOR2XL inst_cellmath__86__86__I2736 (.Y(N15852), .A(inst_cellmath__9[25]), .B(inst_cellmath__9[27]));
NOR2XL inst_cellmath__86__86__I2737 (.Y(N15855), .A(inst_cellmath__9[28]), .B(inst_cellmath__9[23]));
NOR2XL inst_cellmath__86__86__I2738 (.Y(N15858), .A(inst_cellmath__9[29]), .B(inst_cellmath__9[24]));
NOR2XL inst_cellmath__86__86__I2739 (.Y(N15848), .A(inst_cellmath__9[30]), .B(inst_cellmath__9[26]));
AND4XL inst_cellmath__86__86__I2740 (.Y(inst_cellmath__86), .A(N15852), .B(N15858), .C(N15855), .D(N15848));
AND2XL cynw_cm_float_div_ieee_I2741 (.Y(N1678), .A(inst_cellmath__83), .B(inst_cellmath__84));
AND2XL cynw_cm_float_div_ieee_I2742 (.Y(N1679), .A(inst_cellmath__86), .B(inst_cellmath__85));
OR4X1 cynw_cm_float_div_ieee_I2743 (.Y(inst_cellmath__87), .A(N1679), .B(inst_cellmath__79), .C(inst_cellmath__80), .D(N1678));
OR2XL cynw_cm_float_div_ieee_I2744 (.Y(inst_cellmath__88), .A(inst_cellmath__86), .B(inst_cellmath__83));
OR2XL cynw_cm_float_div_ieee_I2745 (.Y(inst_cellmath__89), .A(inst_cellmath__85), .B(inst_cellmath__84));
XOR2XL cynw_cm_float_div_ieee_I2746 (.Y(inst_cellmath__91), .A(inst_cellmath__9[31]), .B(inst_cellmath__8[31]));
OR2XL cynw_cm_float_div_ieee_I2747 (.Y(N1680), .A(inst_cellmath__91), .B(inst_cellmath__87));
NOR2BX1 inst_cellmath__90_2WWMM_I2748 (.Y(N15943), .AN(inst_cellmath__80), .B(inst_cellmath__79));
NOR2XL inst_cellmath__90_2WWMM_I2749 (.Y(N15898), .A(inst_cellmath__80), .B(inst_cellmath__79));
AOI22XL inst_cellmath__90_2WWMM_I2750 (.Y(N15964), .A0(inst_cellmath__8[31]), .A1(inst_cellmath__79), .B0(N15943), .B1(inst_cellmath__9[31]));
AO22XL inst_cellmath__90_2WWMM_I2751 (.Y(N1751), .A0(inst_cellmath__79), .A1(inst_cellmath__8[0]), .B0(N15943), .B1(inst_cellmath__9[0]));
AO22XL inst_cellmath__90_2WWMM_I2752 (.Y(N1752), .A0(inst_cellmath__79), .A1(inst_cellmath__8[1]), .B0(N15943), .B1(inst_cellmath__9[1]));
AO22XL inst_cellmath__90_2WWMM_I2753 (.Y(N1753), .A0(inst_cellmath__79), .A1(inst_cellmath__8[2]), .B0(N15943), .B1(inst_cellmath__9[2]));
AO22XL inst_cellmath__90_2WWMM_I2754 (.Y(N1754), .A0(inst_cellmath__79), .A1(inst_cellmath__8[3]), .B0(N15943), .B1(inst_cellmath__9[3]));
AO22XL inst_cellmath__90_2WWMM_I2755 (.Y(N1755), .A0(inst_cellmath__79), .A1(inst_cellmath__8[4]), .B0(N15943), .B1(inst_cellmath__9[4]));
AO22XL inst_cellmath__90_2WWMM_I2756 (.Y(N1756), .A0(inst_cellmath__79), .A1(inst_cellmath__8[5]), .B0(N15943), .B1(inst_cellmath__9[5]));
AO22XL inst_cellmath__90_2WWMM_I2757 (.Y(N1757), .A0(inst_cellmath__79), .A1(inst_cellmath__8[6]), .B0(N15943), .B1(inst_cellmath__9[6]));
AO22XL inst_cellmath__90_2WWMM_I2758 (.Y(N1758), .A0(inst_cellmath__79), .A1(inst_cellmath__8[7]), .B0(N15943), .B1(inst_cellmath__9[7]));
AO22XL inst_cellmath__90_2WWMM_I2759 (.Y(N1759), .A0(inst_cellmath__79), .A1(inst_cellmath__8[8]), .B0(N15943), .B1(inst_cellmath__9[8]));
AO22XL inst_cellmath__90_2WWMM_I2760 (.Y(N1760), .A0(inst_cellmath__79), .A1(inst_cellmath__8[9]), .B0(N15943), .B1(inst_cellmath__9[9]));
AO22XL inst_cellmath__90_2WWMM_I2761 (.Y(N1761), .A0(inst_cellmath__79), .A1(inst_cellmath__8[10]), .B0(N15943), .B1(inst_cellmath__9[10]));
AO22XL inst_cellmath__90_2WWMM_I2762 (.Y(N1762), .A0(inst_cellmath__79), .A1(inst_cellmath__8[11]), .B0(N15943), .B1(inst_cellmath__9[11]));
AO22XL inst_cellmath__90_2WWMM_I2763 (.Y(N1763), .A0(inst_cellmath__79), .A1(inst_cellmath__8[12]), .B0(N15943), .B1(inst_cellmath__9[12]));
AO22XL inst_cellmath__90_2WWMM_I2764 (.Y(N1764), .A0(inst_cellmath__79), .A1(inst_cellmath__8[13]), .B0(N15943), .B1(inst_cellmath__9[13]));
AO22XL inst_cellmath__90_2WWMM_I2765 (.Y(N1765), .A0(inst_cellmath__79), .A1(inst_cellmath__8[14]), .B0(N15943), .B1(inst_cellmath__9[14]));
AO22XL inst_cellmath__90_2WWMM_I2766 (.Y(N1766), .A0(inst_cellmath__79), .A1(inst_cellmath__8[15]), .B0(N15943), .B1(inst_cellmath__9[15]));
AO22XL inst_cellmath__90_2WWMM_I2767 (.Y(N1767), .A0(inst_cellmath__79), .A1(inst_cellmath__8[16]), .B0(N15943), .B1(inst_cellmath__9[16]));
AO22XL inst_cellmath__90_2WWMM_I2768 (.Y(N1768), .A0(inst_cellmath__79), .A1(inst_cellmath__8[17]), .B0(N15943), .B1(inst_cellmath__9[17]));
AO22XL inst_cellmath__90_2WWMM_I2769 (.Y(N1769), .A0(inst_cellmath__79), .A1(inst_cellmath__8[18]), .B0(N15943), .B1(inst_cellmath__9[18]));
AO22XL inst_cellmath__90_2WWMM_I2770 (.Y(N1770), .A0(inst_cellmath__79), .A1(inst_cellmath__8[19]), .B0(N15943), .B1(inst_cellmath__9[19]));
AO22XL inst_cellmath__90_2WWMM_I2771 (.Y(N1771), .A0(inst_cellmath__79), .A1(inst_cellmath__8[20]), .B0(N15943), .B1(inst_cellmath__9[20]));
AO22XL inst_cellmath__90_2WWMM_I2772 (.Y(N1772), .A0(inst_cellmath__79), .A1(inst_cellmath__8[21]), .B0(N15943), .B1(inst_it2_lookup1_cellmath__53[0]));
OAI2BB1X1 inst_cellmath__90_2WWMM_I2773 (.Y(N1750), .A0N(N15898), .A1N(N1680), .B0(N15964));
NAND3XL hyperpropagate_4_1_A_I9203 (.Y(N28027), .A(inst_cellmath__12[0]), .B(inst_cellmath__12[2]), .C(inst_cellmath__12[1]));
NOR2XL hyperpropagate_4_1_A_I9204 (.Y(inst_cellmath__96), .A(inst_cellmath__12[3]), .B(N28027));
DFFQXL inst_cellmath__98_0_I318 (.Q(inst_cellmath__113[31]), .D(N1750), .CK(clk));
DFFQXL inst_cellmath__100_0_I319 (.Q(inst_cellmath__100), .D(inst_cellmath__87), .CK(clk));
DFFQXL inst_cellmath__101_0_I320 (.Q(inst_cellmath__101), .D(inst_cellmath__88), .CK(clk));
DFFQXL inst_cellmath__102_0_I321 (.Q(inst_cellmath__102), .D(inst_cellmath__89), .CK(clk));
DFFQXL inst_cellmath__103_0_I322 (.Q(inst_cellmath__103), .D(inst_cellmath__69), .CK(clk));
DFFQXL inst_cellmath__104_0_I323 (.Q(inst_cellmath__104), .D(inst_cellmath__73), .CK(clk));
DFFQXL inst_cellmath__105_0_I324 (.Q(inst_cellmath__105), .D(inst_cellmath__70), .CK(clk));
DFFQXL inst_cellmath__106_0_I325 (.Q(inst_cellmath__106), .D(inst_cellmath__74), .CK(clk));
DFFQXL inst_cellmath__110_0_0__I326 (.Q(inst_cellmath__110[0]), .D(inst_cellmath__67[0]), .CK(clk));
DFFQXL inst_cellmath__110_0_1__I327 (.Q(inst_cellmath__110[1]), .D(inst_cellmath__67[1]), .CK(clk));
DFFQXL inst_cellmath__110_0_2__I328 (.Q(inst_cellmath__110[2]), .D(inst_cellmath__67[2]), .CK(clk));
DFFQXL inst_cellmath__110_0_3__I329 (.Q(inst_cellmath__110[3]), .D(inst_cellmath__67[3]), .CK(clk));
DFFQXL inst_cellmath__110_0_4__I330 (.Q(inst_cellmath__110[4]), .D(inst_cellmath__67[4]), .CK(clk));
DFFQXL inst_cellmath__110_0_5__I331 (.Q(inst_cellmath__110[5]), .D(inst_cellmath__67[5]), .CK(clk));
DFFQXL inst_cellmath__110_0_6__I332 (.Q(inst_cellmath__110[6]), .D(inst_cellmath__67[6]), .CK(clk));
DFFQXL inst_cellmath__110_0_7__I333 (.Q(inst_cellmath__110[7]), .D(inst_cellmath__67[7]), .CK(clk));
DFFQXL inst_cellmath__111_0_0__I334 (.Q(inst_cellmath__111[0]), .D(inst_cellmath__68[0]), .CK(clk));
DFFQXL inst_cellmath__111_0_1__I335 (.Q(inst_cellmath__111[1]), .D(inst_cellmath__68[1]), .CK(clk));
DFFQXL inst_cellmath__111_0_2__I336 (.Q(inst_cellmath__111[2]), .D(inst_cellmath__68[2]), .CK(clk));
DFFQXL inst_cellmath__111_0_3__I337 (.Q(inst_cellmath__111[3]), .D(inst_cellmath__68[3]), .CK(clk));
DFFQXL inst_cellmath__111_0_4__I338 (.Q(inst_cellmath__111[4]), .D(inst_cellmath__68[4]), .CK(clk));
DFFQXL inst_cellmath__111_0_5__I339 (.Q(inst_cellmath__111[5]), .D(inst_cellmath__68[5]), .CK(clk));
DFFQXL inst_cellmath__111_0_6__I340 (.Q(inst_cellmath__111[6]), .D(inst_cellmath__68[6]), .CK(clk));
DFFQXL inst_cellmath__111_0_7__I341 (.Q(inst_cellmath__111[7]), .D(inst_cellmath__68[7]), .CK(clk));
DFFQXL inst_cellmath__109_0_I342 (.Q(inst_cellmath__109), .D(inst_cellmath__96), .CK(clk));
INVXL cynw_cm_float_div_ieee_I362 (.Y(N4587), .A(inst_cellmath__109));
INVX2 cynw_cm_float_div_ieee_I369 (.Y(N4594), .A(N4587));
NOR2XL inst_cellmath__135_0_I2778 (.Y(N16019), .A(inst_cellmath__103), .B(inst_cellmath__101));
INVXL inst_cellmath__135_0_I2779 (.Y(N16014), .A(inst_cellmath__100));
NOR3BXL inst_cellmath__135_0_I2780 (.Y(N16016), .AN(N16014), .B(inst_cellmath__105), .C(inst_cellmath__102));
NAND2XL inst_cellmath__135_0_I2781 (.Y(inst_cellmath__135), .A(N16019), .B(N16016));
NOR2XL inst_cellmath__136_0_I2785 (.Y(N16033), .A(inst_cellmath__102), .B(inst_cellmath__101));
NOR3BXL inst_cellmath__136_0_I4157 (.Y(N16030), .AN(N16014), .B(inst_cellmath__106), .C(inst_cellmath__104));
NAND2XL inst_cellmath__136_0_I2788 (.Y(inst_cellmath__136), .A(N16033), .B(N16030));
MX2XL cynw_cm_float_div_ieee_I2789 (.Y(inst_cellmath__137), .A(inst_cellmath__135), .B(inst_cellmath__136), .S0(inst_cellmath__122));
NOR2XL inst_cellmath__113__113__I2790 (.Y(N16067), .A(inst_cellmath__122), .B(inst_cellmath__137));
NOR2BX1 inst_cellmath__113__113__I2791 (.Y(N16083), .AN(inst_cellmath__122), .B(inst_cellmath__137));
AOI22XL inst_cellmath__113__113__I2792 (.Y(N16052), .A0(inst_cellmath__110[0]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[0]));
AOI22XL inst_cellmath__113__113__I2793 (.Y(N16070), .A0(inst_cellmath__110[1]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[1]));
AOI22XL inst_cellmath__113__113__I2794 (.Y(N16086), .A0(inst_cellmath__110[2]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[2]));
AOI22XL inst_cellmath__113__113__I2795 (.Y(N16064), .A0(inst_cellmath__110[3]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[3]));
AOI22XL inst_cellmath__113__113__I2796 (.Y(N16080), .A0(inst_cellmath__110[4]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[4]));
AOI22XL inst_cellmath__113__113__I2797 (.Y(N16059), .A0(inst_cellmath__110[5]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[5]));
AOI22XL inst_cellmath__113__113__I2798 (.Y(N16076), .A0(inst_cellmath__110[6]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[6]));
AOI22XL inst_cellmath__113__113__I2799 (.Y(N16055), .A0(inst_cellmath__110[7]), .A1(N16083), .B0(N16067), .B1(inst_cellmath__111[7]));
OAI31X1 inst_cellmath__113__113__I4158 (.Y(N16051), .A0(inst_cellmath__103), .A1(inst_cellmath__101), .A2(inst_cellmath__100), .B0(inst_cellmath__137));
NAND2XL inst_cellmath__113__113__I2801 (.Y(inst_cellmath__113[23]), .A(N16051), .B(N16052));
NAND2XL inst_cellmath__113__113__I2802 (.Y(inst_cellmath__113[24]), .A(N16051), .B(N16070));
NAND2XL inst_cellmath__113__113__I2803 (.Y(inst_cellmath__113[25]), .A(N16051), .B(N16086));
NAND2XL inst_cellmath__113__113__I2804 (.Y(inst_cellmath__113[26]), .A(N16051), .B(N16064));
NAND2XL inst_cellmath__113__113__I2805 (.Y(inst_cellmath__113[27]), .A(N16051), .B(N16080));
NAND2XL inst_cellmath__113__113__I2806 (.Y(inst_cellmath__113[28]), .A(N16051), .B(N16059));
NAND2XL inst_cellmath__113__113__I2807 (.Y(inst_cellmath__113[29]), .A(N16051), .B(N16076));
NAND2XL inst_cellmath__113__113__I2808 (.Y(inst_cellmath__113[30]), .A(N16051), .B(N16055));
AND2XL inst_cellmath__113__115__U_2WWMM_I2809 (.Y(N16178), .A(inst_cellmath__100), .B(inst_cellmath__137));
INVXL inst_cellmath__113__115__U_2WWMM_I2810 (.Y(N16122), .A(inst_cellmath__137));
AO22XL inst_cellmath__113__115__U_2WWMM_I2811 (.Y(inst_cellmath__113[0]), .A0(N16178), .A1(inst_cellmath__112[0]), .B0(N16122), .B1(N1922));
AO22XL inst_cellmath__113__115__U_2WWMM_I2812 (.Y(inst_cellmath__113[1]), .A0(N16178), .A1(inst_cellmath__112[1]), .B0(N16122), .B1(inst_cellmath__129[1]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2813 (.Y(inst_cellmath__113[2]), .A0(N16178), .A1(inst_cellmath__112[2]), .B0(N16122), .B1(inst_cellmath__129[2]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2814 (.Y(inst_cellmath__113[3]), .A0(N16178), .A1(inst_cellmath__112[3]), .B0(N16122), .B1(inst_cellmath__129[3]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2815 (.Y(inst_cellmath__113[4]), .A0(N16178), .A1(inst_cellmath__112[4]), .B0(N16122), .B1(inst_cellmath__129[4]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2816 (.Y(inst_cellmath__113[5]), .A0(N16178), .A1(inst_cellmath__112[5]), .B0(N16122), .B1(inst_cellmath__129[5]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2817 (.Y(inst_cellmath__113[6]), .A0(N16178), .A1(inst_cellmath__112[6]), .B0(N16122), .B1(inst_cellmath__129[6]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2818 (.Y(inst_cellmath__113[7]), .A0(N16178), .A1(inst_cellmath__112[7]), .B0(N16122), .B1(inst_cellmath__129[7]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2819 (.Y(inst_cellmath__113[8]), .A0(N16178), .A1(inst_cellmath__112[8]), .B0(N16122), .B1(inst_cellmath__129[8]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2820 (.Y(inst_cellmath__113[9]), .A0(N16178), .A1(inst_cellmath__112[9]), .B0(N16122), .B1(inst_cellmath__129[9]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2821 (.Y(inst_cellmath__113[10]), .A0(N16178), .A1(inst_cellmath__112[10]), .B0(N16122), .B1(inst_cellmath__129[10]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2822 (.Y(inst_cellmath__113[11]), .A0(N16178), .A1(inst_cellmath__112[11]), .B0(N16122), .B1(inst_cellmath__129[11]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2823 (.Y(inst_cellmath__113[12]), .A0(N16178), .A1(inst_cellmath__112[12]), .B0(N16122), .B1(inst_cellmath__129[12]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2824 (.Y(inst_cellmath__113[13]), .A0(N16178), .A1(inst_cellmath__112[13]), .B0(N16122), .B1(inst_cellmath__129[13]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2825 (.Y(inst_cellmath__113[14]), .A0(N16178), .A1(inst_cellmath__112[14]), .B0(N16122), .B1(inst_cellmath__129[14]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2826 (.Y(inst_cellmath__113[15]), .A0(N16178), .A1(inst_cellmath__112[15]), .B0(N16122), .B1(inst_cellmath__129[15]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2827 (.Y(inst_cellmath__113[16]), .A0(N16178), .A1(inst_cellmath__112[16]), .B0(N16122), .B1(inst_cellmath__129[16]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2828 (.Y(inst_cellmath__113[17]), .A0(N16178), .A1(inst_cellmath__112[17]), .B0(N16122), .B1(inst_cellmath__129[17]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2829 (.Y(inst_cellmath__113[18]), .A0(N16178), .A1(inst_cellmath__112[18]), .B0(N16122), .B1(inst_cellmath__129[18]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2830 (.Y(inst_cellmath__113[19]), .A0(N16178), .A1(inst_cellmath__112[19]), .B0(N16122), .B1(inst_cellmath__129[19]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2831 (.Y(inst_cellmath__113[20]), .A0(N16178), .A1(inst_cellmath__112[20]), .B0(N16122), .B1(inst_cellmath__129[20]));
AO22XL inst_cellmath__113__115__U_2WWMM_I2832 (.Y(inst_cellmath__113[21]), .A0(N16178), .A1(inst_cellmath__112[21]), .B0(N16122), .B1(inst_cellmath__129[21]));
AO21XL inst_cellmath__113__115__U_2WWMM_I2833 (.Y(inst_cellmath__113[22]), .A0(N16122), .A1(inst_cellmath__129[22]), .B0(N16178));
assign inst_cellmath__9[21] = inst_it2_lookup1_cellmath__53[0];
assign inst_cellmath__9[22] = inst_it2_lookup1_cellmath__53[1];
assign inst_cellmath__14[0] = 1'B0;
assign inst_cellmath__16[0] = 1'B0;
assign inst_cellmath__17[0] = 1'B0;
assign inst_cellmath__22[3] = inst_cellmath__22[4];
assign inst_lookup0_cellmath__27[0] = inst_it2_lookup1_cellmath__53[0];
assign inst_lookup0_cellmath__27[1] = inst_it2_lookup1_cellmath__53[1];
assign inst_lookup0_cellmath__29[0] = inst_cellmath__42[0];
assign inst_cellmath__30[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__30[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__30[2] = inst_cellmath__38__W1[2];
assign inst_cellmath__30[25] = inst_it2_cellmath__60[4];
assign inst_cellmath__31[0] = inst_cellmath__31[1];
assign inst_cellmath__34[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__34[1] = 1'B0;
assign inst_cellmath__34[2] = 1'B0;
assign inst_cellmath__35[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__35[1] = 1'B0;
assign inst_cellmath__35[2] = 1'B0;
assign inst_cellmath__38__W0[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__38__W0[1] = 1'B0;
assign inst_cellmath__38__W0[25] = 1'B0;
assign inst_cellmath__38__W1[0] = inst_it2_cellmath__60[4];
assign inst_cellmath__38__W1[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__39__W0[0] = inst_it2_cellmath__60[3];
assign inst_cellmath__39__W0[1] = inst_it2_cellmath__60[4];
assign inst_cellmath__39__W0[2] = inst_it2_cellmath__60[5];
assign inst_cellmath__39__W0[3] = inst_it2_cellmath__60[6];
assign inst_cellmath__39__W0[4] = inst_it2_cellmath__60[7];
assign inst_cellmath__39__W0[5] = inst_it2_cellmath__60[8];
assign inst_cellmath__39__W0[6] = inst_it2_cellmath__60[9];
assign inst_cellmath__39__W0[7] = inst_it2_cellmath__60[10];
assign inst_cellmath__39__W0[8] = inst_it2_cellmath__60[11];
assign inst_cellmath__39__W0[9] = inst_it2_cellmath__60[12];
assign inst_cellmath__39__W0[10] = inst_it2_cellmath__60[13];
assign inst_cellmath__39__W0[11] = inst_it2_cellmath__60[14];
assign inst_cellmath__39__W0[12] = inst_it2_cellmath__60[15];
assign inst_cellmath__39__W0[13] = inst_it2_cellmath__60[16];
assign inst_cellmath__39__W0[14] = inst_it2_cellmath__60[17];
assign inst_cellmath__39__W0[15] = inst_it2_cellmath__60[18];
assign inst_cellmath__39__W0[16] = inst_it2_cellmath__60[19];
assign inst_cellmath__39__W0[17] = inst_it2_cellmath__60[20];
assign inst_cellmath__39__W0[18] = inst_it2_cellmath__60[21];
assign inst_cellmath__39__W0[19] = inst_it2_cellmath__60[22];
assign inst_cellmath__39__W0[20] = inst_it2_cellmath__60[23];
assign inst_cellmath__39__W0[21] = inst_it2_cellmath__60[24];
assign inst_cellmath__39__W0[22] = inst_it2_cellmath__60[25];
assign inst_cellmath__39__W0[25] = 1'B0;
assign inst_cellmath__39__W1[0] = 1'B0;
assign inst_cellmath__39__W1[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__39__W1[2] = inst_it2_cellmath__61[4];
assign inst_cellmath__39__W1[3] = inst_it2_cellmath__61[5];
assign inst_cellmath__39__W1[4] = inst_it2_cellmath__61[6];
assign inst_cellmath__39__W1[5] = inst_it2_cellmath__61[7];
assign inst_cellmath__39__W1[6] = inst_it2_cellmath__61[8];
assign inst_cellmath__39__W1[7] = inst_it2_cellmath__61[9];
assign inst_cellmath__39__W1[8] = inst_it2_cellmath__61[10];
assign inst_cellmath__39__W1[9] = inst_it2_cellmath__61[11];
assign inst_cellmath__39__W1[10] = inst_it2_cellmath__61[12];
assign inst_cellmath__39__W1[11] = inst_it2_cellmath__61[13];
assign inst_cellmath__39__W1[12] = inst_it2_cellmath__61[14];
assign inst_cellmath__39__W1[13] = inst_it2_cellmath__61[15];
assign inst_cellmath__39__W1[14] = inst_it2_cellmath__61[16];
assign inst_cellmath__39__W1[15] = inst_it2_cellmath__61[17];
assign inst_cellmath__39__W1[16] = inst_it2_cellmath__61[18];
assign inst_cellmath__39__W1[17] = inst_it2_cellmath__61[19];
assign inst_cellmath__39__W1[18] = inst_it2_cellmath__61[20];
assign inst_cellmath__39__W1[19] = inst_it2_cellmath__61[21];
assign inst_cellmath__39__W1[20] = inst_it2_cellmath__61[22];
assign inst_cellmath__39__W1[21] = inst_it2_cellmath__61[23];
assign inst_cellmath__39__W1[22] = inst_it2_cellmath__61[24];
assign inst_cellmath__39__W1[23] = inst_it2_cellmath__61[25];
assign inst_cellmath__42[27] = 1'B0;
assign inst_cellmath__42[28] = 1'B0;
assign inst_cellmath__43[27] = 1'B0;
assign inst_cellmath__43[28] = 1'B0;
assign inst_cellmath__46[25] = 1'B0;
assign inst_cellmath__46[26] = 1'B0;
assign inst_cellmath__46[27] = 1'B0;
assign inst_cellmath__46[28] = 1'B0;
assign inst_cellmath__47[25] = 1'B0;
assign inst_cellmath__47[26] = 1'B0;
assign inst_cellmath__47[27] = 1'B0;
assign inst_cellmath__47[28] = 1'B0;
assign inst_it2_lookup1_cellmath__55[0] = inst_cellmath__40[0];
assign inst_it2_cellmath__56[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__56[1] = inst_it2_cellmath__63__W1[1];
assign inst_it2_cellmath__56[25] = inst_cellmath__14[2];
assign inst_it2_cellmath__57[0] = inst_it2_cellmath__57[1];
assign inst_it2_cellmath__60[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__60[1] = 1'B0;
assign inst_it2_cellmath__60[2] = 1'B0;
assign inst_it2_cellmath__61[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__61[1] = 1'B0;
assign inst_it2_cellmath__61[2] = 1'B0;
assign inst_it2_cellmath__62__W0[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__62__W0[1] = 1'B0;
assign inst_it2_cellmath__62__W0[2] = 1'B0;
assign inst_it2_cellmath__62__W0[25] = 1'B0;
assign inst_it2_cellmath__62__W1[0] = inst_cellmath__14[2];
assign inst_it2_cellmath__62__W1[1] = inst_it2_cellmath__63__W1[1];
assign inst_it2_cellmath__62__W1[2] = 1'B0;
assign inst_it2_cellmath__63__W1[0] = 1'B0;
assign inst_cellmath__67[8] = 1'B0;
assign inst_cellmath__67[9] = 1'B0;
assign inst_cellmath__120[0] = 1'B0;
assign inst_cellmath__124[28] = 1'B0;
endmodule

`ifdef arith_fdrq_A_bdw410776230_bdw_COMPILED
`else
`define arith_fdrq_A_bdw410776230_bdw_COMPILED
module arith_fdrq_A_bdw410776230_bdw (
	r,
	d,
	clk,
	q
	); /* architecture "gate_level" */ 
input  r,
	d;
input  clk;
output  q;
wire  data;
DFFQXL arith_fdrq_A_I0 (.Q(q), .D(data), .CK(clk));
AND2XL arith_fdrq_A_I1 (.Y(data), .A(d), .B(r));
endmodule
`endif //  `ifdef arith_fdrq_A_bdw410776230_bdw_COMPILED

/* CADENCE  urj4SgjfqBg= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



