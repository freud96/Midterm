/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:20:27 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__68,
	inst_cellmath__82;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [20:0] inst_cellmath__197;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire  inst_cellmath__219;
wire N487,N541,N542,N543,N544,N577,N580 
	,N608,N609,N610,N611,N612,N613,N614,N615 
	,N616,N617,N618,N619,N620,N621,N622,N623 
	,N624,N625,N626,N627,N628,N629,N630,N631 
	,N632,N633,N634,N635,N636,N637,N639,N640 
	,N641,N642,N643,N644,N645,N646,N647,N648 
	,N649,N650,N651,N652,N653,N654,N655,N656 
	,N657,N658,N659,N660,N661,N662,N663,N664 
	,N665,N666,N667,N668,N670,N675,N679,N680 
	,N681,N682,N683,N684,N685,N686,N687,N688 
	,N689,N690,N691,N692,N693,N694,N695,N696 
	,N697,N698,N699,N700,N701,N733,N734,N736 
	,N738,N739,N740,N741,N743,N744,N745,N746 
	,N747,N748,N749,N750,N751,N752,N753,N754 
	,N755,N757,N759,N770,N771,N776,N780,N3584 
	,N3657,N3658,N3659,N3660,N3661,N3662,N3665,N3666 
	,N5394,N5396,N5397,N5398,N5399,N5403,N5404,N5406 
	,N5407,N5408,N5409,N5410,N5411,N5413,N5414,N5416 
	,N5417,N5420,N5421,N5422,N5424,N5425,N5426,N5427 
	,N5430,N5431,N5433,N5434,N5435,N5436,N5437,N5438 
	,N5439,N5440,N5441,N5442,N5444,N5445,N5447,N5448 
	,N5450,N5451,N5452,N5453,N5454,N5455,N5457,N5459 
	,N5460,N5461,N5463,N5464,N5467,N5468,N5469,N5471 
	,N5472,N5473,N5475,N5476,N5477,N5478,N5479,N5480 
	,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488 
	,N5490,N5491,N5492,N5493,N5494,N5496,N5497,N5499 
	,N5501,N5503,N5504,N5505,N5507,N5508,N5510,N5512 
	,N5513,N5514,N5516,N5517,N5520,N5521,N5522,N5523 
	,N5524,N5525,N5526,N5528,N5529,N5530,N5532,N5533 
	,N5534,N5535,N5536,N5538,N5539,N5540,N5541,N5542 
	,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5551 
	,N5552,N5554,N5555,N5556,N5557,N5558,N5560,N5562 
	,N5564,N5568,N5569,N5570,N5571,N5573,N5574,N5576 
	,N5577,N5578,N5579,N5580,N5582,N5583,N5584,N5585 
	,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593 
	,N5594,N5595,N5598,N5600,N5603,N5604,N5605,N5606 
	,N5607,N5609,N5610,N5611,N5612,N5613,N5614,N5618 
	,N5619,N5620,N5621,N5622,N5623,N5624,N5626,N5627 
	,N5628,N5631,N5632,N5633,N5635,N5636,N5639,N5640 
	,N5641,N5642,N5643,N5645,N5646,N5648,N5650,N5651 
	,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659 
	,N5660,N5661,N5663,N5664,N5665,N5667,N5668,N5669 
	,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677 
	,N5678,N5680,N5681,N5682,N5683,N5684,N5685,N5686 
	,N5687,N5688,N5692,N5693,N5694,N5695,N5698,N5699 
	,N5700,N5701,N5702,N5703,N5704,N5705,N5707,N5708 
	,N5710,N5711,N5714,N5715,N5717,N5718,N5719,N5720 
	,N5721,N5724,N5725,N5726,N5727,N5729,N5730,N5731 
	,N5732,N5734,N5735,N5736,N5737,N5738,N5739,N5740 
	,N5742,N5744,N5745,N5746,N5747,N5748,N5749,N5751 
	,N5753,N5754,N5756,N5757,N5758,N5759,N5760,N5761 
	,N5764,N5766,N5768,N5769,N5770,N5773,N5774,N5775 
	,N5776,N5777,N5778,N5779,N5780,N5781,N5783,N5784 
	,N5785,N5786,N5787,N5788,N5789,N5791,N5792,N5794 
	,N5795,N5796,N5797,N5798,N5800,N5802,N5805,N5806 
	,N5807,N5808,N5810,N5811,N5812,N5813,N5814,N5815 
	,N5816,N5817,N5818,N5819,N5820,N5821,N5823,N5825 
	,N5826,N5827,N5828,N5829,N5830,N5831,N5833,N5835 
	,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845 
	,N5847,N5848,N5849,N5850,N5851,N5852,N5854,N5856 
	,N5857,N5858,N5859,N5860,N5862,N5863,N5866,N5869 
	,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5878 
	,N5880,N5884,N5885,N5886,N5887,N5888,N5889,N5890 
	,N5891,N5892,N5893,N5895,N5898,N5899,N5900,N5903 
	,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911 
	,N5912,N5913,N5914,N5916,N5917,N5918,N5919,N5920 
	,N5921,N5922,N5924,N5925,N5926,N5927,N5928,N5929 
	,N5931,N5932,N5934,N5935,N5936,N5938,N5939,N5940 
	,N5941,N5942,N5943,N5944,N5945,N5946,N5948,N5950 
	,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958 
	,N5960,N5961,N5962,N5965,N5966,N5967,N5968,N5969 
	,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977 
	,N5978,N5979,N5980,N5983,N5984,N5985,N5986,N5987 
	,N5989,N5990,N5991,N5992,N5993,N5994,N5996,N6000 
	,N6001,N6002,N6004,N6006,N6007,N6008,N6009,N6010 
	,N6011,N6012,N6013,N6014,N6019,N6020,N6021,N6022 
	,N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6033 
	,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6042 
	,N6043,N6044,N6045,N6046,N6047,N6049,N6050,N6051 
	,N6052,N6053,N6054,N6056,N6057,N6058,N6059,N6060 
	,N6061,N6063,N6064,N6066,N6067,N6068,N6069,N6070 
	,N6073,N6075,N6076,N6077,N6078,N6079,N6081,N6082 
	,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090 
	,N6091,N6092,N6093,N6096,N6097,N6098,N6099,N6100 
	,N6101,N6102,N6103,N6105,N6107,N6108,N6110,N6111 
	,N6112,N6113,N6115,N6116,N6117,N6119,N6120,N6121 
	,N6123,N6124,N6125,N6126,N6128,N6130,N6131,N6132 
	,N6133,N6136,N6139,N6140,N6141,N6142,N6143,N6144 
	,N6145,N6146,N6147,N6148,N6150,N6151,N6152,N6153 
	,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162 
	,N6163,N6164,N6165,N6168,N6169,N6171,N6172,N6173 
	,N6174,N6175,N6176,N6177,N6178,N6181,N6182,N6183 
	,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191 
	,N6192,N6193,N6195,N6198,N6199,N6200,N6203,N6205 
	,N6206,N6207,N6208,N6209,N6210,N6211,N6212,N6213 
	,N6214,N6216,N6218,N6219,N6220,N6221,N6222,N6223 
	,N6225,N6226,N6227,N6228,N6230,N6231,N6232,N6234 
	,N6235,N6236,N6237,N6238,N6239,N6240,N6241,N6242 
	,N6243,N6244,N6245,N6248,N6249,N6250,N6251,N6252 
	,N6253,N7100,N7102,N7103,N7107,N7108,N7121,N7123 
	,N7124,N7125,N7127,N7128,N7131,N7132,N7134,N7135 
	,N7136,N7138,N7140,N7144,N7146,N7147,N7149,N7151 
	,N7152,N7154,N7156,N7157,N7160,N7162,N7163,N7165 
	,N7166,N7168,N7169,N7171,N7173,N7175,N7176,N7178 
	,N7179,N7181,N7182,N7184,N7187,N7189,N7190,N7192 
	,N7194,N7195,N7196,N7197,N7200,N7202,N7203,N7204 
	,N7206,N7209,N7210,N7212,N7213,N7215,N7217,N7219 
	,N7220,N7222,N7224,N7225,N7227,N7229,N7230,N7233 
	,N7234,N7236,N7238,N7239,N7243,N7245,N7246,N7248 
	,N7249,N7252,N7255,N7256,N7258,N7259,N7261,N7263 
	,N7265,N7266,N7267,N7269,N7270,N7271,N7273,N7275 
	,N7276,N7278,N7280,N7281,N7283,N7287,N7289,N7290 
	,N7292,N7293,N7295,N7297,N7298,N7299,N7301,N7304 
	,N7306,N7307,N7309,N7310,N7311,N7313,N7315,N7316 
	,N7319,N7321,N7322,N7324,N7325,N7327,N7330,N7331 
	,N7333,N7334,N7335,N7336,N7337,N7339,N7341,N7344 
	,N7346,N7347,N7349,N7350,N7352,N7354,N7355,N7357 
	,N7359,N7361,N7364,N7365,N7367,N7368,N7370,N7371 
	,N7373,N7631,N7669,N7670,N7672,N7673,N7675,N7676 
	,N7677,N7678,N7679,N7680,N7682,N7683,N7684,N7685 
	,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694 
	,N7695,N7696,N7697,N7698,N7699,N7700,N7701,N7703 
	,N7704,N7705,N7706,N7708,N7709,N7710,N7711,N7712 
	,N7715,N7716,N7717,N7718,N7719,N7720,N7721,N7723 
	,N7725,N7726,N7727,N7728,N7729,N7730,N7732,N7733 
	,N7734,N7735,N7736,N7737,N7738,N7739,N7740,N7741 
	,N7742,N7743,N7744,N7746,N7747,N7748,N7749,N7750 
	,N7752,N7753,N7754,N7755,N7757,N7759,N7760,N7761 
	,N7762,N7763,N7764,N7765,N7766,N7767,N7769,N7770 
	,N7771,N7772,N7773,N7775,N7776,N7777,N7778,N7779 
	,N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787 
	,N7788,N7789,N7790,N7791,N7792,N7793,N7794,N7797 
	,N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805 
	,N7806,N7807,N7809,N7810,N7811,N7812,N7813,N7814 
	,N7815,N7816,N7817,N7819,N7820,N7821,N7822,N7823 
	,N7824,N7826,N7827,N7829,N7830,N7831,N7832,N7833 
	,N7834,N7835,N7838,N7839,N7841,N7843,N7844,N7845 
	,N7846,N7848,N7849,N7851,N7852,N7854,N7855,N7856 
	,N7857,N7858,N7859,N7860,N7861,N7862,N7863,N7864 
	,N7865,N7867,N7868,N7870,N7871,N7872,N7873,N7874 
	,N7875,N7876,N7877,N7878,N7881,N7882,N7883,N7884 
	,N7885,N7886,N7887,N7888,N7890,N7891,N7892,N7894 
	,N7896,N7897,N7898,N7899,N7900,N7901,N7902,N7903 
	,N7904,N7906,N7908,N7910,N7911,N7913,N7915,N7916 
	,N7917,N7918,N7919,N7920,N7921,N7923,N7924,N7925 
	,N7926,N7928,N7929,N7930,N7931,N7932,N7933,N7934 
	,N7935,N7936,N7937,N7938,N7939,N7940,N7941,N7942 
	,N7943,N7945,N7946,N7947,N7949,N7950,N7951,N7952 
	,N7953,N7954,N7955,N7956,N7957,N7958,N7959,N7960 
	,N7961,N7962,N7964,N7965,N7966,N7967,N7968,N7969 
	,N7970,N7971,N7972,N7974,N7975,N7976,N7977,N7978 
	,N7979,N7982,N7983,N7985,N7986,N7987,N7988,N7989 
	,N7990,N7991,N7992,N7993,N7994,N7995,N7997,N7998 
	,N7999,N8000,N8001,N8002,N8003,N8004,N8006,N8008 
	,N8009,N8010,N8011,N8012,N8016,N8017,N8018,N8019 
	,N8020,N8021,N8022,N8023,N8025,N8026,N8027,N8028 
	,N8029,N8032,N8033,N8034,N8035,N8036,N8037,N8038 
	,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046 
	,N8047,N8048,N8050,N8052,N8053,N8054,N8055,N8056 
	,N8057,N8058,N8059,N8060,N8061,N8062,N8063,N8064 
	,N8065,N8067,N8068,N8069,N8070,N8071,N8072,N8075 
	,N8076,N8078,N8079,N8080,N8081,N8082,N8083,N8084 
	,N8086,N8087,N8088,N8089,N8090,N8091,N8092,N8093 
	,N8094,N8095,N8097,N8098,N8099,N8101,N8102,N8103 
	,N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111 
	,N8112,N8113,N8115,N8116,N8118,N8119,N8120,N8123 
	,N8124,N8125,N8126,N8127,N8128,N8129,N8130,N8131 
	,N8132,N8133,N8134,N8135,N8136,N8138,N8139,N8140 
	,N8141,N8143,N8144,N8145,N8146,N8147,N8148,N8150 
	,N8151,N8152,N8153,N8154,N8157,N8158,N8160,N8161 
	,N8162,N8163,N8164,N8165,N8166,N8167,N8169,N8170 
	,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178 
	,N8180,N8182,N8183,N8185,N8187,N8188,N8189,N8190 
	,N8191,N8192,N8195,N8196,N8197,N8198,N8200,N8201 
	,N8202,N8204,N8205,N8206,N8207,N8208,N8209,N8210 
	,N8211,N8212,N8213,N8215,N8216,N8217,N8218,N8219 
	,N8223,N8224,N8225,N8226,N8227,N8228,N8229,N8230 
	,N8231,N8232,N8233,N8234,N8235,N8236,N8237,N8238 
	,N8239,N8242,N8243,N8244,N8245,N8246,N8247,N8249 
	,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257 
	,N8258,N8260,N8262,N8263,N8264,N8265,N8267,N8269 
	,N8272,N8273,N8274,N8275,N8276,N8277,N8278,N8280 
	,N8282,N8283,N8284,N8285,N8286,N8287,N8288,N8290 
	,N8291,N8292,N8293,N8294,N8295,N8297,N8298,N8299 
	,N8300,N8301,N8302,N8303,N8304,N8305,N8307,N8308 
	,N8309,N8310,N8312,N8313,N8314,N8315,N8316,N8317 
	,N8319,N8321,N8322,N8323,N8324,N8325,N8326,N8327 
	,N8328,N8329,N8330,N8331,N8334,N8335,N8336,N8338 
	,N8339,N8340,N8341,N8342,N8344,N8345,N8348,N8349 
	,N8350,N8351,N8352,N8354,N8355,N8356,N8358,N8360 
	,N8361,N8362,N8363,N8364,N8365,N8366,N8367,N8370 
	,N8371,N8372,N8373,N8374,N8375,N8376,N8378,N8379 
	,N8380,N8381,N8383,N8384,N8385,N8386,N8388,N8389 
	,N8390,N8391,N8392,N8393,N8394,N8395,N8396,N8397 
	,N8399,N8400,N8401,N8402,N8403,N8405,N8408,N8410 
	,N8413,N8414,N8415,N8416,N8417,N8418,N8419,N8420 
	,N8421,N8422,N8424,N8425,N8426,N8427,N8428,N8429 
	,N8430,N8431,N8432,N8433,N8434,N8435,N8436,N8437 
	,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445 
	,N8446,N8447,N8449,N8450,N8452,N8453,N8454,N8455 
	,N8456,N8457,N8458,N8459,N8460,N8461,N8462,N8463 
	,N8464,N8466,N8467,N8468,N8469,N8470,N8472,N8473 
	,N8474,N8475,N8477,N8478,N8479,N8480,N8481,N8483 
	,N8484,N8485,N8486,N8488,N8489,N8490,N8492,N8493 
	,N8494,N8495,N8497,N8498,N8500,N8501,N8502,N8503 
	,N8504,N8506,N8507,N8509,N8510,N8511,N8512,N8514 
	,N8517,N8518,N8519,N8520,N8521,N8522,N8523,N8524 
	,N8525,N8526,N8527,N8528,N8529,N8531,N8532,N8533 
	,N8534,N8535,N8536,N8537,N8538,N8539,N8540,N8541 
	,N8542,N8543,N8545,N8546,N8547,N8549,N8550,N8552 
	,N8553,N8554,N8555,N8556,N8557,N8558,N8559,N8560 
	,N8561,N8562,N8563,N8564,N8565,N8566,N8567,N8568 
	,N8569,N8571,N8573,N8574,N8575,N8576,N8577,N8578 
	,N8579,N8580,N8581,N8582,N8584,N8585,N8586,N8587 
	,N8589,N8590,N8591,N8593,N8594,N8596,N8597,N8598 
	,N8599,N8601,N8602,N8605,N8606,N8607,N8608,N8609 
	,N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617 
	,N8618,N8620,N8621,N8622,N8624,N8625,N8626,N8627 
	,N8629,N8630,N8632,N8633,N8634,N8636,N8637,N8638 
	,N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8647 
	,N8648,N8649,N8650,N8651,N8652,N8653,N8655,N8656 
	,N8657,N8658,N8659,N8660,N8661,N8662,N8663,N8664 
	,N8665,N8666,N8667,N8669,N8671,N8673,N8674,N8675 
	,N8676,N8677,N8678,N8679,N8681,N8683,N8684,N8685 
	,N8686,N8687,N8688,N8690,N8692,N8694,N8696,N8697 
	,N8698,N8700,N8701,N8702,N8703,N8705,N8706,N8707 
	,N8708,N8709,N8710,N8711,N8712,N8713,N8714,N8715 
	,N8716,N8717,N8719,N8720,N8721,N8722,N8723,N8724 
	,N8725,N8727,N8728,N8729,N8730,N8731,N8732,N8734 
	,N8735,N8736,N8737,N8738,N8739,N8740,N8741,N8742 
	,N8743,N8745,N8746,N8747,N8749,N8752,N8753,N8754 
	,N8755,N8756,N8757,N8759,N8762,N8763,N8764,N8765 
	,N8767,N8768,N8769,N8770,N8771,N8772,N8773,N8774 
	,N8775,N8776,N8777,N8778,N8779,N8781,N8782,N8783 
	,N8784,N8785,N8787,N8788,N9903,N9906,N9907,N9908 
	,N9909,N9911,N9912,N9914,N9915,N9916,N9917,N9918 
	,N9919,N9920,N9922,N9923,N9925,N9927,N9928,N9929 
	,N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937 
	,N9938,N9939,N9940,N9941,N9942,N9943,N9944,N9945 
	,N9946,N9947,N9948,N9951,N9952,N9953,N9954,N9955 
	,N9957,N9958,N9959,N9960,N9961,N9962,N9963,N9964 
	,N9965,N9966,N9967,N9968,N9969,N9970,N9971,N9972 
	,N9973,N9975,N9976,N9977,N9978,N9979,N9980,N9981 
	,N9982,N9983,N9985,N9986,N9987,N9988,N9989,N9990 
	,N9991,N9992,N9993,N9994,N9995,N9996,N9997,N9999 
	,N10000,N10002,N10004,N10006,N10008,N10009,N10010,N10011 
	,N10012,N10013,N10014,N10015,N10016,N10017,N10018,N10020 
	,N10021,N10022,N10023,N10024,N10025,N10029,N10031,N10032 
	,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041 
	,N10042,N10043,N10044,N10046,N10047,N10049,N10050,N10051 
	,N10052,N10054,N10055,N10056,N10058,N10059,N10062,N10063 
	,N10065,N10066,N10068,N10069,N10070,N10071,N10073,N10075 
	,N10076,N10077,N10078,N10079,N10080,N10081,N10082,N10083 
	,N10084,N10085,N10086,N10087,N10089,N10090,N10091,N10092 
	,N10093,N10094,N10096,N10097,N10098,N10099,N10100,N10101 
	,N10102,N10103,N10104,N10105,N10106,N10108,N10109,N10110 
	,N10111,N10112,N10113,N10115,N10117,N10118,N10119,N10120 
	,N10121,N10122,N10123,N10124,N10125,N10126,N10127,N10128 
	,N10129,N10130,N10131,N10132,N10133,N10134,N10136,N10137 
	,N10138,N10140,N10142,N10143,N10144,N10145,N10146,N10147 
	,N10148,N10149,N10150,N10151,N10152,N10154,N10155,N10156 
	,N10157,N10158,N10159,N10161,N10162,N10164,N10166,N10167 
	,N10168,N10169,N10170,N10171,N10172,N10173,N10174,N10175 
	,N10176,N10177,N10178,N10179,N10180,N10181,N10182,N10183 
	,N10185,N10187,N10188,N10189,N10190,N10191,N10192,N10194 
	,N10195,N10196,N10197,N10198,N10199,N10200,N10201,N10202 
	,N10203,N10204,N10205,N10206,N10207,N10208,N10209,N10210 
	,N10211,N10212,N10213,N10214,N10215,N10216,N10218,N10219 
	,N10221,N10222,N10223,N10224,N10226,N10227,N10228,N10229 
	,N10230,N10231,N10232,N10233,N10234,N10235,N10237,N10238 
	,N10239,N10241,N10242,N10243,N10244,N10245,N10246,N10247 
	,N10249,N10252,N10254,N10255,N10256,N10257,N10258,N10260 
	,N10261,N10263,N10264,N10265,N10266,N10267,N10269,N10271 
	,N10273,N10275,N10276,N10277,N10278,N10279,N10280,N10281 
	,N10284,N10285,N10286,N10287,N10288,N10289,N10290,N10291 
	,N10292,N10293,N10294,N10295,N10296,N10298,N10299,N10301 
	,N10302,N10303,N10304,N10305,N10306,N10307,N10308,N10310 
	,N10311,N10312,N10313,N10314,N10315,N10316,N10317,N10318 
	,N10319,N10321,N10322,N10324,N10325,N10326,N10327,N10328 
	,N10329,N10331,N10333,N10334,N10335,N10336,N10337,N10338 
	,N10339,N10341,N10342,N10343,N10344,N10345,N10346,N10347 
	,N10348,N10349,N10351,N10352,N10353,N10354,N10355,N10356 
	,N10357,N10358,N10359,N10361,N10362,N10363,N10364,N10365 
	,N10367,N10368,N10369,N10370,N10371,N10372,N10373,N10374 
	,N10376,N10377,N10378,N10379,N10380,N10381,N10382,N10383 
	,N10384,N10385,N10386,N10387,N10388,N10389,N10390,N10393 
	,N10394,N10395,N10396,N10397,N10399,N10400,N10401,N10402 
	,N10403,N10404,N10405,N10408,N10409,N10410,N10412,N10413 
	,N10414,N10416,N10417,N10418,N10419,N10420,N10421,N10422 
	,N10423,N10424,N10425,N10426,N10427,N10431,N10432,N10433 
	,N10434,N10436,N10437,N10438,N10439,N10440,N10442,N10443 
	,N10445,N10446,N10447,N10448,N10449,N10450,N10451,N10452 
	,N10456,N10457,N10458,N10459,N10460,N10463,N10464,N10465 
	,N10466,N10467,N10468,N10469,N10470,N10471,N10472,N10473 
	,N10475,N10476,N10477,N10478,N10479,N10480,N10481,N10482 
	,N10483,N10484,N10486,N10487,N10488,N10489,N10490,N10491 
	,N10492,N10493,N10494,N10495,N10496,N10497,N10498,N10500 
	,N10502,N10503,N10505,N10506,N10507,N10508,N10509,N10510 
	,N10511,N10512,N10515,N10516,N10518,N10519,N10520,N10521 
	,N10523,N10524,N10525,N10526,N10527,N10528,N10529,N10532 
	,N10533,N10534,N10535,N10536,N10538,N10539,N11160,N11161 
	,N11162,N11163,N11164,N11165,N11166,N11168,N11169,N11170 
	,N11171,N11172,N11173,N11174,N11175,N11176,N11177,N11178 
	,N11179,N11180,N11181,N11182,N11183,N11184,N11185,N11186 
	,N11187,N11188,N11189,N11191,N11192,N11193,N11194,N11195 
	,N11196,N11197,N11199,N11201,N11203,N11205,N11206,N11207 
	,N11208,N11209,N11210,N11211,N11212,N11214,N11215,N11216 
	,N11217,N11218,N11220,N11222,N11223,N11224,N11225,N11226 
	,N11227,N11228,N11230,N11231,N11233,N11234,N11235,N11236 
	,N11237,N11238,N11239,N11240,N11241,N11242,N11244,N11245 
	,N11246,N11247,N11248,N11249,N11251,N11253,N11254,N11255 
	,N11256,N11257,N11258,N11259,N11260,N11261,N11262,N11263 
	,N11264,N11265,N11266,N11267,N11268,N11269,N11270,N11272 
	,N11273,N11274,N11275,N11276,N11277,N11278,N11280,N11281 
	,N11282,N11283,N11284,N11285,N11287,N11288,N11289,N11290 
	,N11291,N11292,N11293,N11294,N11295,N11298,N11299,N11301 
	,N11302,N11303,N11304,N11305,N11306,N11307,N11308,N11309 
	,N11310,N11311,N11312,N11313,N11314,N11316,N11317,N11318 
	,N11319,N11320,N11321,N11322,N11323,N11325,N11326,N11327 
	,N11328,N11329,N11330,N11331,N11332,N11333,N11335,N11336 
	,N11337,N11338,N11339,N11340,N11341,N11342,N11343,N11344 
	,N11345,N11346,N11347,N11349,N11350,N11351,N11352,N11353 
	,N11354,N11355,N11356,N11357,N11360,N11361,N11362,N11363 
	,N11364,N11365,N11367,N11368,N11369,N11370,N11371,N11372 
	,N11373,N11375,N11376,N11377,N11378,N11379,N11380,N11382 
	,N11383,N11385,N11386,N11387,N11388,N11389,N11390,N11391 
	,N11392,N11393,N11395,N11396,N11397,N11398,N11399,N11400 
	,N11401,N11402,N11404,N11405,N11407,N11408,N11409,N11410 
	,N11411,N11412,N11413,N11415,N11416,N11417,N11418,N11419 
	,N11420,N11421,N11423,N11424,N11425,N11427,N11428,N11429 
	,N11430,N11432,N11433,N11434,N11435,N11436,N11437,N11438 
	,N11439,N11440,N11441,N11442,N11443,N11445,N11447,N11448 
	,N11449,N11450,N11451,N11453,N11454,N11456,N11457,N11458 
	,N11459,N11460,N11461,N11462,N11463,N11464,N11465,N11466 
	,N11467,N11468,N11470,N11471,N11472,N11474,N11476,N11477 
	,N11479,N11480,N11481,N11483,N11484,N11485,N11486,N11487 
	,N11488,N11489,N11490,N11491,N11492,N11493,N11494,N11495 
	,N11497,N11498,N11499,N11500,N11501,N11502,N11503,N11504 
	,N11505,N11506,N11507,N11508,N11509,N11511,N11512,N11513 
	,N11514,N11516,N11519,N11520,N11521,N11522,N11523,N11524 
	,N11525,N11526,N11527,N11528,N11529,N11530,N11531,N11532 
	,N11533,N11534,N11535,N11536,N11538,N11539,N11540,N11541 
	,N11542,N11543,N11544,N11545,N11547,N11548,N11549,N11550 
	,N11551,N11552,N11553,N11554,N11555,N11556,N11557,N11558 
	,N11559,N11560,N11561,N11562,N11563,N11564,N11565,N11566 
	,N11567,N11568,N11569,N11570,N11571,N11572,N11574,N11575 
	,N11576,N11577,N11578,N11579,N11580,N11582,N11583,N11584 
	,N11585,N11588,N11589,N11590,N11591,N11592,N11593,N11594 
	,N11595,N11598,N11599,N11600,N11601,N11602,N11603,N11605 
	,N11606,N11607,N11610,N11611,N11612,N11613,N11614,N11615 
	,N11616,N11617,N11618,N11619,N11620,N11621,N11622,N11623 
	,N11624,N11625,N11626,N11627,N11628,N11630,N11631,N11632 
	,N11633,N11634,N11635,N11636,N11637,N11638,N11639,N11640 
	,N11641,N11642,N11643,N11644,N11645,N11646,N11647,N11648 
	,N11649,N11650,N11652,N11653,N11654,N11655,N11657,N11658 
	,N11659,N11660,N11662,N11663,N11664,N11665,N11666,N11667 
	,N11668,N11670,N11671,N11672,N11673,N11674,N11675,N11676 
	,N11677,N11678,N11679,N11680,N11681,N11682,N11683,N11684 
	,N11685,N11686,N11687,N11688,N11690,N11691,N11692,N11694 
	,N11695,N11696,N11697,N11698,N11700,N11701,N11702,N11703 
	,N11704,N11705,N11706,N11707,N11708,N11709,N11710,N11711 
	,N11712,N11713,N11715,N11716,N11718,N11719,N11720,N11721 
	,N11722,N11723,N11724,N11725,N11727,N11728,N11729,N11730 
	,N11731,N11732,N11733,N11734,N11737,N11739,N11740,N11741 
	,N11742,N11743,N11744,N11745,N11746,N11747,N11748,N11749 
	,N11750,N11752,N11753,N11754,N11755,N11756,N11757,N11758 
	,N11760,N11761,N11762,N11763,N11764,N11765,N11767,N11768 
	,N11770,N11771,N11772,N11773,N11774,N11775,N11776,N11777 
	,N11778,N11780,N11781,N11782,N11783,N11784,N11785,N11786 
	,N11788,N11790,N11791,N11792,N11793,N11794,N11795,N11796 
	,N11799,N11800,N11801,N11802,N11803,N11804,N11805,N11806 
	,N11809,N11810,N11811,N11812,N11813,N11814,N11816,N11819 
	,N11820,N11821,N11823,N11824,N11825,N11826,N11827,N11828 
	,N11829,N11830,N11832,N11833,N11834,N11835,N11836,N11837 
	,N11839,N11840,N11842,N11843,N11844,N11845,N11846,N11847 
	,N11848,N11849,N11850,N11851,N11852,N11853,N11854,N11855 
	,N11856,N11858,N11859,N11861,N11862,N11863,N11864,N11867 
	,N11868,N11869,N11870,N11871,N11872,N11873,N11874,N11875 
	,N11876,N11877,N11878,N11879,N11880,N11881,N11882,N11884 
	,N11885,N11886,N11887,N11888,N11889,N11890,N11891,N11892 
	,N11894,N11895,N11896,N11897,N11899,N11900,N11901,N11902 
	,N11904,N11905,N11906,N11909,N11910,N11911,N11912,N11913 
	,N11914,N11915,N11916,N11917,N11918,N11919,N11920,N11921 
	,N11922,N11923,N11924,N11925,N11926,N11927,N11929,N11930 
	,N11931,N11932,N11933,N11934,N11936,N11937,N11938,N11939 
	,N11940,N11941,N11943,N11944,N11945,N11946,N11947,N11948 
	,N11949,N11950,N11951,N11952,N11953,N11954,N11955,N11956 
	,N11957,N11958,N11959,N11960,N11961,N11962,N11963,N11965 
	,N11966,N11967,N11968,N11969,N11970,N11971,N11972,N11973 
	,N11976,N11977,N11978,N11979,N11980,N11982,N11983,N11984 
	,N11985,N11986,N11987,N11988,N11989,N11990,N11991,N11992 
	,N11993,N11994,N11995,N11998,N11999,N12000,N12001,N12003 
	,N12004,N12007,N12008,N12009,N12010,N12011,N12012,N12013 
	,N12014,N12015,N12016,N12017,N12018,N12019,N12020,N12021 
	,N12022,N12023,N12024,N12025,N12026,N12028,N12029,N12030 
	,N12032,N12033,N12034,N12035,N12036,N12037,N12038,N12039 
	,N12040,N12042,N12043,N12044,N12045,N12046,N12047,N12050 
	,N12051,N12052,N12053,N12054,N12055,N12056,N12058,N12059 
	,N12060,N12061,N12062,N12064,N12065,N12066,N12067,N12068 
	,N12070,N12071,N12072,N12073,N12074,N12075,N12076,N12077 
	,N12078,N12079,N12080,N12081,N12082,N12083,N12084,N12085 
	,N12086,N12087,N12088,N12089,N12090,N12091,N12093,N12094 
	,N12095,N12096,N12097,N12099,N12100,N12101,N12102,N12103 
	,N12104,N12105,N12106,N12107,N12108,N12109,N12110,N12111 
	,N12113,N12114,N12115,N12116,N12117,N12118,N12119,N12120 
	,N12121,N12122,N12123,N12124,N12125,N12128,N12129,N12130 
	,N12133,N12134,N12135,N12136,N12137,N12138,N12139,N12140 
	,N12141,N12142,N12143,N12144,N12145,N12146,N12148,N12149 
	,N12150,N12151,N12153,N12154,N12155,N12156,N12158,N12159 
	,N12161,N12162,N12163,N12164,N12165,N12166,N12167,N12168 
	,N12169,N12170,N12171,N12172,N12173,N12174,N12175,N12176 
	,N12177,N12178,N12179,N12181,N12182,N12183,N12184,N12185 
	,N12186,N12188,N12190,N12191,N12192,N12194,N12196,N12198 
	,N12199,N12200,N12201,N12202,N12204,N12205,N12206,N12207 
	,N12208,N12209,N12210,N12211,N12212,N12213,N12214,N12216 
	,N12218,N12219,N12220,N12221,N12223,N12224,N12226,N12227 
	,N12228,N12229,N12230,N12231,N12232,N12233,N12234,N12235 
	,N12236,N12237,N12238,N12239,N12240,N12242,N12243,N12244 
	,N12245,N12246,N12247,N12250,N12252,N12253,N12254,N12255 
	,N12256,N12257,N12258,N12259,N12260,N12261,N12262,N12263 
	,N12264,N12265,N12267,N12268,N12269,N12270,N12271,N12272 
	,N12273,N12274,N12275,N12276,N12277,N12279,N12280,N12281 
	,N12283,N12284,N12286,N12288,N12290,N12291,N12292,N12293 
	,N12294,N12295,N12296,N12297,N12298,N12299,N12300,N12301 
	,N12302,N12303,N12304,N12305,N12306,N12307,N12308,N12309 
	,N12310,N12311,N12313,N12314,N12315,N12316,N12318,N12319 
	,N12320,N12321,N12322,N12323,N12324,N12325,N12326,N12327 
	,N12328,N12329,N12330,N12331,N12332,N12333,N12334,N12335 
	,N12336,N12337,N12338,N12339,N12340,N12341,N12343,N12344 
	,N12345,N12346,N12348,N12350,N12351,N12352,N12353,N12354 
	,N12355,N12356,N12357,N12358,N12359,N12360,N12361,N12362 
	,N12363,N12364,N12365,N12366,N12367,N12368,N12370,N12371 
	,N12373,N12374,N12375,N12376,N12379,N12381,N12382,N12383 
	,N12384,N12385,N12386,N12387,N12388,N12389,N12390,N12391 
	,N12392,N12393,N12394,N12395,N12396,N12398,N12399,N12400 
	,N12401,N12402,N12403,N12405,N12406,N12407,N12408,N12410 
	,N12411,N12412,N12414,N12415,N12416,N12418,N12419,N12420 
	,N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428 
	,N12429,N12430,N12431,N12432,N12433,N12435,N12436,N12437 
	,N12438,N12440,N12441,N12442,N12443,N12444,N12445,N12446 
	,N12447,N12448,N12449,N12450,N12451,N12452,N12453,N12454 
	,N12455,N12456,N12458,N12459,N12460,N12461,N12462,N12464 
	,N12465,N12466,N12467,N12468,N12469,N12470,N12471,N12472 
	,N12473,N12474,N12475,N12477,N12478,N12479,N12480,N12481 
	,N12482,N12483,N12484,N12485,N12486,N12487,N12488,N12489 
	,N12490,N12491,N12492,N12493,N12494,N12496,N12497,N12498 
	,N12499,N12502,N12503,N12504,N12505,N12506,N12507,N12508 
	,N12509,N12510,N12511,N12512,N12513,N12514,N12515,N12516 
	,N12517,N12518,N12519,N12520,N12522,N12523,N12524,N12525 
	,N12526,N12527,N12529,N12530,N12531,N12532,N12533,N12534 
	,N12535,N12536,N12537,N12538,N12539,N12540,N12541,N12542 
	,N12543,N12544,N12545,N12546,N12547,N12548,N12549,N12550 
	,N12551,N12552,N12554,N12555,N12556,N12557,N12558,N12559 
	,N12561,N12562,N12563,N12565,N12566,N12567,N12568,N12569 
	,N12570,N12571,N12572,N12573,N12574,N12575,N12576,N12578 
	,N12579,N12580,N12581,N12582,N12584,N12586,N12587,N12588 
	,N12589,N12590,N12591,N12592,N12593,N12594,N12595,N12596 
	,N12597,N12599,N12600,N12601,N12602,N12603,N12604,N12606 
	,N12607,N12608,N12609,N12611,N12612,N12613,N12614,N12615 
	,N12616,N12617,N12618,N12619,N12620,N12621,N12622,N12623 
	,N12625,N12626,N12627,N12628,N12629,N12630,N12632,N12634 
	,N12635,N12636,N12637,N12638,N12639,N12641,N12642,N12643 
	,N12647,N12648,N12649,N12650,N12651,N12652,N12653,N12655 
	,N12656,N12657,N12658,N12659,N12660,N12661,N12662,N12663 
	,N12664,N12665,N12667,N12668,N12669,N12670,N12671,N12673 
	,N12674,N12675,N12676,N12677,N12678,N12679,N12680,N12681 
	,N12682,N12683,N12684,N12685,N12686,N12687,N12688,N12689 
	,N12690,N12691,N12692,N12693,N12695,N12696,N12697,N12700 
	,N12701,N12702,N12703,N12704,N12705,N12706,N12707,N12708 
	,N12709,N12710,N12711,N12712,N12713,N12714,N12715,N12716 
	,N12717,N12719,N12720,N12721,N12722,N12723,N12725,N12728 
	,N12729,N12730,N12731,N12732,N12733,N12734,N12735,N12736 
	,N12737,N12739,N12740,N12741,N12742,N12743,N12744,N12745 
	,N12746,N12747,N12748,N12749,N12750,N12751,N12752,N12753 
	,N12754,N12756,N12757,N12758,N12759,N12760,N12761,N12763 
	,N12764,N12765,N12767,N12768,N12769,N12770,N12771,N12772 
	,N12773,N12775,N12776,N12777,N12778,N12779,N12780,N12782 
	,N12783,N12784,N12785,N12786,N12788,N12789,N12791,N12792 
	,N12793,N12794,N12796,N12797,N12798,N12799,N12800,N12801 
	,N12802,N12803,N12804,N12805,N12806,N12807,N12808,N12809 
	,N12810,N12813,N12814,N12815,N12816,N12817,N12819,N12820 
	,N12821,N12822,N12823,N12824,N12825,N12826,N12828,N12829 
	,N12830,N12831,N12832,N12833,N12834,N12835,N12836,N12837 
	,N12838,N12839,N12840,N12841,N12842,N12843,N12844,N12846 
	,N12847,N12848,N12849,N12850,N12851,N12852,N12854,N12856 
	,N12857,N12858,N12859,N12860,N12862,N12863,N12864,N12865 
	,N12866,N12867,N12868,N12869,N12870,N12871,N12872,N12874 
	,N12875,N14515,N14520,N14521,N14522,N14525,N14526,N14528 
	,N14529,N14530,N14531,N14534,N14535,N14536,N14537,N14541 
	,N14542,N14543,N14545,N14550,N14551,N14554,N14555,N14556 
	,N14557,N14558,N14562,N14563,N14564,N14565,N14566,N14571 
	,N14572,N14577,N14578,N14579,N14580,N14582,N14583,N14585 
	,N14586,N14587,N14588,N14589,N14590,N14594,N14595,N14596 
	,N14599,N14600,N14601,N14602,N14604,N14605,N14607,N14608 
	,N14609,N14610,N14614,N14615,N14616,N14617,N14619,N14620 
	,N14621,N14622,N14623,N14625,N14627,N14628,N14629,N14630 
	,N14631,N14634,N14635,N14638,N14640,N14641,N14643,N14644 
	,N14645,N14646,N14649,N14650,N14651,N14652,N14653,N14655 
	,N14658,N14660,N14661,N14662,N14663,N14665,N14666,N14667 
	,N14669,N14671,N14672,N14673,N14679,N14680,N14682,N14683 
	,N14687,N14688,N14689,N14690,N14692,N14693,N14694,N14697 
	,N14699,N14700,N14701,N14703,N14704,N14706,N14707,N14710 
	,N14711,N14712,N14714,N14716,N14718,N14719,N14722,N14724 
	,N14725,N14728,N14729,N14733,N14736,N14737,N14738,N14739 
	,N14745,N14746,N14749,N14750,N14751,N14752,N14753,N14756 
	,N14758,N14759,N14760,N14761,N14763,N14767,N14768,N14771 
	,N14772,N14773,N14774,N14775,N14777,N14779,N14780,N14782 
	,N14783,N14787,N14788,N14789,N14792,N14794,N14795,N14797 
	,N14799,N14801,N14802,N14803,N14807,N14808,N14810,N14812 
	,N14813,N14814,N14817,N14821,N14822,N14823,N14824,N14826 
	,N14827,N14830,N14832,N14834,N14836,N14837,N14838,N14840 
	,N14841,N14843,N14845,N14846,N14847,N14849,N14853,N14855 
	,N14856,N14858,N14859,N14861,N14865,N14866,N14867,N14869 
	,N14871,N14872,N14874,N14875,N14877,N14878,N14881,N14882 
	,N14883,N14885,N14886,N14887,N14888,N14893,N14895,N14896 
	,N14897,N14899,N14900,N14902,N14903,N14904,N14908,N14909 
	,N14910,N14911,N14914,N14915,N14918,N14922,N14923,N14924 
	,N14927,N14928,N14929,N14931,N14934,N14935,N14938,N14940 
	,N14943,N14944,N14945,N14948,N14949,N14950,N14951,N14954 
	,N14956,N14957,N14958,N14959,N14963,N14964,N14965,N14966 
	,N14967,N14970,N14971,N14972,N14974,N14975,N14977,N14978 
	,N14979,N14980,N14982,N14985,N14986,N14987,N14988,N14990 
	,N14992,N14994,N14998,N14999,N15000,N15001,N15003,N15006 
	,N15010,N15011,N15012,N15014,N15015,N15016,N15020,N15022 
	,N15023,N15024,N15025,N15028,N15031,N15033,N15034,N15036 
	,N15038,N15039,N15040,N15041,N15043,N15045,N15048,N15050 
	,N15052,N15055,N15057,N15058,N15059,N15061,N15063,N15066 
	,N15067,N15069,N15070,N15072,N15074,N15075,N15076,N15079 
	,N15080,N15083,N15084,N15087,N15088,N15089,N15737,N15744 
	,N15746,N15749,N15763,N15767,N15769,N15771,N15773,N15777 
	,N15780,N15784,N15788,N15790,N15794,N15796,N15798,N15804 
	,N15829,N15832,N15839,N15854,N15863,N15867,N15891,N15898 
	,N15911,N15913,N15917,N15920,N15921,N15923,N15926,N15928 
	,N15931,N15934,N15935,N15937,N15938,N15941,N15944,N15945 
	,N15946,N15949,N15950,N15952,N15953,N15954,N15956,N15958 
	,N15959,N15960,N15962,N15963,N15967,N15969,N15970,N15972 
	,N15976,N15978,N15980,N15982,N15983,N15984,N15987,N15989 
	,N15990,N15992,N15994,N15996,N16062,N16063,N16065,N16069 
	,N16072,N16087,N16090,N16091,N16092,N16093,N16096,N16098 
	,N16099,N16100,N16103,N16104,N16105,N16107,N16108,N16109 
	,N16111,N16113,N16114,N16115,N16118,N16119,N16120,N16121 
	,N16124,N16125,N16126,N16129,N16130,N16131,N16132,N16133 
	,N16136,N16138,N16139,N16140,N16142,N16144,N16145,N16146 
	,N16147,N16150,N16151,N16153,N16154,N16155,N16158,N16159 
	,N16161,N16162,N16163,N16166,N16168,N16169,N16170,N16172 
	,N16175,N16176,N16178,N16180,N16181,N16182,N16183,N16186 
	,N16187,N16188,N16189,N16192,N16195,N16196,N16197,N16200 
	,N16201,N16202,N16203,N16206,N16207,N16208,N16212,N16213 
	,N16214,N16216,N16218,N16219,N16220,N16221,N16222,N16225 
	,N16228,N16229,N16230,N16231,N16234,N16235,N16236,N16239 
	,N16240,N16241,N16391,N16405,N16422,N16426,N16436,N16449 
	,N16452,N16468,N16482,N16530,N16532,N16534,N16535,N16540 
	,N16542,N16545,N16547,N16556,N16557,N16558,N16560,N16563 
	,N16565,N16568,N16570,N16572,N16575,N16576,N16578,N16607 
	,N16612,N16646,N22540,N22553,N22556,N22561,N22566,N22567 
	,N22568,N22572,N22573,N22574,N22577,N22578,N22579,N22580 
	,N22581,N22582,N22583,N22584,N22585,N22586,N22587,N22588 
	,N22589,N22590,N22592,N22593,N22595,N22596,N22597,N22598 
	,N22599,N22600,N22602,N22608,N22635,N22642,N22651,N22659 
	,N22699,N22705,N22714,N22721,N22732,N22738,N22746,N22752 
	,N22759,N43233,N43236,N43240,N43242,N43245,N43246,N43251 
	,N43255,N43261,N43262,N43266,N43267,N43268,N43271,N43280 
	,N43285,N43287,N43288,N43289,N43335,N43337,N43345,N43346 
	,N43353,N43361,N43365,N43367,N43395,N43396,N43404,N43412 
	,N43414,N43424,N43426,N43432,N43433,N43434,N43438,N43441 
	,N43446,N43448,N43449,N43467,N43470,N43473,N43474,N43477 
	,N43481,N43482,N43485,N43488,N43489,N43492,N43495,N43498 
	,N43503,N43506,N43511,N43514,N43517,N43520,N43523,N43526 
	,N43527,N43530,N43689,N43693,N43696,N43706,N43708,N43713 
	,N43715,N43717,N43739,N43743,N43747,N43755,N43757,N43761 
	,N43769,N43770,N43775,N43800,N43804,N43808,N43811,N43813 
	,N43817,N43831,N43834,N43837,N43838,N43841,N43845,N43846 
	,N43849,N43852,N43853,N43856,N43859,N43862,N43867,N43870 
	,N43875,N43878,N43881,N43884,N43887,N43890,N43891,N43894 
	,N43935,N43938,N43941,N43944,N43947,N43949,N43954,N43957 
	,N43960,N43963,N43964,N43967,N43970,N43973,N43976,N43982 
	,N43985,N43987,N43990,N43993,N43994,N43997,N44036,N44043 
	,N44049,N44056,N44063,N44070,N44079,N44087,N44095,N44103 
	,N44110,N44116,N44122,N44129;
INVX2 inst_blk01_cellmath__39_I440 (.Y(N5580), .A(a_man[0]));
CLKINVX12 inst_blk01_cellmath__39_I441 (.Y(N5560), .A(a_man[1]));
CLKINVX6 inst_blk01_cellmath__39_I442 (.Y(N5956), .A(a_man[2]));
CLKINVX4 inst_blk01_cellmath__39_I443 (.Y(N5551), .A(a_man[3]));
CLKINVX8 inst_blk01_cellmath__39_I444 (.Y(N5833), .A(a_man[4]));
CLKINVX6 inst_blk01_cellmath__39_I445 (.Y(N6212), .A(a_man[5]));
CLKINVX6 inst_blk01_cellmath__39_I446 (.Y(N5760), .A(a_man[6]));
BUFX2 inst_blk01_cellmath__39_I10021 (.Y(N22553), .A(N5760));
CLKINVX6 inst_blk01_cellmath__39_I447 (.Y(N6105), .A(a_man[7]));
CLKINVX4 inst_blk01_cellmath__39_I448 (.Y(N5612), .A(a_man[8]));
CLKINVX6 inst_blk01_cellmath__39_I449 (.Y(N5993), .A(a_man[9]));
INVX12 inst_blk01_cellmath__39_I450 (.Y(N5496), .A(a_man[10]));
INVX3 inst_blk01_cellmath__39_I451 (.Y(N5878), .A(a_man[11]));
INVX3 inst_blk01_cellmath__39_I452 (.Y(N5399), .A(a_man[12]));
CLKINVX6 inst_blk01_cellmath__39_I453 (.Y(N5761), .A(a_man[13]));
CLKINVX4 inst_blk01_cellmath__39_I454 (.Y(N6147), .A(a_man[14]));
INVX2 inst_blk01_cellmath__39_I455 (.Y(N5659), .A(a_man[15]));
INVX3 inst_blk01_cellmath__39_I456 (.Y(N6040), .A(a_man[16]));
INVX3 inst_blk01_cellmath__39_I457 (.Y(N5541), .A(a_man[17]));
INVX2 inst_blk01_cellmath__39_I458 (.Y(N5926), .A(a_man[18]));
INVX2 inst_blk01_cellmath__39_I459 (.Y(N5437), .A(a_man[19]));
INVX2 inst_blk01_cellmath__39_I460 (.Y(N5816), .A(a_man[20]));
INVX2 inst_blk01_cellmath__39_I461 (.Y(N6190), .A(a_man[21]));
INVX1 inst_blk01_cellmath__39_I462 (.Y(N5703), .A(a_man[22]));
BUFX2 inst_blk01_cellmath__39_I463 (.Y(N5934), .A(N5703));
XNOR2X1 inst_blk01_cellmath__39_I464 (.Y(N5815), .A(a_man[9]), .B(a_man[2]));
OR2XL inst_blk01_cellmath__39_I465 (.Y(N6009), .A(a_man[9]), .B(a_man[2]));
ADDFX1 inst_blk01_cellmath__39_I466 (.CO(N5891), .S(N5705), .A(a_man[3]), .B(a_man[10]), .CI(N5560));
ADDFXL inst_blk01_cellmath__39_I467 (.CO(N5411), .S(N6088), .A(a_man[4]), .B(a_man[11]), .CI(N5956));
ADDFX1 inst_blk01_cellmath__39_I468 (.CO(N5781), .S(N5592), .A(a_man[5]), .B(a_man[12]), .CI(N5551));
ADDFX1 inst_blk01_cellmath__39_I469 (.CO(N6160), .S(N5972), .A(a_man[6]), .B(a_man[13]), .CI(N5833));
XNOR2X1 inst_blk01_cellmath__39_I470 (.Y(N5484), .A(a_man[14]), .B(a_man[7]));
OR2XL inst_blk01_cellmath__39_I471 (.Y(N5674), .A(a_man[14]), .B(a_man[7]));
ADDHX1 inst_blk01_cellmath__39_I472 (.CO(N5556), .S(N6241), .A(N6212), .B(N5580));
XNOR2X1 inst_blk01_cellmath__39_I473 (.Y(N5746), .A(a_man[15]), .B(a_man[8]));
OR2XL inst_blk01_cellmath__39_I474 (.Y(N5941), .A(a_man[15]), .B(a_man[8]));
ADDFHXL inst_blk01_cellmath__39_I475 (.CO(N5829), .S(N5642), .A(N5760), .B(N5496), .CI(N5560));
XNOR2X1 inst_blk01_cellmath__39_I476 (.Y(N6025), .A(a_man[16]), .B(a_man[9]));
OR2XL inst_blk01_cellmath__39_I477 (.Y(N6209), .A(a_man[16]), .B(a_man[9]));
ADDFXL inst_blk01_cellmath__39_I478 (.CO(N6100), .S(N5909), .A(a_man[0]), .B(N5956), .CI(N6105));
ADDHX1 inst_blk01_cellmath__39_I479 (.CO(N5610), .S(N5425), .A(N5703), .B(N5878));
XNOR2X1 inst_blk01_cellmath__39_I480 (.Y(N5795), .A(a_man[17]), .B(a_man[10]));
OR2XL inst_blk01_cellmath__39_I481 (.Y(N5990), .A(a_man[17]), .B(a_man[10]));
ADDFXL inst_blk01_cellmath__39_I482 (.CO(N5876), .S(N5687), .A(N5551), .B(a_man[1]), .CI(N5612));
ADDHX1 inst_blk01_cellmath__39_I483 (.CO(N5397), .S(N6066), .A(N5399), .B(N5816));
ADDFX1 inst_blk01_cellmath__39_I484 (.CO(N5758), .S(N5574), .A(a_man[11]), .B(a_man[18]), .CI(a_man[2]));
ADDFHXL inst_blk01_cellmath__39_I485 (.CO(N6145), .S(N5955), .A(N5993), .B(N5761), .CI(N5833));
OR2XL inst_blk01_cellmath__39_I487 (.Y(N5656), .A(a_man[19]), .B(a_man[12]));
OR2XL inst_blk01_cellmath__39_I491 (.Y(N5434), .A(a_man[20]), .B(a_man[13]));
ADDFHX1 inst_blk01_cellmath__39_I494 (.CO(N6085), .S(N5889), .A(a_man[14]), .B(a_man[21]), .CI(a_man[0]));
ADDFHXL inst_blk01_cellmath__39_I495 (.CO(N5590), .S(N5408), .A(a_man[5]), .B(a_man[2]), .CI(N6105));
ADDHX1 inst_blk01_cellmath__39_I496 (.CO(N5969), .S(N5775), .A(N5399), .B(N6040));
XNOR2X1 inst_blk01_cellmath__39_I497 (.Y(N6156), .A(a_man[22]), .B(a_man[15]));
OR2XL inst_blk01_cellmath__39_I498 (.Y(N5478), .A(a_man[22]), .B(a_man[15]));
ADDFX1 inst_blk01_cellmath__39_I499 (.CO(N6237), .S(N6054), .A(a_man[3]), .B(a_man[1]), .CI(a_man[6]));
ADDFX1 inst_blk01_cellmath__39_I505 (.CO(N5905), .S(N5715), .A(a_man[4]), .B(a_man[18]), .CI(a_man[6]));
ADDHX1 inst_blk01_cellmath__39_I506 (.CO(N5421), .S(N6097), .A(a_man[9]), .B(N5878));
ADDFX1 inst_blk01_cellmath__39_I507 (.CO(N5792), .S(N5605), .A(a_man[5]), .B(a_man[19]), .CI(a_man[7]));
ADDHX1 inst_blk01_cellmath__39_I508 (.CO(N6173), .S(N5985), .A(a_man[10]), .B(N5399));
ADDFX1 inst_blk01_cellmath__39_I509 (.CO(N5683), .S(N5491), .A(a_man[6]), .B(a_man[20]), .CI(a_man[8]));
ADDHX1 inst_blk01_cellmath__39_I510 (.CO(N6064), .S(N5872), .A(N5761), .B(a_man[11]));
ADDFX1 inst_blk01_cellmath__39_I511 (.CO(N5571), .S(N6252), .A(a_man[7]), .B(a_man[21]), .CI(a_man[9]));
XNOR2X1 inst_blk01_cellmath__39_I512 (.Y(N5754), .A(a_man[22]), .B(a_man[8]));
OR2XL inst_blk01_cellmath__39_I513 (.Y(N5951), .A(a_man[22]), .B(a_man[8]));
XNOR2X1 inst_blk01_cellmath__39_I514 (.Y(N5651), .A(a_man[5]), .B(N5580));
OR2XL inst_blk01_cellmath__39_I515 (.Y(N5840), .A(a_man[5]), .B(N5580));
ADDFX1 inst_blk01_cellmath__39_I516 (.CO(N5726), .S(N5534), .A(N5560), .B(a_man[6]), .CI(N5659));
ADDFX1 inst_blk01_cellmath__39_I517 (.CO(N6113), .S(N5919), .A(a_man[0]), .B(a_man[7]), .CI(N5956));
ADDHX1 inst_blk01_cellmath__39_I518 (.CO(N5620), .S(N5431), .A(N5761), .B(N6040));
ADDFX1 inst_blk01_cellmath__39_I519 (.CO(N6001), .S(N5808), .A(a_man[1]), .B(a_man[8]), .CI(N5551));
ADDFX1 inst_blk01_cellmath__39_I520 (.CO(N5505), .S(N6183), .A(N5541), .B(N5878), .CI(N6147));
ADDFX1 inst_blk01_cellmath__39_I521 (.CO(N5886), .S(N5695), .A(N5580), .B(N5926), .CI(N5833));
ADDFX1 inst_blk01_cellmath__39_I522 (.CO(N5404), .S(N6079), .A(N5815), .B(N5659), .CI(N5399));
ADDFX1 inst_blk01_cellmath__39_I523 (.CO(N5770), .S(N5585), .A(N6040), .B(N5437), .CI(N6212));
ADDFX1 inst_blk01_cellmath__39_I524 (.CO(N6152), .S(N5961), .A(N6009), .B(N5705), .CI(N5761));
ADDFX1 inst_blk01_cellmath__39_I525 (.CO(N5664), .S(N5473), .A(N22553), .B(N5816), .CI(N5541));
ADDFXL inst_blk01_cellmath__39_I526 (.CO(N6047), .S(N5851), .A(N6147), .B(N5891), .CI(N6088));
ADDFX1 inst_blk01_cellmath__39_I527 (.CO(N5549), .S(N6231), .A(N6190), .B(N5926), .CI(N6105));
ADDFXL inst_blk01_cellmath__39_I528 (.CO(N5932), .S(N5740), .A(N5411), .B(N5659), .CI(N5592));
ADDFX1 inst_blk01_cellmath__39_I529 (.CO(N5445), .S(N6126), .A(N5437), .B(N5934), .CI(N5612));
ADDFHXL inst_blk01_cellmath__39_I530 (.CO(N5820), .S(N5632), .A(N5781), .B(N6040), .CI(N5972));
ADDFX1 inst_blk01_cellmath__39_I531 (.CO(N6199), .S(N6014), .A(N5541), .B(N5816), .CI(N5993));
ADDFX1 inst_blk01_cellmath__39_I532 (.CO(N5711), .S(N5517), .A(N5484), .B(N6160), .CI(N6241));
ADDFX1 inst_blk01_cellmath__39_I533 (.CO(N6093), .S(N5900), .A(N5926), .B(N6190), .CI(N5674));
ADDFX1 inst_blk01_cellmath__39_I534 (.CO(N5600), .S(N5417), .A(N5746), .B(N5556), .CI(N5642));
ADDFHXL inst_blk01_cellmath__39_I535 (.CO(N5980), .S(N5788), .A(N5941), .B(N5437), .CI(N5829));
ADDFX1 inst_blk01_cellmath__39_I536 (.CO(N5488), .S(N6169), .A(N6025), .B(N5425), .CI(N5909));
ADDHX1 inst_blk01_cellmath__39_I27980 (.CO(N5700), .S(N43517), .A(N5878), .B(N5659));
ADDFXL inst_blk01_cellmath__39_I27979 (.CO(N6188), .S(N43488), .A(a_man[4]), .B(a_man[1]), .CI(N5760));
ADDHX1 inst_blk01_cellmath__39_I28121 (.CO(N5522), .S(N43881), .A(N5496), .B(a_man[8]));
ADDFX1 inst_blk01_cellmath__39_I553 (.CO(N5847), .S(N5661), .A(N5522), .B(N5816), .CI(N6040));
ADDFX1 inst_blk01_cellmath__39_I28120 (.CO(N6021), .S(N43852), .A(a_man[3]), .B(a_man[17]), .CI(a_man[5]));
ADDFX1 inst_blk01_cellmath__39_I554 (.CO(N6227), .S(N6043), .A(N6097), .B(N6021), .CI(N5715));
ADDFX1 inst_blk01_cellmath__39_I555 (.CO(N5736), .S(N5544), .A(N5421), .B(N6190), .CI(N5541));
ADDFX1 inst_blk01_cellmath__39_I556 (.CO(N6123), .S(N5929), .A(N5905), .B(N5985), .CI(N5605));
ADDFX1 inst_blk01_cellmath__39_I557 (.CO(N5627), .S(N5441), .A(N5934), .B(N5926), .CI(N6173));
ADDFXL inst_blk01_cellmath__39_I558 (.CO(N6011), .S(N5818), .A(N5872), .B(N5792), .CI(N5491));
ADDFX1 inst_blk01_cellmath__39_I559 (.CO(N5514), .S(N6193), .A(N5437), .B(a_man[12]), .CI(N6147));
ADDFX1 inst_blk01_cellmath__39_I560 (.CO(N5895), .S(N5708), .A(N5683), .B(N6064), .CI(N6252));
ADDFX1 inst_blk01_cellmath__39_I561 (.CO(N5414), .S(N6090), .A(a_man[13]), .B(a_man[10]), .CI(N5659));
ADDFX1 inst_blk01_cellmath__39_I562 (.CO(N5783), .S(N5595), .A(N5754), .B(N5571), .CI(N5816));
ADDFX1 inst_blk01_cellmath__39_I563 (.CO(N6163), .S(N5975), .A(a_man[11]), .B(a_man[9]), .CI(a_man[14]));
ADDFX1 inst_blk01_cellmath__39_I564 (.CO(N5676), .S(N5485), .A(N5951), .B(N6190), .CI(N6040));
ADDFX1 inst_blk01_cellmath__39_I565 (.CO(N6059), .S(N5862), .A(a_man[12]), .B(a_man[10]), .CI(a_man[15]));
ADDHX1 inst_blk01_cellmath__39_I566 (.CO(N5558), .S(N6243), .A(N5541), .B(N5934));
ADDFX1 inst_blk01_cellmath__39_I567 (.CO(N5944), .S(N5748), .A(a_man[13]), .B(a_man[11]), .CI(a_man[16]));
XNOR2X1 inst_blk01_cellmath__39_I568 (.Y(N6132), .A(a_man[12]), .B(a_man[14]));
OR2XL inst_blk01_cellmath__39_I569 (.Y(N5454), .A(a_man[12]), .B(a_man[14]));
XNOR2X1 inst_blk01_cellmath__39_I570 (.Y(N6028), .A(a_man[13]), .B(a_man[15]));
OR2XL inst_blk01_cellmath__39_I571 (.Y(N6211), .A(a_man[13]), .B(a_man[15]));
XNOR2X1 inst_blk01_cellmath__39_I572 (.Y(N5912), .A(a_man[14]), .B(a_man[16]));
OR2XL inst_blk01_cellmath__39_I573 (.Y(N6103), .A(a_man[14]), .B(a_man[16]));
XNOR2X1 inst_blk01_cellmath__39_I574 (.Y(N5798), .A(a_man[15]), .B(a_man[17]));
OR2XL inst_blk01_cellmath__39_I575 (.Y(N5992), .A(a_man[15]), .B(a_man[17]));
INVXL inst_blk01_cellmath__39_I576 (.Y(N5577), .A(N22553));
ADDHX1 inst_blk01_cellmath__39_I577 (.CO(N5658), .S(N5464), .A(N5833), .B(N6105));
ADDHX1 inst_blk01_cellmath__39_I578 (.CO(N6039), .S(N5845), .A(N6212), .B(N5612));
ADDFX1 inst_blk01_cellmath__39_I579 (.CO(N5538), .S(N6225), .A(a_man[0]), .B(N5993), .CI(N22553));
ADDFX1 inst_blk01_cellmath__39_I580 (.CO(N5924), .S(N5731), .A(N6105), .B(a_man[1]), .CI(N5496));
ADDFX1 inst_blk01_cellmath__39_I581 (.CO(N5436), .S(N6120), .A(a_man[2]), .B(N5878), .CI(N5612));
ADDFX1 inst_blk01_cellmath__39_I582 (.CO(N5813), .S(N5624), .A(N5399), .B(a_man[3]), .CI(N5993));
ADDFX1 inst_blk01_cellmath__39_I583 (.CO(N6189), .S(N6007), .A(N5761), .B(a_man[4]), .CI(N5496));
ADDFX1 inst_blk01_cellmath__39_I584 (.CO(N5702), .S(N5510), .A(N5878), .B(N6147), .CI(N5612));
ADDFX1 inst_blk01_cellmath__39_I585 (.CO(N6086), .S(N5890), .A(N5399), .B(N5840), .CI(N5993));
ADDFX1 inst_blk01_cellmath__39_I586 (.CO(N5591), .S(N5409), .A(N5431), .B(N5726), .CI(N5496));
ADDFX1 inst_blk01_cellmath__39_I587 (.CO(N5970), .S(N5779), .A(N6113), .B(N5620), .CI(N5808));
ADDFX1 inst_blk01_cellmath__39_I588 (.CO(N5481), .S(N6159), .A(N5505), .B(N6001), .CI(N5695));
ADDFX1 inst_blk01_cellmath__39_I589 (.CO(N5858), .S(N5672), .A(N5886), .B(N5585), .CI(N5404));
ADDFHXL inst_blk01_cellmath__39_I590 (.CO(N6239), .S(N6056), .A(N5770), .B(N5473), .CI(N6152));
ADDFXL inst_blk01_cellmath__39_I591 (.CO(N5744), .S(N5555), .A(N6231), .B(N5664), .CI(N6047));
ADDFXL inst_blk01_cellmath__39_I592 (.CO(N6130), .S(N5939), .A(N6126), .B(N5549), .CI(N5932));
ADDFHXL inst_blk01_cellmath__39_I593 (.CO(N5640), .S(N5451), .A(N6014), .B(N5445), .CI(N5820));
ADDFX1 inst_blk01_cellmath__39_I594 (.CO(N6023), .S(N5826), .A(N5900), .B(N6199), .CI(N5711));
ADDFHXL inst_blk01_cellmath__39_I595 (.CO(N5523), .S(N6207), .A(N6093), .B(N5788), .CI(N5600));
ADDFXL inst_blk01_cellmath__39_I27981 (.CO(N43495), .S(N5678), .A(N5610), .B(N6209), .CI(N6100));
ADDFXL inst_blk01_cellmath__39_I596 (.CO(N5907), .S(N5718), .A(N5678), .B(N5980), .CI(N5488));
XNOR2X1 inst_blk01_cellmath__39_I27978 (.Y(N43473), .A(a_man[20]), .B(a_man[13]));
ADDFX1 inst_blk01_cellmath__39_I27988 (.CO(N5914), .S(N43482), .A(N43473), .B(N43517), .CI(N43488));
ADDHX1 inst_blk01_cellmath__39_I27977 (.CO(N43526), .S(N43511), .A(N5496), .B(N6147));
ADDFHXL inst_blk01_cellmath__39_I27976 (.CO(N43498), .S(N43481), .A(a_man[3]), .B(a_man[0]), .CI(N6212));
ADDFX1 inst_blk01_cellmath__39_I27987 (.CO(N5530), .S(N43520), .A(N43526), .B(N5656), .CI(N43498));
ADDFXL inst_blk01_cellmath__39_I28122 (.CO(N43859), .S(N6108), .A(N5700), .B(N5434), .CI(N6188));
ADDFXL inst_blk01_cellmath__39_I600 (.CO(N5685), .S(N5493), .A(N5914), .B(N5530), .CI(N6108));
ADDFHXL inst_blk01_cellmath__39_I28118 (.CO(N43875), .S(N43862), .A(a_man[2]), .B(a_man[16]), .CI(a_man[4]));
ADDFXL inst_blk01_cellmath__39_I28128 (.CO(N5957), .S(N43884), .A(N5437), .B(N5659), .CI(N43875));
ADDFHXL inst_blk01_cellmath__39_I28119 (.CO(N43837), .S(N43890), .A(N6147), .B(a_man[7]), .CI(N5993));
ADDFX1 inst_blk01_cellmath__39_I28129 (.CO(N5468), .S(N43846), .A(N43837), .B(N43881), .CI(N43852));
ADDFXL inst_blk01_cellmath__39_I604 (.CO(N5460), .S(N6143), .A(N5661), .B(N5957), .CI(N5468));
ADDFHXL inst_blk01_cellmath__39_I605 (.CO(N5842), .S(N5654), .A(N5544), .B(N5847), .CI(N6227));
ADDFXL inst_blk01_cellmath__39_I606 (.CO(N6221), .S(N6036), .A(N5441), .B(N5736), .CI(N6123));
ADDFXL inst_blk01_cellmath__39_I607 (.CO(N5727), .S(N5535), .A(N5627), .B(N6193), .CI(N6011));
ADDFHXL inst_blk01_cellmath__39_I608 (.CO(N6115), .S(N5921), .A(N6090), .B(N5514), .CI(N5895));
ADDFX1 inst_blk01_cellmath__39_I609 (.CO(N5621), .S(N5433), .A(N5975), .B(N5414), .CI(N5783));
ADDFX1 inst_blk01_cellmath__39_I610 (.CO(N6004), .S(N5810), .A(N6243), .B(N6163), .CI(N5862));
ADDFX1 inst_blk01_cellmath__39_I611 (.CO(N5507), .S(N6185), .A(N5558), .B(N5926), .CI(N6059));
ADDFX1 inst_blk01_cellmath__39_I612 (.CO(N5887), .S(N5699), .A(N5437), .B(a_man[17]), .CI(N5944));
ADDFX1 inst_blk01_cellmath__39_I613 (.CO(N5406), .S(N6083), .A(a_man[18]), .B(N5816), .CI(N5454));
ADDFX1 inst_blk01_cellmath__39_I614 (.CO(N5773), .S(N5587), .A(N6190), .B(a_man[19]), .CI(N6211));
ADDFX1 inst_blk01_cellmath__39_I615 (.CO(N6155), .S(N5966), .A(N6103), .B(a_man[20]), .CI(N5934));
ADDFX1 inst_blk01_cellmath__39_I616 (.CO(N5668), .S(N5476), .A(a_man[21]), .B(a_man[18]), .CI(N6040));
ADDFX1 inst_blk01_cellmath__39_I617 (.CO(N6051), .S(N5854), .A(a_man[19]), .B(a_man[17]), .CI(a_man[22]));
INVXL inst_blk01_cellmath__39_I618 (.Y(N6235), .A(N5551));
ADDHX1 inst_blk01_cellmath__39_I619 (.CO(N5448), .S(N6128), .A(N5560), .B(N5833));
ADDHX1 inst_blk01_cellmath__39_I620 (.CO(N5823), .S(N5636), .A(N6212), .B(N5956));
ADDFX1 inst_blk01_cellmath__39_I621 (.CO(N6203), .S(N6019), .A(N5577), .B(N5580), .CI(N5551));
ADDFX1 inst_blk01_cellmath__39_I622 (.CO(N5714), .S(N5520), .A(N22553), .B(N5464), .CI(N5560));
ADDFX1 inst_blk01_cellmath__39_I623 (.CO(N6096), .S(N5904), .A(N5845), .B(N5658), .CI(N5956));
ADDFX1 inst_blk01_cellmath__39_I624 (.CO(N5603), .S(N5420), .A(N6039), .B(N5551), .CI(N6225));
ADDFX1 inst_blk01_cellmath__39_I625 (.CO(N5984), .S(N5791), .A(N5731), .B(N5538), .CI(N5833));
ADDFX1 inst_blk01_cellmath__39_I626 (.CO(N5490), .S(N6172), .A(N6120), .B(N5924), .CI(N6212));
ADDFXL inst_blk01_cellmath__39_I627 (.CO(N5871), .S(N5681), .A(N5624), .B(N5436), .CI(N22553));
ADDFX1 inst_blk01_cellmath__39_I628 (.CO(N6249), .S(N6063), .A(N6007), .B(N5813), .CI(N6105));
ADDFX1 inst_blk01_cellmath__39_I629 (.CO(N5753), .S(N5569), .A(N5651), .B(N6189), .CI(N5510));
ADDFX1 inst_blk01_cellmath__39_I630 (.CO(N6140), .S(N5950), .A(N5534), .B(N5702), .CI(N5890));
ADDFX1 inst_blk01_cellmath__39_I631 (.CO(N5650), .S(N5459), .A(N6086), .B(N5919), .CI(N5409));
ADDFX1 inst_blk01_cellmath__39_I632 (.CO(N6033), .S(N5839), .A(N5591), .B(N6183), .CI(N5779));
ADDFX1 inst_blk01_cellmath__39_I633 (.CO(N5533), .S(N6218), .A(N6079), .B(N5970), .CI(N6159));
ADDFXL inst_blk01_cellmath__39_I634 (.CO(N5917), .S(N5724), .A(N5961), .B(N5481), .CI(N5672));
ADDFHXL inst_blk01_cellmath__39_I635 (.CO(N5430), .S(N6111), .A(N5858), .B(N5851), .CI(N6056));
ADDFHXL inst_blk01_cellmath__39_I636 (.CO(N5806), .S(N5619), .A(N6239), .B(N5740), .CI(N5555));
ADDFXL inst_blk01_cellmath__39_I637 (.CO(N6182), .S(N6000), .A(N5744), .B(N5632), .CI(N5939));
ADDFXL inst_blk01_cellmath__39_I638 (.CO(N5693), .S(N5504), .A(N6130), .B(N5517), .CI(N5451));
ADDFX1 inst_blk01_cellmath__39_I639 (.CO(N6078), .S(N5885), .A(N5640), .B(N5417), .CI(N5826));
ADDFHXL inst_blk01_cellmath__39_I640 (.CO(N5583), .S(N5403), .A(N6023), .B(N6169), .CI(N6207));
ADDFXL inst_blk01_cellmath__39_I27982 (.CO(N43523), .S(N6061), .A(N5795), .B(N6066), .CI(N5687));
ADDFHX1 inst_blk01_cellmath__39_I641 (.CO(N5960), .S(N5768), .A(N5523), .B(N6061), .CI(N5718));
ADDFX1 inst_blk01_cellmath__39_I27984 (.CO(N43514), .S(N5946), .A(N5574), .B(N5876), .CI(N5955));
ADDFX1 inst_blk01_cellmath__39_I27983 (.CO(N43485), .S(N43470), .A(N5990), .B(N6190), .CI(N5397));
ADDFXL inst_blk01_cellmath__39_I27989 (.CO(N43527), .S(N6098), .A(N43495), .B(N43470), .CI(N43523));
ADDFHX1 inst_blk01_cellmath__39_I642 (.CO(N5471), .S(N6151), .A(N5907), .B(N5946), .CI(N6098));
ADDFHXL inst_blk01_cellmath__39_I27985 (.CO(N43477), .S(N43530), .A(N5758), .B(N5934), .CI(N6145));
XNOR2X1 inst_blk01_cellmath__39_I27975 (.Y(N43467), .A(a_man[19]), .B(a_man[12]));
ADDFHXL inst_blk01_cellmath__39_I27986 (.CO(N43506), .S(N43492), .A(N43511), .B(N43467), .CI(N43481));
ADDFHXL inst_blk01_cellmath__39_I27991 (.CO(N6174), .S(N43503), .A(N43477), .B(N43506), .CI(N43520));
ADDFX1 inst_blk01_cellmath__39_I28123 (.CO(N43887), .S(N5614), .A(N5408), .B(N5775), .CI(N5889));
ADDFXL inst_blk01_cellmath__39_I645 (.CO(N5739), .S(N5546), .A(N6174), .B(N5614), .CI(N5493));
ADDFXL inst_blk01_cellmath__39_I28117 (.CO(N43845), .S(N43831), .A(N5612), .B(N5541), .CI(N5761));
ADDFX1 inst_blk01_cellmath__39_I28125 (.CO(N43878), .S(N5499), .A(N6156), .B(N6054), .CI(N43831));
ADDFHXL inst_blk01_cellmath__39_I28124 (.CO(N43849), .S(N43834), .A(N5969), .B(N6085), .CI(N5590));
ADDFHXL inst_blk01_cellmath__39_I28130 (.CO(N43891), .S(N5874), .A(N43859), .B(N43834), .CI(N43887));
ADDFHX1 inst_blk01_cellmath__39_I646 (.CO(N6125), .S(N5931), .A(N5685), .B(N5499), .CI(N5874));
ADDFX1 inst_blk01_cellmath__39_I28126 (.CO(N43841), .S(N43894), .A(N5478), .B(N5926), .CI(N6237));
ADDFXL inst_blk01_cellmath__39_I28127 (.CO(N43870), .S(N43856), .A(N43862), .B(N43845), .CI(N43890));
ADDFXL inst_blk01_cellmath__39_I28132 (.CO(N5953), .S(N43867), .A(N43841), .B(N43884), .CI(N43870));
ADDFX1 inst_blk01_cellmath__39_I649 (.CO(N5516), .S(N6198), .A(N5953), .B(N6043), .CI(N6143));
ADDFHXL inst_blk01_cellmath__39_I650 (.CO(N5898), .S(N5710), .A(N5460), .B(N5929), .CI(N5654));
ADDFXL inst_blk01_cellmath__39_I651 (.CO(N5416), .S(N6091), .A(N5842), .B(N5818), .CI(N6036));
ADDFHXL inst_blk01_cellmath__39_I652 (.CO(N5787), .S(N5598), .A(N5708), .B(N6221), .CI(N5535));
ADDFHXL inst_blk01_cellmath__39_I653 (.CO(N6168), .S(N5977), .A(N5727), .B(N5595), .CI(N5921));
ADDFX1 inst_blk01_cellmath__39_I654 (.CO(N5677), .S(N5486), .A(N5433), .B(N5485), .CI(N6115));
ADDFX1 inst_blk01_cellmath__39_I655 (.CO(N6060), .S(N5866), .A(N5810), .B(N5676), .CI(N5621));
ADDFX1 inst_blk01_cellmath__39_I656 (.CO(N5562), .S(N6245), .A(N6185), .B(N5748), .CI(N6004));
ADDFX1 inst_blk01_cellmath__39_I657 (.CO(N5945), .S(N5749), .A(N5507), .B(N6132), .CI(N5699));
ADDFX1 inst_blk01_cellmath__39_I658 (.CO(N5455), .S(N6136), .A(N5887), .B(N6028), .CI(N6083));
ADDFX1 inst_blk01_cellmath__39_I659 (.CO(N5835), .S(N5645), .A(N5406), .B(N5912), .CI(N5587));
ADDFX1 inst_blk01_cellmath__39_I660 (.CO(N6213), .S(N6029), .A(N5773), .B(N5798), .CI(N5966));
ADDFX1 inst_blk01_cellmath__39_I661 (.CO(N5721), .S(N5528), .A(N5476), .B(N5992), .CI(N6155));
ADDFX1 inst_blk01_cellmath__39_I662 (.CO(N6107), .S(N5913), .A(N5668), .B(a_man[16]), .CI(N5854));
ADDFX1 inst_blk01_cellmath__39_I663 (.CO(N5613), .S(N5427), .A(a_man[20]), .B(a_man[18]), .CI(N6051));
ADDHX1 inst_blk01_cellmath__39_I664 (.CO(N5994), .S(N5802), .A(a_man[19]), .B(a_man[21]));
ADDHX1 inst_blk01_cellmath__39_I665 (.CO(N5497), .S(N6177), .A(a_man[20]), .B(a_man[22]));
NOR2XL inst_blk01_cellmath__39_I668 (.Y(N6148), .A(N5580), .B(N6235));
NAND2XL inst_blk01_cellmath__39_I669 (.Y(N5467), .A(N5580), .B(N6235));
NOR2XL inst_blk01_cellmath__39_I670 (.Y(N5660), .A(N5551), .B(N6128));
NOR2XL inst_blk01_cellmath__39_I672 (.Y(N6042), .A(N5448), .B(N5636));
NAND2XL inst_blk01_cellmath__39_I673 (.Y(N6226), .A(N5448), .B(N5636));
NOR2XL inst_blk01_cellmath__39_I674 (.Y(N5542), .A(N5823), .B(N6019));
NAND2XL inst_blk01_cellmath__39_I675 (.Y(N5734), .A(N5823), .B(N6019));
NOR2XL inst_blk01_cellmath__39_I676 (.Y(N5928), .A(N6203), .B(N5520));
NOR2XL inst_blk01_cellmath__39_I678 (.Y(N5439), .A(N5714), .B(N5904));
NAND2XL inst_blk01_cellmath__39_I679 (.Y(N5626), .A(N5714), .B(N5904));
NOR2XL inst_blk01_cellmath__39_I680 (.Y(N5817), .A(N6096), .B(N5420));
NAND2XL inst_blk01_cellmath__39_I681 (.Y(N6010), .A(N6096), .B(N5420));
NOR2XL inst_blk01_cellmath__39_I682 (.Y(N6192), .A(N5603), .B(N5791));
NAND2XL inst_blk01_cellmath__39_I683 (.Y(N5512), .A(N5603), .B(N5791));
NOR2XL inst_blk01_cellmath__39_I684 (.Y(N5707), .A(N5984), .B(N6172));
NOR2XL inst_blk01_cellmath__39_I686 (.Y(N6089), .A(N5490), .B(N5681));
NAND2XL inst_blk01_cellmath__39_I687 (.Y(N5413), .A(N5490), .B(N5681));
NOR2XL inst_blk01_cellmath__39_I688 (.Y(N5594), .A(N5871), .B(N6063));
NOR2XL inst_blk01_cellmath__39_I690 (.Y(N5973), .A(N6249), .B(N5569));
NAND2XL inst_blk01_cellmath__39_I691 (.Y(N6162), .A(N6249), .B(N5569));
NAND3XL inst_blk01_cellmath__39_I28160 (.Y(N6026), .A(N5560), .B(N5956), .C(N5580));
AOI21XL inst_blk01_cellmath__39_I694 (.Y(N6176), .A0(N5467), .A1(N6026), .B0(N6148));
AOI21XL inst_blk01_cellmath__39_I695 (.Y(N6068), .A0(N6226), .A1(N5660), .B0(N6042));
OAI2BB1X1 inst_blk01_cellmath__39_I10023 (.Y(N5398), .A0N(N5551), .A1N(N6128), .B0(N6226));
OAI21XL inst_blk01_cellmath__39_I697 (.Y(N5730), .A0(N5398), .A1(N6176), .B0(N6068));
AOI21XL inst_blk01_cellmath__39_I698 (.Y(N5778), .A0(N5734), .A1(N5730), .B0(N5542));
AOI21XL inst_blk01_cellmath__39_I699 (.Y(N5671), .A0(N5626), .A1(N5928), .B0(N5439));
OAI2BB1X1 inst_blk01_cellmath__39_I10024 (.Y(N5857), .A0N(N6203), .A1N(N5520), .B0(N5626));
OAI21X1 inst_blk01_cellmath__39_I701 (.Y(N5606), .A0(N5778), .A1(N5857), .B0(N5671));
INVXL gen2_alt_A_I28612 (.Y(N44036), .A(N6192));
OAI2BB1X1 gen2_alt_A_I28613 (.Y(N5503), .A0N(N5512), .A1N(N5817), .B0(N44036));
CLKAND2X2 inst_blk01_cellmath__39_I703 (.Y(N5692), .A(N5512), .B(N6010));
AOI21X2 inst_blk01_cellmath__39_I709 (.Y(N6081), .A0(N5606), .A1(N5692), .B0(N5503));
AOI21XL inst_blk01_cellmath__39_I710 (.Y(N5965), .A0(N5413), .A1(N5707), .B0(N6089));
OAI2BB1X1 inst_blk01_cellmath__39_I10026 (.Y(N6153), .A0N(N5984), .A1N(N6172), .B0(N5413));
AOI21XL inst_blk01_cellmath__39_I713 (.Y(N5852), .A0(N6162), .A1(N5594), .B0(N5973));
OAI2BB1X1 inst_blk01_cellmath__39_I10027 (.Y(N6050), .A0N(N5871), .A1N(N6063), .B0(N6162));
OA21X1 inst_blk01_cellmath__39_I719 (.Y(N5786), .A0(N5965), .A1(N6050), .B0(N5852));
OR2XL inst_blk01_cellmath__39_I720 (.Y(N5976), .A(N6050), .B(N6153));
OAI21X2 inst_blk01_cellmath__39_I724 (.Y(N5540), .A0(N5976), .A1(N6081), .B0(N5786));
NOR2XL inst_blk01_cellmath__39_I751 (.Y(N5927), .A(N5753), .B(N5950));
NAND2XL inst_blk01_cellmath__39_I752 (.Y(N6121), .A(N5753), .B(N5950));
NOR2XL inst_blk01_cellmath__39_I753 (.Y(N5438), .A(N6140), .B(N5459));
NOR2XL inst_blk01_cellmath__39_I755 (.Y(N5814), .A(N5650), .B(N5839));
NAND2XL inst_blk01_cellmath__39_I756 (.Y(N6008), .A(N5650), .B(N5839));
NOR2XL inst_blk01_cellmath__39_I757 (.Y(N6191), .A(N6033), .B(N6218));
NOR2XL inst_blk01_cellmath__39_I759 (.Y(N5704), .A(N5533), .B(N5724));
NAND2X1 inst_blk01_cellmath__39_I760 (.Y(N5893), .A(N5533), .B(N5724));
NOR2X1 inst_blk01_cellmath__39_I761 (.Y(N6087), .A(N5917), .B(N6111));
NAND2X2 inst_blk01_cellmath__39_I762 (.Y(N5410), .A(N5917), .B(N6111));
NOR2XL inst_blk01_cellmath__39_I763 (.Y(N5593), .A(N5430), .B(N5619));
NAND2X4 inst_blk01_cellmath__39_I764 (.Y(N5780), .A(N5430), .B(N5619));
NOR2X2 inst_blk01_cellmath__39_I765 (.Y(N5971), .A(N5806), .B(N6000));
NAND2XL inst_blk01_cellmath__39_I766 (.Y(N6161), .A(N5806), .B(N6000));
NOR2XL inst_blk01_cellmath__39_I767 (.Y(N5483), .A(N6182), .B(N5504));
NAND2X2 inst_blk01_cellmath__39_I768 (.Y(N5673), .A(N6182), .B(N5504));
NOR2X1 inst_blk01_cellmath__39_I769 (.Y(N5860), .A(N5693), .B(N5885));
NAND2X2 inst_blk01_cellmath__39_I770 (.Y(N6057), .A(N5693), .B(N5885));
NOR2X1 inst_blk01_cellmath__39_I771 (.Y(N6240), .A(N5403), .B(N6078));
NAND2X4 inst_blk01_cellmath__39_I772 (.Y(N5557), .A(N6078), .B(N5403));
NOR2X2 inst_blk01_cellmath__39_I773 (.Y(N5745), .A(N5583), .B(N5768));
NAND2X2 inst_blk01_cellmath__39_I774 (.Y(N5940), .A(N5583), .B(N5768));
NOR2X1 inst_blk01_cellmath__39_I775 (.Y(N6131), .A(N5960), .B(N6151));
NAND2X4 inst_blk01_cellmath__39_I776 (.Y(N5452), .A(N5960), .B(N6151));
ADDFHXL inst_blk01_cellmath__39_I27990 (.CO(N43489), .S(N43474), .A(N43485), .B(N43530), .CI(N43514));
ADDFHX1 inst_blk01_cellmath__39_I27992 (.CO(N5850), .S(N5663), .A(N43527), .B(N43492), .CI(N43474));
NOR2X2 inst_blk01_cellmath__39_I777 (.Y(N5641), .A(N5471), .B(N5663));
NAND2X2 inst_blk01_cellmath__39_I778 (.Y(N5830), .A(N5471), .B(N5663));
ADDFHXL inst_blk01_cellmath__39_I27993 (.CO(N6230), .S(N6046), .A(N43482), .B(N43489), .CI(N43503));
NOR2X1 inst_blk01_cellmath__39_I779 (.Y(N6024), .A(N5850), .B(N6046));
NAND2X4 inst_blk01_cellmath__39_I27994 (.Y(N6208), .A(N5850), .B(N6046));
NOR2X2 inst_blk01_cellmath__39_I781 (.Y(N5525), .A(N6230), .B(N5546));
NAND2X1 inst_blk01_cellmath__39_I782 (.Y(N5719), .A(N6230), .B(N5546));
NOR2X1 inst_blk01_cellmath__39_I783 (.Y(N5908), .A(N5739), .B(N5931));
NAND2X4 inst_blk01_cellmath__39_I784 (.Y(N6102), .A(N5739), .B(N5931));
ADDFHXL inst_blk01_cellmath__39_I28131 (.CO(N43853), .S(N43838), .A(N43894), .B(N43849), .CI(N43878));
ADDFHXL inst_blk01_cellmath__39_I28133 (.CO(N5631), .S(N5444), .A(N43856), .B(N43891), .CI(N43838));
NOR2X1 inst_blk01_cellmath__39_I785 (.Y(N5424), .A(N6125), .B(N5444));
NAND2X2 inst_blk01_cellmath__39_I786 (.Y(N5609), .A(N6125), .B(N5444));
ADDFHX1 inst_blk01_cellmath__39_I28134 (.CO(N6012), .S(N5819), .A(N43846), .B(N43853), .CI(N43867));
NOR2XL inst_blk01_cellmath__39_I787 (.Y(N5797), .A(N5819), .B(N5631));
NAND2X4 inst_blk01_cellmath__39_I28135 (.Y(N5989), .A(N5631), .B(N5819));
NOR2X2 inst_blk01_cellmath__39_I789 (.Y(N6175), .A(N6012), .B(N6198));
NAND2X2 inst_blk01_cellmath__39_I790 (.Y(N5494), .A(N6012), .B(N6198));
NOR2X1 inst_blk01_cellmath__39_I791 (.Y(N5686), .A(N5516), .B(N5710));
NAND2X4 inst_blk01_cellmath__39_I792 (.Y(N5875), .A(N5516), .B(N5710));
NOR2X1 inst_blk01_cellmath__39_I793 (.Y(N6067), .A(N5898), .B(N6091));
NAND2X2 inst_blk01_cellmath__39_I794 (.Y(N5396), .A(N5898), .B(N6091));
NOR2XL inst_blk01_cellmath__39_I795 (.Y(N5573), .A(N5416), .B(N5598));
NAND2X2 inst_blk01_cellmath__39_I796 (.Y(N5759), .A(N5416), .B(N5598));
NOR2X1 inst_blk01_cellmath__39_I797 (.Y(N5954), .A(N5787), .B(N5977));
NAND2X1 inst_blk01_cellmath__39_I798 (.Y(N6144), .A(N5787), .B(N5977));
NOR2XL inst_blk01_cellmath__39_I799 (.Y(N5463), .A(N6168), .B(N5486));
NAND2X2 inst_blk01_cellmath__39_I800 (.Y(N5655), .A(N6168), .B(N5486));
NOR2XL inst_blk01_cellmath__39_I801 (.Y(N5843), .A(N5677), .B(N5866));
NAND2XL inst_blk01_cellmath__39_I802 (.Y(N6037), .A(N5677), .B(N5866));
NOR2XL inst_blk01_cellmath__39_I803 (.Y(N6223), .A(N6245), .B(N6060));
NAND2X1 inst_blk01_cellmath__39_I804 (.Y(N5536), .A(N6245), .B(N6060));
NOR2XL inst_blk01_cellmath__39_I805 (.Y(N5729), .A(N5562), .B(N5749));
NAND2XL inst_blk01_cellmath__39_I806 (.Y(N5922), .A(N5562), .B(N5749));
NOR2XL inst_blk01_cellmath__39_I807 (.Y(N6117), .A(N5945), .B(N6136));
NAND2XL inst_blk01_cellmath__39_I808 (.Y(N5435), .A(N5945), .B(N6136));
NOR2XL inst_blk01_cellmath__39_I809 (.Y(N5623), .A(N5455), .B(N5645));
NAND2XL inst_blk01_cellmath__39_I810 (.Y(N5811), .A(N5455), .B(N5645));
NOR2XL inst_blk01_cellmath__39_I811 (.Y(N6006), .A(N5835), .B(N6029));
NAND2XL inst_blk01_cellmath__39_I812 (.Y(N6187), .A(N5835), .B(N6029));
NOR2XL inst_blk01_cellmath__39_I813 (.Y(N5508), .A(N6213), .B(N5528));
NAND2XL inst_blk01_cellmath__39_I814 (.Y(N5701), .A(N6213), .B(N5528));
NOR2XL inst_blk01_cellmath__39_I815 (.Y(N5888), .A(N5721), .B(N5913));
NAND2XL inst_blk01_cellmath__39_I816 (.Y(N6084), .A(N5721), .B(N5913));
NOR2XL inst_blk01_cellmath__39_I817 (.Y(N5407), .A(N5427), .B(N6107));
NAND2XL inst_blk01_cellmath__39_I818 (.Y(N5589), .A(N5427), .B(N6107));
NOR2XL inst_blk01_cellmath__39_I819 (.Y(N5774), .A(N5802), .B(N5613));
NAND2XL inst_blk01_cellmath__39_I820 (.Y(N5968), .A(N5802), .B(N5613));
NOR2XL inst_blk01_cellmath__39_I821 (.Y(N6158), .A(N5994), .B(N6177));
NAND2XL inst_blk01_cellmath__39_I822 (.Y(N5477), .A(N5994), .B(N6177));
NOR2XL inst_blk01_cellmath__39_I823 (.Y(N5670), .A(N6190), .B(N5497));
NAND2XL inst_blk01_cellmath__39_I824 (.Y(N5856), .A(N6190), .B(N5497));
NOR2XL inst_blk01_cellmath__39_I825 (.Y(N6053), .A(a_man[22]), .B(a_man[21]));
NAND2XL inst_blk01_cellmath__39_I826 (.Y(N6236), .A(a_man[22]), .B(a_man[21]));
AOI21X1 inst_blk01_cellmath__39_I827 (.Y(N5936), .A0(N6121), .A1(N5540), .B0(N5927));
AOI21XL inst_blk01_cellmath__39_I828 (.Y(N5825), .A0(N6008), .A1(N5438), .B0(N5814));
OAI2BB1X1 inst_blk01_cellmath__39_I10029 (.Y(N6020), .A0N(N6140), .A1N(N5459), .B0(N6008));
OAI21X2 inst_blk01_cellmath__39_I830 (.Y(N5604), .A0(N6020), .A1(N5936), .B0(N5825));
AOI21X1 inst_blk01_cellmath__39_I831 (.Y(N5492), .A0(N6191), .A1(N5893), .B0(N5704));
OAI2BB1X1 inst_blk01_cellmath__39_I10031 (.Y(N5682), .A0N(N6033), .A1N(N6218), .B0(N5893));
AOI21X2 inst_blk01_cellmath__39_I834 (.Y(N6251), .A0(N5780), .A1(N6087), .B0(N5593));
NAND2X4 inst_blk01_cellmath__39_I835 (.Y(N5570), .A(N5780), .B(N5410));
OAI21X4 inst_blk01_cellmath__39_I836 (.Y(N6034), .A0(N5570), .A1(N5492), .B0(N6251));
NOR2X4 inst_blk01_cellmath__39_I837 (.Y(N6220), .A(N5682), .B(N5570));
AOI21X2 inst_blk01_cellmath__39_I838 (.Y(N5918), .A0(N5673), .A1(N5971), .B0(N5483));
NAND2X2 inst_blk01_cellmath__39_I839 (.Y(N6112), .A(N6161), .B(N5673));
INVXL inst_blk01_cellmath__39_I840 (.Y(N5800), .A(N6057));
AOI21X4 inst_blk01_cellmath__39_I841 (.Y(N5807), .A0(N5860), .A1(N5557), .B0(N6240));
NAND2X4 inst_blk01_cellmath__39_I842 (.Y(N6002), .A(N6057), .B(N5557));
OAI21X4 inst_blk01_cellmath__39_I843 (.Y(N5584), .A0(N6002), .A1(N5918), .B0(N5807));
NOR2X4 inst_blk01_cellmath__39_I844 (.Y(N5769), .A(N6002), .B(N6112));
AOI21X4 inst_blk01_cellmath__39_I845 (.Y(N5472), .A0(N5452), .A1(N5745), .B0(N6131));
NAND2X4 inst_blk01_cellmath__39_I846 (.Y(N5665), .A(N5940), .B(N5452));
INVXL inst_blk01_cellmath__39_I847 (.Y(N5579), .A(N5830));
AOI21X4 inst_blk01_cellmath__39_I848 (.Y(N6232), .A0(N5641), .A1(N6208), .B0(N6024));
NAND2X4 inst_blk01_cellmath__39_I849 (.Y(N5548), .A(N6208), .B(N5830));
OAI21X4 inst_blk01_cellmath__39_I850 (.Y(N6013), .A0(N5548), .A1(N5472), .B0(N6232));
NOR2X6 inst_blk01_cellmath__39_I851 (.Y(N6200), .A(N5665), .B(N5548));
AOI21X4 inst_blk01_cellmath__39_I852 (.Y(N5899), .A0(N5525), .A1(N6102), .B0(N5908));
NAND2X2 inst_blk01_cellmath__39_I853 (.Y(N6092), .A(N5719), .B(N6102));
INVXL inst_blk01_cellmath__39_I854 (.Y(N5732), .A(N5609));
AOI21X2 inst_blk01_cellmath__39_I855 (.Y(N5789), .A0(N5989), .A1(N5424), .B0(N5797));
NAND2X4 inst_blk01_cellmath__39_I856 (.Y(N5979), .A(N5989), .B(N5609));
OAI21X4 inst_blk01_cellmath__39_I857 (.Y(N5564), .A0(N5979), .A1(N5899), .B0(N5789));
NOR2X6 inst_blk01_cellmath__39_I858 (.Y(N5751), .A(N5979), .B(N6092));
AOI21X4 inst_blk01_cellmath__39_I859 (.Y(N5457), .A0(N6175), .A1(N5875), .B0(N5686));
NAND2X4 inst_blk01_cellmath__39_I860 (.Y(N5646), .A(N5875), .B(N5494));
INVXL inst_blk01_cellmath__39_I861 (.Y(N5892), .A(N5396));
AOI21X2 inst_blk01_cellmath__39_I862 (.Y(N6214), .A0(N6067), .A1(N5759), .B0(N5573));
NAND2X4 inst_blk01_cellmath__39_I863 (.Y(N5529), .A(N5759), .B(N5396));
OAI21X4 inst_blk01_cellmath__39_I864 (.Y(N5996), .A0(N5529), .A1(N5457), .B0(N6214));
NOR2X4 inst_blk01_cellmath__39_I865 (.Y(N6178), .A(N5529), .B(N5646));
AOI21X2 inst_blk01_cellmath__39_I866 (.Y(N5880), .A0(N5655), .A1(N5954), .B0(N5463));
NAND2X2 inst_blk01_cellmath__39_I867 (.Y(N6073), .A(N5655), .B(N6144));
INVXL inst_blk01_cellmath__39_I868 (.Y(N5675), .A(N6037));
AOI21XL inst_blk01_cellmath__39_I869 (.Y(N5764), .A0(N5536), .A1(N5843), .B0(N6223));
NAND2X1 inst_blk01_cellmath__39_I870 (.Y(N5958), .A(N5536), .B(N6037));
OAI21X2 inst_blk01_cellmath__39_I871 (.Y(N5543), .A0(N5958), .A1(N5880), .B0(N5764));
NOR2X2 inst_blk01_cellmath__39_I872 (.Y(N5735), .A(N5958), .B(N6073));
AOI21X1 inst_blk01_cellmath__39_I873 (.Y(N5440), .A0(N5435), .A1(N5729), .B0(N6117));
NAND2X1 inst_blk01_cellmath__39_I874 (.Y(N5628), .A(N5435), .B(N5922));
INVXL inst_blk01_cellmath__39_I875 (.Y(N5453), .A(N5811));
AOI21XL inst_blk01_cellmath__39_I876 (.Y(N6195), .A0(N6187), .A1(N5623), .B0(N6006));
NAND2XL inst_blk01_cellmath__39_I877 (.Y(N5513), .A(N6187), .B(N5811));
OAI21XL inst_blk01_cellmath__39_I878 (.Y(N5974), .A0(N5513), .A1(N5440), .B0(N6195));
NOR2XL inst_blk01_cellmath__39_I879 (.Y(N6165), .A(N5513), .B(N5628));
AOI21XL inst_blk01_cellmath__39_I880 (.Y(N5863), .A0(N6084), .A1(N5508), .B0(N5888));
NAND2XL inst_blk01_cellmath__39_I881 (.Y(N6058), .A(N6084), .B(N5701));
INVXL inst_blk01_cellmath__39_I882 (.Y(N5910), .A(N5407));
INVXL inst_blk01_cellmath__39_I883 (.Y(N6101), .A(N5589));
AOI21XL inst_blk01_cellmath__39_I884 (.Y(N5747), .A0(N5968), .A1(N5407), .B0(N5774));
NAND2XL inst_blk01_cellmath__39_I885 (.Y(N5943), .A(N5968), .B(N5589));
INVXL inst_blk01_cellmath__39_I886 (.Y(N5796), .A(N5863));
INVXL inst_blk01_cellmath__39_I887 (.Y(N5991), .A(N6058));
OAI21XL inst_blk01_cellmath__39_I888 (.Y(N6027), .A0(N6101), .A1(N5863), .B0(N5910));
NOR2XL inst_blk01_cellmath__39_I889 (.Y(N6210), .A(N6101), .B(N6058));
OAI21XL inst_blk01_cellmath__39_I890 (.Y(N5526), .A0(N5943), .A1(N5863), .B0(N5747));
NOR2XL inst_blk01_cellmath__39_I891 (.Y(N5720), .A(N5943), .B(N6058));
AOI21XL inst_blk01_cellmath__39_I892 (.Y(N5688), .A0(N5701), .A1(N5974), .B0(N5508));
AOI21XL inst_blk01_cellmath__39_I893 (.Y(N6070), .A0(N5991), .A1(N5974), .B0(N5796));
AOI21XL inst_blk01_cellmath__39_I894 (.Y(N5576), .A0(N6210), .A1(N5974), .B0(N6027));
AOI21XL inst_blk01_cellmath__39_I895 (.Y(N5844), .A0(N5856), .A1(N6158), .B0(N5670));
NAND2XL inst_blk01_cellmath__39_I896 (.Y(N6038), .A(N5856), .B(N5477));
INVXL inst_blk01_cellmath__39_I897 (.Y(N5657), .A(N6236));
AO21XL inst_blk01_cellmath__39_I898 (.Y(N5776), .A0(N5720), .A1(N5974), .B0(N5526));
AND2X1 inst_blk01_cellmath__39_I899 (.Y(N5967), .A(N6165), .B(N5720));
INVXL inst_blk01_cellmath__39_I900 (.Y(N6157), .A(N5604));
AOI21X4 inst_blk01_cellmath__39_I901 (.Y(N5938), .A0(N5604), .A1(N6220), .B0(N6034));
AOI21X4 inst_blk01_cellmath__39_I902 (.Y(N5450), .A0(N5769), .A1(N6034), .B0(N5584));
NAND2X4 inst_blk01_cellmath__39_I903 (.Y(N5639), .A(N5769), .B(N6220));
AOI21X4 inst_blk01_cellmath__39_I904 (.Y(N5828), .A0(N6200), .A1(N5584), .B0(N6013));
NAND2X4 inst_blk01_cellmath__39_I905 (.Y(N6022), .A(N6200), .B(N5769));
AOI21X4 inst_blk01_cellmath__39_I906 (.Y(N6206), .A0(N5751), .A1(N6013), .B0(N5564));
NAND2X4 inst_blk01_cellmath__39_I907 (.Y(N5524), .A(N5751), .B(N6200));
AOI21X4 inst_blk01_cellmath__39_I908 (.Y(N5717), .A0(N6178), .A1(N5564), .B0(N5996));
NAND2X4 inst_blk01_cellmath__39_I909 (.Y(N5906), .A(N6178), .B(N5751));
AOI21X2 inst_blk01_cellmath__39_I910 (.Y(N6099), .A0(N5735), .A1(N5996), .B0(N5543));
NAND2X2 inst_blk01_cellmath__39_I911 (.Y(N5422), .A(N5735), .B(N6178));
AOI21X2 inst_blk01_cellmath__39_I912 (.Y(N5607), .A0(N5967), .A1(N5543), .B0(N5776));
NAND2X2 inst_blk01_cellmath__39_I913 (.Y(N5794), .A(N5967), .B(N5735));
INVXL inst_blk01_cellmath__39_I914 (.Y(N5479), .A(N6157));
INVX1 inst_blk01_cellmath__39_I915 (.Y(N5669), .A(N5938));
OAI21X4 inst_blk01_cellmath__39_I916 (.Y(N5873), .A0(N5639), .A1(N6157), .B0(N5450));
OAI21X4 inst_blk01_cellmath__39_I917 (.Y(N5394), .A0(N5938), .A1(N6022), .B0(N5828));
OAI21X1 inst_blk01_cellmath__39_I918 (.Y(N5757), .A0(N5524), .A1(N5450), .B0(N6206));
NOR2X1 inst_blk01_cellmath__39_I919 (.Y(N5952), .A(N5524), .B(N5639));
OAI21X2 inst_blk01_cellmath__39_I920 (.Y(N6142), .A0(N5906), .A1(N5828), .B0(N5717));
NOR2X2 inst_blk01_cellmath__39_I921 (.Y(N5461), .A(N5906), .B(N6022));
OAI21X2 inst_blk01_cellmath__39_I922 (.Y(N5653), .A0(N5422), .A1(N6206), .B0(N6099));
NOR2X2 inst_blk01_cellmath__39_I923 (.Y(N5841), .A(N5422), .B(N5524));
OAI21X4 inst_blk01_cellmath__39_I924 (.Y(N6035), .A0(N5794), .A1(N5717), .B0(N5607));
NOR2X2 inst_blk01_cellmath__39_I925 (.Y(N6222), .A(N5794), .B(N5906));
INVXL inst_blk01_cellmath__39_I928 (.Y(N6238), .A(N5873));
AOI21X4 inst_blk01_cellmath__39_I931 (.Y(N5698), .A0(N5461), .A1(N5669), .B0(N6142));
AOI21X4 inst_blk01_cellmath__39_I932 (.Y(N6082), .A0(N5841), .A1(N5873), .B0(N5653));
AOI21X4 inst_blk01_cellmath__39_I933 (.Y(N5588), .A0(N6222), .A1(N5394), .B0(N6035));
NOR2XL inst_blk01_cellmath__39_I938 (.Y(N6075), .A(N5800), .B(N5918));
NOR2XL inst_blk01_cellmath__39_I939 (.Y(N5986), .A(N6075), .B(N5860));
NOR2XL inst_blk01_cellmath__39_I940 (.Y(N5737), .A(N5579), .B(N5472));
NOR2XL inst_blk01_cellmath__39_I941 (.Y(N6253), .A(N5737), .B(N5641));
NOR2XL andori2bb1_A_I28614 (.Y(N44043), .A(N5732), .B(N5899));
NOR2XL andori2bb1_A_I28615 (.Y(N5652), .A(N44043), .B(N5424));
NOR2X1 inst_blk01_cellmath__39_I944 (.Y(N5784), .A(N5892), .B(N5457));
NOR2XL inst_blk01_cellmath__39_I945 (.Y(N5920), .A(N6067), .B(N5784));
NOR2XL inst_blk01_cellmath__39_I946 (.Y(N6244), .A(N5675), .B(N5880));
NOR2XL inst_blk01_cellmath__39_I947 (.Y(N6184), .A(N6244), .B(N5843));
NOR2XL inst_blk01_cellmath__39_I948 (.Y(N5831), .A(N5453), .B(N5440));
NOR2XL inst_blk01_cellmath__39_I949 (.Y(N5586), .A(N5831), .B(N5623));
INVXL inst_blk01_cellmath__39_I950 (.Y(N5962), .A(N5974));
NOR2XL inst_blk01_cellmath__39_I951 (.Y(N5426), .A(N5657), .B(N5844));
NOR2XL inst_blk01_cellmath__39_I952 (.Y(N5633), .A(N5426), .B(N6053));
OR2XL inst_blk01_cellmath__39_I953 (.Y(N5821), .A(N5657), .B(N6038));
NAND2BXL inst_blk01_cellmath__39_I964 (.Y(N6228), .AN(N6240), .B(N5557));
NAND2BXL inst_blk01_cellmath__39_I965 (.Y(N6242), .AN(N5745), .B(N5940));
NAND2BXL inst_blk01_cellmath__39_I966 (.Y(N5942), .AN(N6131), .B(N5452));
NAND2BXL inst_blk01_cellmath__39_I967 (.Y(N6164), .AN(N5641), .B(N5830));
NAND2BXL inst_blk01_cellmath__39_I968 (.Y(N5643), .AN(N6024), .B(N6208));
NAND2BXL inst_blk01_cellmath__39_I969 (.Y(N5911), .AN(N5525), .B(N5719));
NAND2BXL inst_blk01_cellmath__39_I970 (.Y(N5611), .AN(N5908), .B(N6102));
NAND2BXL inst_blk01_cellmath__39_I971 (.Y(N5578), .AN(N5424), .B(N5609));
NAND2BXL inst_blk01_cellmath__39_I972 (.Y(N5925), .AN(N5797), .B(N5989));
NAND2BXL inst_blk01_cellmath__39_I974 (.Y(N6146), .AN(N5686), .B(N5875));
NAND2BXL inst_blk01_cellmath__39_I975 (.Y(N5859), .AN(N6067), .B(N5396));
NAND2BXL inst_blk01_cellmath__39_I976 (.Y(N6205), .AN(N5573), .B(N5759));
NAND2BXL inst_blk01_cellmath__39_I977 (.Y(N6119), .AN(N5954), .B(N6144));
NAND2BXL inst_blk01_cellmath__39_I978 (.Y(N5812), .AN(N5463), .B(N5655));
NAND2BXL inst_blk01_cellmath__39_I979 (.Y(N6141), .AN(N5843), .B(N6037));
NAND2BXL inst_blk01_cellmath__39_I980 (.Y(N5622), .AN(N6223), .B(N5536));
NAND2BXL inst_blk01_cellmath__39_I981 (.Y(N5777), .AN(N5729), .B(N5922));
NAND2BXL inst_blk01_cellmath__39_I982 (.Y(N5480), .AN(N6117), .B(N5435));
NAND2BXL inst_blk01_cellmath__39_I983 (.Y(N5552), .AN(N5623), .B(N5811));
NAND2BXL inst_blk01_cellmath__39_I984 (.Y(N5903), .AN(N6006), .B(N6187));
NAND2BXL inst_blk01_cellmath__39_I985 (.Y(N6250), .AN(N5508), .B(N5701));
NAND2BXL inst_blk01_cellmath__39_I986 (.Y(N5725), .AN(N5888), .B(N6084));
NAND2BXL inst_blk01_cellmath__39_I987 (.Y(N6077), .AN(N5407), .B(N5589));
NAND2BXL inst_blk01_cellmath__39_I988 (.Y(N5547), .AN(N5774), .B(N5968));
NAND2BXL inst_blk01_cellmath__39_I989 (.Y(N5987), .AN(N6158), .B(N5477));
NAND2BXL inst_blk01_cellmath__39_I990 (.Y(N5684), .AN(N5670), .B(N5856));
NAND2BXL inst_blk01_cellmath__39_I991 (.Y(N5487), .AN(N6053), .B(N6236));
XNOR2X1 inst_blk01_cellmath__39_I997 (.Y(N609), .A(N6242), .B(N6238));
INVX1 inst_cellmath__48_I27883 (.Y(N5554), .A(N5394));
XNOR2X1 inst_blk01_cellmath__39_I998 (.Y(N613), .A(N5911), .B(N5554));
XNOR2X1 inst_blk01_cellmath__39_I1000 (.Y(N621), .A(N6119), .B(N5698));
XNOR2X1 inst_blk01_cellmath__39_I1001 (.Y(N625), .A(N5777), .B(N6082));
XNOR2X1 inst_blk01_cellmath__39_I1002 (.Y(N633), .A(N5987), .B(N5588));
XOR2XL inst_blk01_cellmath__39_I1021 (.Y(N5475), .A(N6228), .B(N5986));
OAI21XL inst_blk01_cellmath__39_I1022 (.Y(N5848), .A0(N5800), .A1(N6112), .B0(N5986));
XNOR2X1 inst_blk01_cellmath__39_I1023 (.Y(N5667), .A(N6228), .B(N5848));
MXI2XL inst_blk01_cellmath__39_I1024 (.Y(N608), .A(N5475), .B(N5667), .S0(N5669));
XNOR2X1 inst_blk01_cellmath__39_I1025 (.Y(N6234), .A(N5940), .B(N5942));
XNOR2X1 inst_blk01_cellmath__39_I1026 (.Y(N6049), .A(N5745), .B(N5942));
MXI2XL inst_blk01_cellmath__39_I1027 (.Y(N610), .A(N6234), .B(N6049), .S0(N6238));
XOR2XL inst_blk01_cellmath__39_I1028 (.Y(N5742), .A(N5472), .B(N6164));
NAND2XL inst_blk01_cellmath__39_I1029 (.Y(N5785), .A(N5665), .B(N5472));
XNOR2X1 inst_blk01_cellmath__39_I1030 (.Y(N5935), .A(N6164), .B(N5785));
MXI2XL inst_blk01_cellmath__39_I1031 (.Y(N611), .A(N5935), .B(N5742), .S0(N6238));
XOR2XL inst_blk01_cellmath__39_I1032 (.Y(N5447), .A(N5643), .B(N6253));
OAI21XL inst_blk01_cellmath__39_I1033 (.Y(N6133), .A0(N5579), .A1(N5665), .B0(N6253));
INVXL xnor2_A_I28616 (.Y(N44049), .A(N5643));
MXI2XL xnor2_A_I28617 (.Y(N5635), .A(N5643), .B(N44049), .S0(N6133));
MXI2XL inst_blk01_cellmath__39_I1035 (.Y(N612), .A(N5635), .B(N5447), .S0(N6238));
NAND2XL inst_blk01_cellmath__39_I1040 (.Y(N6069), .A(N6092), .B(N5899));
OAI21X1 inst_blk01_cellmath__39_I1044 (.Y(N5539), .A0(N6092), .A1(N5732), .B0(N5652));
XNOR2X1 inst_blk01_cellmath__39_I1047 (.Y(N6171), .A(N6146), .B(N5494));
XNOR2X1 inst_blk01_cellmath__39_I1048 (.Y(N5983), .A(N6146), .B(N6175));
AOI21X2 inst_cellmath__48_I27884 (.Y(N6186), .A0(N5952), .A1(N5479), .B0(N5757));
MXI2XL inst_blk01_cellmath__39_I1049 (.Y(N618), .A(N6171), .B(N5983), .S0(N6186));
XOR2XL inst_blk01_cellmath__39_I1050 (.Y(N5680), .A(N5859), .B(N5457));
NAND2XL inst_blk01_cellmath__39_I1051 (.Y(N5482), .A(N5646), .B(N5457));
XNOR2X1 inst_blk01_cellmath__39_I1052 (.Y(N5869), .A(N5859), .B(N5482));
MXI2XL inst_blk01_cellmath__39_I1053 (.Y(N619), .A(N5869), .B(N5680), .S0(N6186));
XOR2XL inst_blk01_cellmath__39_I1054 (.Y(N6248), .A(N6205), .B(N5920));
OAI21XL inst_blk01_cellmath__39_I1055 (.Y(N5827), .A0(N5892), .A1(N5646), .B0(N5920));
XNOR2X1 inst_blk01_cellmath__39_I1056 (.Y(N5568), .A(N6205), .B(N5827));
MXI2X1 inst_blk01_cellmath__39_I1057 (.Y(N620), .A(N5568), .B(N6248), .S0(N6186));
XNOR2X1 inst_blk01_cellmath__39_I1058 (.Y(N6139), .A(N6144), .B(N5812));
XNOR2X1 inst_blk01_cellmath__39_I1059 (.Y(N5948), .A(N5812), .B(N5954));
MXI2X1 inst_blk01_cellmath__39_I1060 (.Y(N622), .A(N6139), .B(N5948), .S0(N5698));
XOR2XL inst_blk01_cellmath__39_I1061 (.Y(N5648), .A(N5880), .B(N6141));
NAND2XL inst_blk01_cellmath__39_I1062 (.Y(N5756), .A(N6073), .B(N5880));
XNOR2X1 inst_blk01_cellmath__39_I1063 (.Y(N5838), .A(N6141), .B(N5756));
MXI2X1 inst_blk01_cellmath__39_I1064 (.Y(N623), .A(N5838), .B(N5648), .S0(N5698));
XOR2XL inst_blk01_cellmath__39_I1065 (.Y(N6216), .A(N6184), .B(N5622));
OAI21XL inst_blk01_cellmath__39_I1066 (.Y(N6116), .A0(N5675), .A1(N6073), .B0(N6184));
XNOR2X1 inst_blk01_cellmath__39_I1067 (.Y(N5532), .A(N5622), .B(N6116));
MXI2X1 inst_blk01_cellmath__39_I1068 (.Y(N624), .A(N5532), .B(N6216), .S0(N5698));
XNOR2X1 inst_blk01_cellmath__39_I1069 (.Y(N6110), .A(N5480), .B(N5922));
XNOR2X1 inst_blk01_cellmath__39_I1070 (.Y(N5916), .A(N5480), .B(N5729));
MXI2X1 inst_blk01_cellmath__39_I1071 (.Y(N626), .A(N6110), .B(N5916), .S0(N6082));
XOR2XL inst_blk01_cellmath__39_I1072 (.Y(N5618), .A(N5552), .B(N5440));
NAND2XL inst_blk01_cellmath__39_I1073 (.Y(N6052), .A(N5628), .B(N5440));
XNOR2X1 inst_blk01_cellmath__39_I1074 (.Y(N5805), .A(N5552), .B(N6052));
MXI2XL inst_blk01_cellmath__39_I1075 (.Y(N627), .A(N5805), .B(N5618), .S0(N6082));
XOR2XL inst_blk01_cellmath__39_I1076 (.Y(N6181), .A(N5903), .B(N5586));
OAI21XL inst_blk01_cellmath__39_I1077 (.Y(N5521), .A0(N5453), .A1(N5628), .B0(N5586));
XNOR2X1 inst_blk01_cellmath__39_I1078 (.Y(N5501), .A(N5903), .B(N5521));
MXI2XL inst_blk01_cellmath__39_I1079 (.Y(N628), .A(N5501), .B(N6181), .S0(N6082));
XOR2XL inst_blk01_cellmath__39_I1080 (.Y(N5884), .A(N6250), .B(N5962));
NAND2BXL inst_blk01_cellmath__39_I1081 (.Y(N5870), .AN(N6165), .B(N5962));
XNOR2X1 inst_blk01_cellmath__39_I1082 (.Y(N6076), .A(N6250), .B(N5870));
MXI2XL inst_blk01_cellmath__39_I1083 (.Y(N629), .A(N6076), .B(N5884), .S0(N6082));
XOR2XL inst_blk01_cellmath__39_I1084 (.Y(N5582), .A(N5725), .B(N5688));
OAI2BB1X1 inst_blk01_cellmath__39_I1085 (.Y(N6219), .A0N(N5701), .A1N(N6165), .B0(N5688));
XNOR2X1 inst_blk01_cellmath__39_I1086 (.Y(N5766), .A(N5725), .B(N6219));
MXI2XL inst_blk01_cellmath__39_I1087 (.Y(N630), .A(N5766), .B(N5582), .S0(N6082));
XOR2XL inst_blk01_cellmath__39_I1088 (.Y(N6150), .A(N6077), .B(N6070));
OAI2BB1X1 inst_blk01_cellmath__39_I1089 (.Y(N5694), .A0N(N5991), .A1N(N6165), .B0(N6070));
XNOR2X1 inst_blk01_cellmath__39_I1090 (.Y(N5469), .A(N6077), .B(N5694));
MXI2X1 inst_blk01_cellmath__39_I1091 (.Y(N631), .A(N5469), .B(N6150), .S0(N6082));
XOR2XL inst_blk01_cellmath__39_I1092 (.Y(N5849), .A(N5547), .B(N5576));
OAI2BB1X1 inst_blk01_cellmath__39_I1093 (.Y(N6045), .A0N(N6210), .A1N(N6165), .B0(N5576));
XNOR2X1 inst_blk01_cellmath__39_I1094 (.Y(N6044), .A(N5547), .B(N6045));
MXI2X1 inst_blk01_cellmath__39_I1095 (.Y(N632), .A(N6044), .B(N5849), .S0(N6082));
XNOR2X1 inst_blk01_cellmath__39_I1096 (.Y(N5738), .A(N5684), .B(N5477));
XNOR2X1 inst_blk01_cellmath__39_I1097 (.Y(N5545), .A(N5684), .B(N6158));
MXI2X1 inst_blk01_cellmath__39_I1098 (.Y(N634), .A(N5738), .B(N5545), .S0(N5588));
XOR2XL inst_blk01_cellmath__39_I1099 (.Y(N6124), .A(N5487), .B(N5844));
NAND2XL inst_blk01_cellmath__39_I1100 (.Y(N5978), .A(N6038), .B(N5844));
XNOR2X1 inst_blk01_cellmath__39_I1101 (.Y(N5442), .A(N5487), .B(N5978));
MXI2X1 inst_blk01_cellmath__39_I1102 (.Y(N635), .A(N5442), .B(N6124), .S0(N5588));
OA21XL inst_blk01_cellmath__39_I1103 (.Y(N637), .A0(N5821), .A1(N5588), .B0(N5633));
INVXL inst_blk01_cellmath__39_I1104 (.Y(N636), .A(N637));
INVXL inst_cellmath__42_0_I1107 (.Y(N7100), .A(a_exp[2]));
INVXL inst_cellmath__42_0_I1108 (.Y(N7107), .A(a_exp[3]));
INVXL inst_cellmath__48_I27903 (.Y(N7103), .A(a_exp[1]));
OAI21XL inst_cellmath__42_0_I1109 (.Y(N7102), .A0(N7100), .A1(N7103), .B0(N7107));
NOR2XL inst_cellmath__42_0_I1112 (.Y(N7108), .A(N7100), .B(N7103));
XOR2X4 inst_cellmath__42_0_I1114 (.Y(inst_cellmath__42[4]), .A(a_exp[4]), .B(N7102));
MXI2XL inst_cellmath__48_I1125 (.Y(N7163), .A(N609), .B(N608), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1126 (.Y(N7219), .A(N610), .B(N609), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1127 (.Y(N7275), .A(N611), .B(N610), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1128 (.Y(N7331), .A(N612), .B(N611), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1129 (.Y(N7132), .A(N613), .B(N612), .S0(a_exp[0]));
XNOR2X1 inst_cellmath__48_I27890 (.Y(N43267), .A(N5719), .B(N5611));
XNOR2X1 inst_cellmath__48_I27891 (.Y(N43280), .A(N5525), .B(N5611));
MXI2XL inst_cellmath__48_I27892 (.Y(N614), .A(N43267), .B(N43280), .S0(N5554));
MXI2XL inst_cellmath__48_I1130 (.Y(N7187), .A(N614), .B(N613), .S0(a_exp[0]));
XNOR2X1 inst_cellmath__48_I27897 (.Y(N43240), .A(N5925), .B(N5539));
XOR2XL inst_cellmath__48_I27896 (.Y(N43285), .A(N5925), .B(N5652));
MXI2X1 inst_cellmath__48_I27902 (.Y(N616), .A(N43240), .B(N43285), .S0(N5554));
XNOR2X1 inst_cellmath__48_I27894 (.Y(N43262), .A(N5578), .B(N6069));
XOR2XL inst_cellmath__48_I27893 (.Y(N43246), .A(N5899), .B(N5578));
MXI2XL inst_cellmath__48_I27895 (.Y(N615), .A(N43262), .B(N43246), .S0(N5554));
MXI2XL inst_cellmath__48_I1132 (.Y(N7298), .A(N616), .B(N615), .S0(a_exp[0]));
NAND2BXL inst_cellmath__48_I27885 (.Y(N43242), .AN(N6175), .B(N5494));
XNOR2X1 inst_cellmath__48_I27889 (.Y(N617), .A(N43242), .B(N6186));
MXI2XL inst_cellmath__48_I1134 (.Y(N7154), .A(N618), .B(N617), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1135 (.Y(N7210), .A(N619), .B(N618), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1136 (.Y(N7266), .A(N620), .B(N619), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1137 (.Y(N7322), .A(N621), .B(N620), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1138 (.Y(N7124), .A(N622), .B(N621), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1139 (.Y(N7176), .A(N623), .B(N622), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1140 (.Y(N7234), .A(N624), .B(N623), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1141 (.Y(N7289), .A(N625), .B(N624), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1142 (.Y(N7346), .A(N626), .B(N625), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1143 (.Y(N7147), .A(N627), .B(N626), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1144 (.Y(N7203), .A(N628), .B(N627), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1145 (.Y(N7256), .A(N629), .B(N628), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1146 (.Y(N7311), .A(N630), .B(N629), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1147 (.Y(N7367), .A(N631), .B(N630), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1148 (.Y(N7168), .A(N632), .B(N631), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1149 (.Y(N7225), .A(N633), .B(N632), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1150 (.Y(N7281), .A(N634), .B(N633), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1151 (.Y(N7335), .A(N635), .B(N634), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1152 (.Y(N7136), .A(N636), .B(N635), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1153 (.Y(N7192), .A(N637), .B(N636), .S0(a_exp[0]));
NAND2XL inst_cellmath__48_I1154 (.Y(N7248), .A(a_exp[0]), .B(N637));
NAND2XL inst_cellmath__48_I27886 (.Y(N43236), .A(N43242), .B(N6186));
OR2XL inst_cellmath__48_I28173 (.Y(N43289), .A(N43242), .B(N6186));
NOR2BX1 inst_cellmath__48_I28175 (.Y(N43266), .AN(N43240), .B(N5554));
INVXL inst_cellmath__48_I27904 (.Y(inst_cellmath__42[1]), .A(N7103));
MX2XL inst_cellmath__48_I28176 (.Y(N43261), .A(N43267), .B(N43280), .S0(N5554));
NOR2BX1 inst_cellmath__48_I27908 (.Y(N43287), .AN(a_exp[0]), .B(N43261));
MX2XL inst_cellmath__48_I28177 (.Y(N43255), .A(N43262), .B(N43246), .S0(N5554));
NOR2X1 inst_cellmath__48_I27912 (.Y(N43245), .A(a_exp[0]), .B(N43255));
MXI2XL inst_cellmath__48_I27913 (.Y(N7243), .A(N615), .B(N614), .S0(a_exp[0]));
INVXL inst_cellmath__48_I27914 (.Y(N43288), .A(a_exp[0]));
AOI211XL inst_cellmath__48_I28178 (.Y(N43251), .A0(N5554), .A1(N43285), .B0(N43288), .C0(N43266));
AOI21X1 inst_cellmath__48_I27916 (.Y(N43268), .A0(N43236), .A1(N43289), .B0(a_exp[0]));
MXI2XL inst_cellmath__48_I27917 (.Y(N7354), .A(N616), .B(N617), .S0(N43288));
BUFX6 inst_cellmath__48_I27918 (.Y(N7336), .A(inst_cellmath__42[1]));
NOR3BXL inst_cellmath__48_I28179 (.Y(N43271), .AN(N7336), .B(N43268), .C(N43251));
NOR3XL inst_cellmath__48_I27921 (.Y(N43233), .A(N7336), .B(N43245), .C(N43287));
NOR2XL inst_cellmath__48_I27922 (.Y(N7287), .A(N43233), .B(N43271));
MXI2XL inst_cellmath__48_I1162 (.Y(N7209), .A(N7163), .B(N7275), .S0(N7336));
MXI2XL inst_cellmath__48_I1163 (.Y(N7265), .A(N7219), .B(N7331), .S0(N7336));
MXI2XL inst_cellmath__48_I1164 (.Y(N7319), .A(N7275), .B(N7132), .S0(N7336));
MXI2XL inst_cellmath__48_I1165 (.Y(N7121), .A(N7331), .B(N7187), .S0(N7336));
MXI2XL inst_cellmath__48_I1166 (.Y(N7175), .A(N7132), .B(N7243), .S0(N7336));
MXI2XL inst_cellmath__48_I1167 (.Y(N7233), .A(N7187), .B(N7298), .S0(N7336));
MXI2XL inst_cellmath__48_I1169 (.Y(N7344), .A(N7298), .B(N7154), .S0(N7336));
MXI2XL inst_cellmath__48_I1170 (.Y(N7144), .A(N7354), .B(N7210), .S0(N7336));
MXI2XL inst_cellmath__48_I1171 (.Y(N7200), .A(N7154), .B(N7266), .S0(N7336));
MXI2X1 inst_cellmath__48_I1172 (.Y(N7255), .A(N7210), .B(N7322), .S0(N7336));
MXI2XL inst_cellmath__48_I1173 (.Y(N7310), .A(N7266), .B(N7124), .S0(N7336));
MXI2XL inst_cellmath__48_I1174 (.Y(N7365), .A(N7322), .B(N7176), .S0(N7336));
MXI2XL inst_cellmath__48_I1175 (.Y(N7166), .A(N7124), .B(N7234), .S0(N7336));
MXI2XL inst_cellmath__48_I1176 (.Y(N7222), .A(N7176), .B(N7289), .S0(N7336));
MXI2XL inst_cellmath__48_I1177 (.Y(N7278), .A(N7234), .B(N7346), .S0(N7336));
MXI2XL inst_cellmath__48_I1178 (.Y(N7334), .A(N7289), .B(N7147), .S0(N7336));
MXI2XL inst_cellmath__48_I1179 (.Y(N7135), .A(N7346), .B(N7203), .S0(N7336));
MXI2XL inst_cellmath__48_I1180 (.Y(N7190), .A(N7147), .B(N7256), .S0(N7336));
MXI2XL inst_cellmath__48_I1181 (.Y(N7246), .A(N7203), .B(N7311), .S0(N7336));
MXI2XL inst_cellmath__48_I1182 (.Y(N7301), .A(N7256), .B(N7367), .S0(N7336));
MXI2XL inst_cellmath__48_I1183 (.Y(N7357), .A(N7311), .B(N7168), .S0(N7336));
MXI2X1 inst_cellmath__48_I1184 (.Y(N7157), .A(N7367), .B(N7225), .S0(N7336));
MXI2X1 inst_cellmath__48_I1185 (.Y(N7213), .A(N7168), .B(N7281), .S0(N7336));
MXI2XL inst_cellmath__48_I1186 (.Y(N7270), .A(N7225), .B(N7335), .S0(N7336));
MXI2X1 inst_cellmath__48_I1187 (.Y(N7325), .A(N7281), .B(N7136), .S0(N7336));
MXI2XL inst_cellmath__48_I1188 (.Y(N7128), .A(N7335), .B(N7192), .S0(N7336));
MXI2X1 inst_cellmath__48_I1189 (.Y(N7181), .A(N7136), .B(N7248), .S0(N7336));
NOR2XL inst_cellmath__48_I1190 (.Y(N7239), .A(N7336), .B(N7192));
NOR2XL inst_cellmath__48_I1191 (.Y(N7350), .A(N7336), .B(N7248));
CLKMX2X4 inst_cellmath__48_I10039 (.Y(N7271), .A(N7103), .B(inst_cellmath__42[1]), .S0(N7100));
MXI2XL inst_cellmath__48_I1200 (.Y(N7309), .A(N7175), .B(N7209), .S0(N7271));
MXI2XL inst_cellmath__48_I1201 (.Y(N7364), .A(N7233), .B(N7265), .S0(N7271));
MXI2XL inst_cellmath__48_I1202 (.Y(N7165), .A(N7287), .B(N7319), .S0(N7271));
MXI2XL inst_cellmath__48_I1203 (.Y(N7220), .A(N7344), .B(N7121), .S0(N7271));
MXI2XL inst_cellmath__48_I1204 (.Y(N7276), .A(N7144), .B(N7175), .S0(N7271));
MXI2XL inst_cellmath__48_I1205 (.Y(N7333), .A(N7200), .B(N7233), .S0(N7271));
MXI2XL inst_cellmath__48_I1206 (.Y(N7134), .A(N7255), .B(N7287), .S0(N7271));
MXI2XL inst_cellmath__48_I1207 (.Y(N7189), .A(N7310), .B(N7344), .S0(N7271));
MXI2X1 inst_cellmath__48_I1208 (.Y(N7245), .A(N7365), .B(N7144), .S0(N7271));
INVXL mx2i_A_I28618 (.Y(N44056), .A(N7271));
AOI22XL mx2i_A_I28619 (.Y(N7299), .A0(N44056), .A1(N7166), .B0(N7200), .B1(N7271));
MXI2X1 inst_cellmath__48_I1210 (.Y(N7355), .A(N7222), .B(N7255), .S0(N7271));
MXI2X1 inst_cellmath__48_I1211 (.Y(N7156), .A(N7278), .B(N7310), .S0(N7271));
MXI2X1 inst_cellmath__48_I1212 (.Y(N7212), .A(N7334), .B(N7365), .S0(N7271));
MXI2XL inst_cellmath__48_I1213 (.Y(N7269), .A(N7135), .B(N7166), .S0(N7271));
MXI2XL inst_cellmath__48_I1214 (.Y(N7324), .A(N7190), .B(N7222), .S0(N7271));
MXI2XL inst_cellmath__48_I1215 (.Y(N7125), .A(N7246), .B(N7278), .S0(N7271));
MXI2XL inst_cellmath__48_I1216 (.Y(N7179), .A(N7301), .B(N7334), .S0(N7271));
MXI2XL inst_cellmath__48_I1217 (.Y(N7238), .A(N7357), .B(N7135), .S0(N7271));
MXI2X1 inst_cellmath__48_I1218 (.Y(N7292), .A(N7157), .B(N7190), .S0(N7271));
MXI2XL inst_cellmath__48_I1219 (.Y(N7349), .A(N7213), .B(N7246), .S0(N7271));
MXI2XL inst_cellmath__48_I1220 (.Y(N7149), .A(N7270), .B(N7301), .S0(N7271));
MXI2XL inst_cellmath__48_I1221 (.Y(N7204), .A(N7325), .B(N7357), .S0(N7271));
MXI2X1 inst_cellmath__48_I1222 (.Y(N7259), .A(N7128), .B(N7157), .S0(N7271));
MXI2X1 inst_cellmath__48_I1223 (.Y(N7315), .A(N7181), .B(N7213), .S0(N7271));
MXI2XL inst_cellmath__48_I1224 (.Y(N7370), .A(N7239), .B(N7270), .S0(N7271));
MXI2XL inst_cellmath__48_I1225 (.Y(N7171), .A(N7350), .B(N7325), .S0(N7271));
NAND2XL inst_cellmath__48_I1226 (.Y(N7227), .A(N7271), .B(N7128));
NAND2XL inst_cellmath__48_I1227 (.Y(N7337), .A(N7181), .B(N7271));
NAND2XL inst_cellmath__48_I1228 (.Y(N7194), .A(N7271), .B(N7239));
NAND2XL inst_cellmath__48_I1229 (.Y(N7304), .A(N7350), .B(N7271));
MXI2XL inst_cellmath__48_I1240 (.Y(N7267), .A(N7309), .B(N7179), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I28180 (.Y(N7321), .A(N7364), .B(N7238), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1242 (.Y(N7123), .A(N7165), .B(N7292), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I1243 (.Y(N7178), .A(N7220), .B(N7349), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I1244 (.Y(N7236), .A(N7276), .B(N7149), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I1245 (.Y(N7290), .A(N7333), .B(N7204), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I1246 (.Y(N7347), .A(N7134), .B(N7259), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I1247 (.Y(N7146), .A(N7189), .B(N7315), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1248 (.Y(N7202), .A(N7245), .B(N7370), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1249 (.Y(N7258), .A(N7299), .B(N7171), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1250 (.Y(N7313), .A(N7355), .B(N7227), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1251 (.Y(N7368), .A(N7156), .B(N7337), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1252 (.Y(N7169), .A(N7212), .B(N7194), .S0(inst_cellmath__42[4]));
MXI2X1 inst_cellmath__48_I1253 (.Y(N7224), .A(N7269), .B(N7304), .S0(inst_cellmath__42[4]));
NOR2X1 inst_cellmath__48_I1254 (.Y(N7280), .A(inst_cellmath__42[4]), .B(N7324));
NOR2X1 inst_cellmath__48_I1255 (.Y(N7138), .A(inst_cellmath__42[4]), .B(N7125));
NOR2XL inst_cellmath__48_I1256 (.Y(N7249), .A(inst_cellmath__42[4]), .B(N7179));
NOR2XL inst_cellmath__48_I1257 (.Y(N7359), .A(inst_cellmath__42[4]), .B(N7238));
NOR2XL inst_cellmath__48_I1258 (.Y(N7215), .A(inst_cellmath__42[4]), .B(N7292));
NOR2XL inst_cellmath__48_I1259 (.Y(N7327), .A(inst_cellmath__42[4]), .B(N7349));
NOR2X1 inst_cellmath__48_I1260 (.Y(N7184), .A(inst_cellmath__42[4]), .B(N7149));
NOR2X1 inst_cellmath__48_I1261 (.Y(N7295), .A(inst_cellmath__42[4]), .B(N7204));
NOR2XL inst_cellmath__48_I1262 (.Y(N7152), .A(inst_cellmath__42[4]), .B(N7259));
NOR2X2 inst_cellmath__48_I1263 (.Y(N7263), .A(inst_cellmath__42[4]), .B(N7315));
NOR2XL inst_cellmath__48_I1264 (.Y(N7373), .A(inst_cellmath__42[4]), .B(N7370));
NOR2XL inst_cellmath__48_I1265 (.Y(N7230), .A(inst_cellmath__42[4]), .B(N7171));
NOR2XL inst_cellmath__48_I1266 (.Y(N7341), .A(inst_cellmath__42[4]), .B(N7227));
NOR2XL inst_cellmath__48_I1267 (.Y(N7197), .A(inst_cellmath__42[4]), .B(N7337));
NOR2X1 inst_cellmath__48_I1268 (.Y(N7307), .A(inst_cellmath__42[4]), .B(N7194));
NOR2XL inst_cellmath__48_I1269 (.Y(N7162), .A(inst_cellmath__42[4]), .B(N7304));
XOR2X4 inst_cellmath__48_I10040 (.Y(N7196), .A(N7107), .B(N7108));
MXI2XL inst_cellmath__48_I1277 (.Y(N7127), .A(N7202), .B(N7267), .S0(N7196));
MXI2X1 inst_cellmath__48_I1278 (.Y(N7182), .A(N7258), .B(N7321), .S0(N7196));
MXI2XL inst_cellmath__48_I1280 (.Y(N7293), .A(N7368), .B(N7178), .S0(N7196));
MXI2XL inst_cellmath__48_I1281 (.Y(N7352), .A(N7169), .B(N7236), .S0(N7196));
MXI2XL inst_cellmath__48_I1282 (.Y(N7151), .A(N7224), .B(N7290), .S0(N7196));
MXI2XL inst_cellmath__48_I1283 (.Y(N7206), .A(N7280), .B(N7347), .S0(N7196));
MXI2XL inst_cellmath__48_I1284 (.Y(N7261), .A(N7138), .B(N7146), .S0(N7196));
MXI2XL inst_cellmath__48_I1285 (.Y(N7316), .A(N7249), .B(N7202), .S0(N7196));
MXI2XL inst_cellmath__48_I1286 (.Y(N7371), .A(N7359), .B(N7258), .S0(N7196));
MXI2XL inst_cellmath__48_I1287 (.Y(N7173), .A(N7215), .B(N7313), .S0(N7196));
MXI2XL inst_cellmath__48_I1288 (.Y(N7229), .A(N7327), .B(N7368), .S0(N7196));
MXI2X1 inst_cellmath__48_I1289 (.Y(N7283), .A(N7184), .B(N7169), .S0(N7196));
MXI2X1 inst_cellmath__48_I1290 (.Y(N7339), .A(N7295), .B(N7224), .S0(N7196));
MXI2XL inst_cellmath__48_I1291 (.Y(N7140), .A(N7152), .B(N7280), .S0(N7196));
MXI2XL inst_cellmath__48_I1292 (.Y(N7195), .A(N7263), .B(N7138), .S0(N7196));
MXI2XL inst_cellmath__48_I1293 (.Y(N7252), .A(N7373), .B(N7249), .S0(N7196));
MXI2X1 inst_cellmath__48_I1294 (.Y(N7306), .A(N7230), .B(N7359), .S0(N7196));
INVXL mx2i_A_I28620 (.Y(N44063), .A(N7196));
AOI22XL mx2i_A_I28621 (.Y(N7361), .A0(N44063), .A1(N7341), .B0(N7215), .B1(N7196));
MXI2XL inst_cellmath__48_I1296 (.Y(N7160), .A(N7197), .B(N7327), .S0(N7196));
INVXL mx2i_A_I10810 (.Y(N22759), .A(N7196));
AOI22XL mx2i_A_I10811 (.Y(N7217), .A0(N7307), .A1(N22759), .B0(N7196), .B1(N7184));
MXI2XL inst_cellmath__48_I1298 (.Y(N7273), .A(N7162), .B(N7295), .S0(N7196));
NAND2XL inst_cellmath__48_I1299 (.Y(N7330), .A(N7152), .B(N7196));
NAND2XL inst_cellmath__48_I1301 (.Y(N7297), .A(N7373), .B(N7196));
MXI2X1 inst_cellmath__48_I27951 (.Y(N43414), .A(N7313), .B(N7123), .S0(N7196));
NOR2XL node_cs_const1_cs_A_I28622 (.Y(N44070), .A(a_exp[4]), .B(N7102));
XNOR2X1 node_cs_const1_cs_A_I28623 (.Y(N7131), .A(a_exp[5]), .B(N44070));
NOR2X1 inst_cellmath__48_I27953 (.Y(N43404), .A(N7131), .B(N43414));
NAND3BX4 inst_cellmath__48_I27954 (.Y(N43412), .AN(N7131), .B(N7196), .C(N7263));
INVX3 inst_cellmath__48_I27955 (.Y(N7631), .A(N43412));
CLKXOR2X1 inst_cellmath__48_I27956 (.Y(inst_cellmath__61[2]), .A(N7631), .B(N43404));
INVX3 inst_cellmath__48_I27957 (.Y(N3661), .A(inst_cellmath__61[2]));
NOR2XL inst_cellmath__48_I1310 (.Y(N733), .A(N7131), .B(N7127));
NOR2X1 inst_cellmath__48_I1311 (.Y(N734), .A(N7131), .B(N7182));
NOR2XL inst_cellmath__48_I1313 (.Y(N736), .A(N7131), .B(N7293));
NOR2XL inst_cellmath__48_I1315 (.Y(N738), .A(N7131), .B(N7151));
NOR2XL inst_cellmath__48_I1316 (.Y(N739), .A(N7131), .B(N7206));
NOR2XL inst_cellmath__48_I1317 (.Y(N740), .A(N7131), .B(N7261));
NOR2XL inst_cellmath__48_I1318 (.Y(N741), .A(N7131), .B(N7316));
NOR2XL inst_cellmath__48_I1320 (.Y(N743), .A(N7131), .B(N7173));
NOR2XL inst_cellmath__48_I1321 (.Y(N744), .A(N7131), .B(N7229));
NOR2X1 inst_cellmath__48_I1322 (.Y(N745), .A(N7131), .B(N7283));
NOR2X1 inst_cellmath__48_I1323 (.Y(N746), .A(N7131), .B(N7339));
NOR2X1 inst_cellmath__48_I1324 (.Y(N747), .A(N7131), .B(N7140));
NOR2X1 inst_cellmath__48_I1325 (.Y(N748), .A(N7131), .B(N7195));
NOR2XL inst_cellmath__48_I1326 (.Y(N749), .A(N7131), .B(N7252));
NOR2X1 inst_cellmath__48_I1327 (.Y(N750), .A(N7131), .B(N7306));
NOR2XL inst_cellmath__48_I1328 (.Y(N751), .A(N7131), .B(N7361));
NOR2X1 inst_cellmath__48_I1329 (.Y(N752), .A(N7131), .B(N7160));
NOR2XL inst_cellmath__48_I1330 (.Y(N753), .A(N7131), .B(N7217));
NOR2X1 inst_cellmath__48_I1331 (.Y(N754), .A(N7131), .B(N7273));
NOR2XL inst_cellmath__48_I1332 (.Y(N755), .A(N7330), .B(N7131));
NOR2XL inst_cellmath__48_I1334 (.Y(N757), .A(N7297), .B(N7131));
CLKXOR2X1 cynw_cm_float_sin_I1339 (.Y(inst_cellmath__61[1]), .A(N7631), .B(N734));
CLKXOR2X1 cynw_cm_float_sin_I10513 (.Y(inst_cellmath__61[5]), .A(N7631), .B(N738));
CLKXOR2X1 cynw_cm_float_sin_I1344 (.Y(inst_cellmath__61[6]), .A(N7631), .B(N739));
CLKXOR2X1 cynw_cm_float_sin_I1348 (.Y(inst_cellmath__61[10]), .A(N7631), .B(N743));
CLKXOR2X1 cynw_cm_float_sin_I1349 (.Y(inst_cellmath__61[11]), .A(N7631), .B(N744));
CLKXOR2X1 cynw_cm_float_sin_I1350 (.Y(inst_cellmath__61[12]), .A(N7631), .B(N745));
CLKXOR2X1 cynw_cm_float_sin_I1351 (.Y(inst_cellmath__61[13]), .A(N7631), .B(N746));
CLKXOR2X1 cynw_cm_float_sin_I1352 (.Y(inst_cellmath__61[14]), .A(N7631), .B(N747));
CLKXOR2X1 cynw_cm_float_sin_I9898 (.Y(inst_cellmath__61[15]), .A(N7631), .B(N748));
CLKXOR2X1 cynw_cm_float_sin_I1355 (.Y(inst_cellmath__61[17]), .A(N7631), .B(N750));
CLKXOR2X1 cynw_cm_float_sin_I1356 (.Y(inst_cellmath__61[18]), .A(N7631), .B(N751));
CLKXOR2X1 cynw_cm_float_sin_I1357 (.Y(inst_cellmath__61[19]), .A(N7631), .B(N752));
CLKXOR2X1 cynw_cm_float_sin_I1358 (.Y(inst_cellmath__61[20]), .A(N7631), .B(N753));
CLKXOR2X1 cynw_cm_float_sin_I1359 (.Y(inst_cellmath__61[21]), .A(N7631), .B(N754));
CLKXOR2X1 cynw_cm_float_sin_I1360 (.Y(inst_cellmath__61[22]), .A(N7631), .B(N755));
INVX2 cynw_cm_float_sin_I296 (.Y(N3657), .A(inst_cellmath__61[10]));
INVXL cynw_cm_float_sin_I297 (.Y(N3658), .A(N3657));
INVX2 cynw_cm_float_sin_I298 (.Y(N3659), .A(inst_cellmath__61[6]));
INVXL cynw_cm_float_sin_I299 (.Y(N3660), .A(N3659));
INVXL cynw_cm_float_sin_I301 (.Y(N3662), .A(N3661));
XNOR2X1 cynw_cm_float_sin_I10044 (.Y(N3665), .A(N7631), .B(N741));
INVXL cynw_cm_float_sin_I305 (.Y(N3666), .A(N3665));
XNOR2X1 cynw_cm_float_sin_I10045 (.Y(inst_cellmath__115__W1[0]), .A(N7631), .B(N749));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1361 (.Y(N8384), .A(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1362 (.Y(N8665), .A(inst_cellmath__61[21]), .B(inst_cellmath__61[20]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10046 (.Y(N8493), .A(N8384), .B(N8665));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1366 (.Y(N8108), .A(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1367 (.Y(N8274), .A(inst_cellmath__61[18]), .B(inst_cellmath__61[17]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10047 (.Y(N8202), .A(N8108), .B(N8274));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1371 (.Y(N8253), .A(N8202), .B(N8493));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1372 (.Y(N7906), .A(inst_cellmath__61[17]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1373 (.Y(N8130), .A(inst_cellmath__61[18]), .B(N7906));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1374 (.Y(N8162), .A(N8130), .B(N8108));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1375 (.Y(N8657), .A(N8162));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1377 (.Y(N8617), .A(N8493), .B(N8657));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1378 (.Y(N7746), .A(inst_cellmath__61[18]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1379 (.Y(N8000), .A(N7746), .B(inst_cellmath__61[17]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10049 (.Y(N8749), .A(N8108), .B(N8000));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1383 (.Y(N8481), .A(N8493), .B(N8749));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1384 (.Y(N8720), .A(N7746), .B(N7906));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I9982 (.Y(N22608), .A(N8108), .B(N8720));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1389 (.Y(N8095), .A(N8493), .B(N22608));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1390 (.Y(N7988), .A(N8274), .B(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1391 (.Y(N8462), .A(N8493), .B(N7988));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1392 (.Y(N8707), .A(N8130), .B(inst_cellmath__61[19]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1393 (.Y(N8087), .A(N8707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1395 (.Y(N7959), .A(N8493), .B(N8087));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10051 (.Y(N7689), .A(inst_cellmath__61[19]), .B(N8000));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1399 (.Y(N8441), .A(N8493), .B(N7689));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10200 (.Y(N8425), .A(inst_cellmath__61[19]), .B(N8720));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1404 (.Y(N7813), .A(N8493), .B(N8425));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1405 (.Y(N8060), .A(inst_cellmath__61[20]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1406 (.Y(N8290), .A(inst_cellmath__61[21]), .B(N8060));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10053 (.Y(N8534), .A(N8384), .B(N8290));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1410 (.Y(N8776), .A(N8202), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1411 (.Y(N7921), .A(N8657), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1412 (.Y(N8150), .A(N8749), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1413 (.Y(N8397), .A(N22608), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1414 (.Y(N8637), .A(N7988), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1415 (.Y(N8660), .A(N8534), .B(N8087));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1416 (.Y(N8017), .A(N7689), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1417 (.Y(N8256), .A(N8425), .B(N8534));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1418 (.Y(N8500), .A(inst_cellmath__61[21]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1419 (.Y(N8739), .A(N8500), .B(inst_cellmath__61[20]));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10315 (.Y(N8489), .A(N8384), .B(N8739));
OR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1423 (.Y(N8728), .A(N8489), .B(N8202));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1424 (.Y(N7870), .A(N8728));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1425 (.Y(N8349), .A(N8489), .B(N8657));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1426 (.Y(N8598), .A(N8489), .B(N8749));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1427 (.Y(N7719), .A(N8489), .B(N22608));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1428 (.Y(N7900), .A(N8489), .B(N7988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1429 (.Y(N8211), .A(N8489), .B(N8087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1430 (.Y(N8364), .A(N8489), .B(N7689));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1431 (.Y(N8688), .A(N8489), .B(N8425));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1432 (.Y(N7832), .A(N8500), .B(N8060));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10055 (.Y(N7822), .A(N8384), .B(N7832));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1436 (.Y(N8305), .A(N8202), .B(N7822));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1437 (.Y(N8228), .A(N7822), .B(N8657));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1438 (.Y(N7676), .A(N8749), .B(N7822));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1439 (.Y(N7939), .A(N22608), .B(N7822));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1440 (.Y(N8170), .A(N7988), .B(N7822));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1441 (.Y(N8414), .A(N7822), .B(N8087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1442 (.Y(N8663), .A(N7822), .B(N7689));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1443 (.Y(N7787), .A(N7822), .B(N8425));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10056 (.Y(N7929), .A(inst_cellmath__61[22]), .B(N8665));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1447 (.Y(N8090), .A(N8202), .B(N7929));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1448 (.Y(N8521), .A(N7929), .B(N8657));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1449 (.Y(N8756), .A(N7929), .B(N8749));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1450 (.Y(N7901), .A(N7929), .B(N22608));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1451 (.Y(N8128), .A(N7988), .B(N7929));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1452 (.Y(N8366), .A(N7929), .B(N8087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1453 (.Y(N8613), .A(N7929), .B(N7689));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1454 (.Y(N7739), .A(N7929), .B(N8425));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1455 (.Y(N8574), .A(inst_cellmath__61[22]), .B(N8290));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1456 (.Y(N8231), .A(N8202), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1457 (.Y(N8475), .A(N8657), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1458 (.Y(N8715), .A(N8749), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1459 (.Y(N7856), .A(N22608), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1460 (.Y(N8091), .A(N7988), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1461 (.Y(N8327), .A(N8087), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1462 (.Y(N8577), .A(N7689), .B(N8574));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1463 (.Y(N7699), .A(N8425), .B(N8574));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10202 (.Y(N8745), .A(inst_cellmath__61[22]), .B(N8739));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1467 (.Y(N8431), .A(N8202), .B(N8745));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1468 (.Y(N8433), .A(N8745), .B(N8657));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1469 (.Y(N8674), .A(N8749), .B(N8745));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1470 (.Y(N7807), .A(N8745), .B(N22608));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1471 (.Y(N7804), .A(N7988), .B(N8745));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1472 (.Y(N8286), .A(N8745), .B(N8087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1473 (.Y(N8539), .A(N7689), .B(N8745));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1474 (.Y(N8285), .A(N8425), .B(N8745));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10058 (.Y(N8080), .A(inst_cellmath__61[22]), .B(N7832));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1478 (.Y(N8148), .A(N8202), .B(N8080));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1479 (.Y(N8389), .A(N8080), .B(N8657));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1480 (.Y(N8632), .A(N8749), .B(N8080));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1481 (.Y(N7759), .A(N8080), .B(N22608));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1482 (.Y(N8145), .A(N7988), .B(N8080));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1483 (.Y(N8629), .A(N8080), .B(N8087));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1484 (.Y(N8497), .A(N7689), .B(N8080));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1485 (.Y(N8736), .A(N8425), .B(N8080));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1486 (.Y(N8177), .A(N8253));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1487 (.Y(N8526), .A(N8617));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10059 (.Y(N8373), .A(N8253), .B(N8617));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1491 (.Y(N8236), .A(N8481));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1492 (.Y(N8097), .A(N8095));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10060 (.Y(N7704), .A(N8481), .B(N8095));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1497 (.Y(N7876), .A(N7959), .B(N8462));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1498 (.Y(N8777), .A(N7959));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1499 (.Y(N8640), .A(N8462));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1500 (.Y(N8502), .A(N8441));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1501 (.Y(N8350), .A(N7813));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10061 (.Y(N7977), .A(N8441), .B(N7813));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10062 (.Y(N8307), .A(N8776), .B(N7921));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1508 (.Y(N8171), .A(N8776));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1509 (.Y(N8043), .A(N7921));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1510 (.Y(N8201), .A(N8397), .B(N8150));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1511 (.Y(N8615), .A(N8397));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1513 (.Y(N8478), .A(N8150));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1514 (.Y(N8329), .A(N8660));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1515 (.Y(N8435), .A(N8637));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1516 (.Y(N8675), .A(N8637), .B(N8660));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1517 (.Y(N8057), .A(N8675));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1519 (.Y(N8392), .A(N8017));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10063 (.Y(N8250), .A(N8017), .B(N8256));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1524 (.Y(N8110), .A(N8256));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1525 (.Y(N8554), .A(N8349), .B(N7870));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1526 (.Y(N7937), .A(N8349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1527 (.Y(N7780), .A(N7719));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1528 (.Y(N8518), .A(N7719), .B(N8598));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1529 (.Y(N8363), .A(N8598));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1530 (.Y(N8408), .A(N7900), .B(N8211));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1531 (.Y(N8712), .A(N7900));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1532 (.Y(N7692), .A(N8211));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1533 (.Y(N7803), .A(N8688));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1534 (.Y(N8769), .A(N8364));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10064 (.Y(N8383), .A(N8688), .B(N8364));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1538 (.Y(N8245), .A(N8228));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1539 (.Y(N8106), .A(N8305));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10065 (.Y(N8456), .A(N8305), .B(N8228));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1543 (.Y(N7933), .A(N7939));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1544 (.Y(N7775), .A(N7939), .B(N7676));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1545 (.Y(N8514), .A(N7676));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1546 (.Y(N7985), .A(N8414), .B(N8170));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1547 (.Y(N7848), .A(N8414));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1548 (.Y(N7687), .A(N8170));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1549 (.Y(N8606), .A(N7787), .B(N8663));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1551 (.Y(N8378), .A(N7787));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1552 (.Y(N7987), .A(N8521), .B(N8090));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1553 (.Y(N8488), .A(N8090));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1555 (.Y(N8338), .A(N7901));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1556 (.Y(N8195), .A(N8756));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1557 (.Y(N8067), .A(N7901), .B(N8756));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1558 (.Y(N8781), .A(N8128));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10066 (.Y(N8648), .A(N8128), .B(N8366));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1561 (.Y(N8506), .A(N8366));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1562 (.Y(N8115), .A(N8613), .B(N7739));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1565 (.Y(N8312), .A(N8613));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1566 (.Y(N8176), .A(N8231));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1567 (.Y(N8666), .A(N8475), .B(N8231));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1568 (.Y(N8524), .A(N8475));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1569 (.Y(N8371), .A(N7856));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1570 (.Y(N8721), .A(N8715));
OR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1572 (.Y(N7864), .A(N7856), .B(N8715));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1573 (.Y(N8331), .A(N7864));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1575 (.Y(N8442), .A(N8091));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1576 (.Y(N8291), .A(N8327));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10067 (.Y(N8638), .A(N8091), .B(N8327));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1580 (.Y(N8501), .A(N7699));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1581 (.Y(N8050), .A(N8577), .B(N7699));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1582 (.Y(N7720), .A(N8577));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1583 (.Y(N7833), .A(N8433));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10068 (.Y(N7677), .A(N8433), .B(N8431));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1588 (.Y(N8415), .A(N8431));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1589 (.Y(N8041), .A(N8674), .B(N7807));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1590 (.Y(N7902), .A(N7807));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1591 (.Y(N7740), .A(N8674));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10069 (.Y(N8716), .A(N7804), .B(N8286));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1595 (.Y(N8578), .A(N7804));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1596 (.Y(N7700), .A(N8286));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1597 (.Y(N7754), .A(N8539), .B(N8285));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1598 (.Y(N8774), .A(N8285));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1599 (.Y(N8633), .A(N8539));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1600 (.Y(N8737), .A(N8148));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10070 (.Y(N8593), .A(N8148), .B(N8389));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1604 (.Y(N8458), .A(N8389));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1606 (.Y(N8683), .A(N7759), .B(N8632));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1607 (.Y(N7826), .A(N8683));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1608 (.Y(N8164), .A(N8632));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1609 (.Y(N8037), .A(N7759));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1610 (.Y(N7897), .A(N8629));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1612 (.Y(N8223), .A(N8629), .B(N8145));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1613 (.Y(N8089), .A(N8145));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1614 (.Y(N7949), .A(N8736));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10203 (.Y(N7800), .A(N8736), .B(N8497));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1618 (.Y(N8768), .A(N8497));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1619 (.Y(N8427), .A(N8177), .B(N8728));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1620 (.Y(N7801), .A(N8781), .B(N8442));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1621 (.Y(N8052), .A(N8176), .B(N7897));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1622 (.Y(N8283), .AN(N7856), .B(N7803));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1623 (.Y(N8535), .A(N8338), .B(N8236));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1624 (.Y(N7967), .A(N8245), .B(N7833));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1626 (.Y(N8627), .A(N8201), .B(N7754));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1627 (.Y(N8450), .A(N7987), .B(N7876));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1628 (.Y(N7821), .AN(N8683), .B(N8041));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1630 (.Y(N8732), .A(N8535), .B(N8627));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1631 (.Y(N7874), .A(N7801), .B(N8450));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1632 (.Y(N7960), .A(N8307), .B(N8606));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1633 (.Y(N8342), .A(N7821), .B(N7960));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28186 (.Y(N8590), .A(N8427), .B(N7939), .C(N8052), .D(N8283));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1635 (.Y(N7711), .A(N8732), .B(N7874));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1636 (.Y(N7744), .A(N8392), .B(N8408), .C(N8342));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1637 (.Y(N8454), .A(N7967), .B(N7744));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1638 (.Y(N8198), .A(N8590), .B(N7711));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1640 (.Y(N7932), .A(N8488), .B(N8728));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1641 (.Y(N8158), .A(N8712), .B(N8737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1642 (.Y(N8405), .A(N8106), .B(N8171));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1643 (.Y(N8651), .A(N7897), .B(N7803));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1644 (.Y(N7772), .A(N8502), .B(N8291));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1645 (.Y(N8028), .A(N8371), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1646 (.Y(N8265), .A(N7985), .B(N7933));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1647 (.Y(N8298), .A(N7780), .B(N8716));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1648 (.Y(N8747), .A(N8115), .B(N8666));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1649 (.Y(N7892), .A(N8250), .B(N7677));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1650 (.Y(N8119), .A(N8606));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1651 (.Y(N8105), .A(N7826));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1652 (.Y(N7983), .A(N7772), .B(N8405));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1653 (.Y(N8219), .A(N8747), .B(N7892));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1654 (.Y(N8470), .A(N8298), .B(N8651));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1655 (.Y(N8703), .A(N8265), .B(N8028));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1656 (.Y(N8084), .A(N8470), .B(N8703));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1657 (.Y(N7684), .AN(N7826), .B(N8119), .C(N7932), .D(N8158));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1658 (.Y(N8546), .A(N7983), .B(N8219));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1659 (.Y(N8568), .A(N8084), .B(N8546));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1661 (.Y(N8764), .A(N8615), .B(N8774));
INVXL cynw_cm_float_sin_I28137 (.Y(N8531), .A(N8663));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1662 (.Y(N8134), .A(N8531), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1663 (.Y(N8375), .A(N8350), .B(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1664 (.Y(N8620), .A(N8408), .B(N7985));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1665 (.Y(N7748), .A(N8638), .B(N8593));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1666 (.Y(N8004), .A(N8554), .B(N8307));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1667 (.Y(N8239), .A(N8648), .B(N8666));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1668 (.Y(N8485), .A(N8456), .B(N7775));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1669 (.Y(N8785), .A(N7826), .B(N8518));
INVX1 cynw_cm_float_sin_I28138 (.Y(N8215), .A(N7739));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1670 (.Y(N7868), .AN(N8764), .B(N8215), .C(N8721));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1671 (.Y(N8099), .A(N7748), .B(N7901));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1672 (.Y(N8336), .A(N8375), .B(N8485));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1673 (.Y(N8585), .A(N8620), .B(N8004));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1674 (.Y(N7706), .A(N8239), .B(N8134));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1675 (.Y(N8064), .A(N8785), .B(N7868));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1676 (.Y(N8446), .A(N8099), .B(N8336));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1677 (.Y(N8679), .A(N8585), .B(N7706));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1678 (.Y(N7817), .A(N8446), .B(N8679));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1680 (.Y(N7767), .AN(N8211), .B(N7897));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1681 (.Y(N8023), .A(N7803), .B(N7848));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1682 (.Y(N7989), .A(N8291), .B(N8371));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1683 (.Y(N8504), .A(N7937), .B(N8774));
INVX1 cynw_cm_float_sin_I27997 (.Y(N8727), .A(N8521));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1684 (.Y(N8742), .A(N8777), .B(N8727));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1685 (.Y(N8765), .A(N8215), .B(N8501));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1686 (.Y(N8126), .A(N8392), .B(N7949));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1687 (.Y(N8197), .A(N7775));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1688 (.Y(N8213), .A(N8197), .B(N8148));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1689 (.Y(N8580), .A(N8201), .B(N8506), .C(N8716));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1690 (.Y(N7838), .A(N8756), .B(N8580));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1691 (.Y(N8075), .A(N8504), .B(N8765));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1692 (.Y(N8310), .A(N7967), .B(N8126));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1693 (.Y(N8561), .A(N7989), .B(N7767));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1694 (.Y(N7679), .A(N8023));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1695 (.Y(N7942), .A(N7679), .B(N7838));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1696 (.Y(N8174), .A(N8075), .B(N8213));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1697 (.Y(N8418), .A(N8310), .B(N8561));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1698 (.Y(N7790), .A(N8105), .B(N8742), .C(N8174));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1699 (.Y(N8045), .A(N8418), .B(N7942));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1701 (.Y(N7863), .A(N8640), .B(N8171));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1702 (.Y(N7957), .A(N8638), .B(N8164));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1703 (.Y(N7816), .A(N7977), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1704 (.Y(N8022), .A(N7687), .B(N8176));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1705 (.Y(N7811), .A(N7863), .B(N8022));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1706 (.Y(N8541), .A(N8633), .B(N7833), .C(N7811));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1707 (.Y(N8636), .AN(N8371), .BN(N7692), .C(N7957), .D(N7816));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1708 (.Y(N8394), .AN(N8329), .B(N7676), .C(N8541), .D(N8119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1710 (.Y(N8596), .A(N8578), .B(N8435));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1711 (.Y(N8157), .AN(N8539), .B(N8338));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1712 (.Y(N8209), .A(N8458), .B(N8777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1713 (.Y(N8687), .A(N8715), .B(N8596));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1714 (.Y(N7831), .A(N8245), .B(N8392));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1715 (.Y(N8649), .A(N7902), .B(N7985));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1716 (.Y(N8559), .A(N8115), .B(N7800));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1717 (.Y(N7931), .A(N8518));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1718 (.Y(N7938), .A(N7931), .B(N8209));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1719 (.Y(N8169), .A(N8559), .B(N8649));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1720 (.Y(N7784), .A(N8687), .B(N8169));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1721 (.Y(N7978), .A(N8164), .B(N8554), .C(N7938));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1722 (.Y(N8754), .A(N8157), .B(N7978));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1723 (.Y(N8520), .AN(N8291), .BN(N8171), .C(N7784), .D(N7831));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1725 (.Y(N8229), .A(N8177), .B(N8578));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1726 (.Y(N8714), .A(N8640), .B(N8737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1727 (.Y(N8576), .A(N8291), .B(N8478));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1728 (.Y(N7696), .A(N8721), .B(N8727));
NAND2BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1729 (.Y(N7952), .AN(N8675), .B(N8195));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1730 (.Y(N8376), .A(N8097), .B(N8524));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1731 (.Y(N8432), .A(N8501), .B(N7833));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1732 (.Y(N7806), .A(N7933), .B(N8037));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1733 (.Y(N8056), .A(N8554), .B(N7977));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1734 (.Y(N8538), .A(N8714), .B(N7952));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1735 (.Y(N8309), .A(N8378), .B(N7949));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1736 (.Y(N8772), .A(N8056), .B(N8309));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I1737 (.Y(N8147), .AN(N8613), .BN(N8229), .C(N8518), .D(N8250));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1738 (.Y(N7789), .A(N7687), .B(N7692));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1739 (.Y(N8386), .A(N7696), .B(N7789));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1740 (.Y(N8630), .A(N7806), .B(N8376));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1741 (.Y(N8249), .A(N8386), .B(N8630));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1742 (.Y(N8370), .A(N8538), .B(N8772));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1743 (.Y(N8495), .A(N8147), .B(N8370));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1744 (.Y(N7878), .A(N8432), .B(N8576), .C(N8249));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1747 (.Y(N7962), .A(N8777), .B(N8057));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1748 (.Y(N7670), .A(N7985), .B(N8164));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1749 (.Y(N8025), .A(N8067), .B(N8201));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1750 (.Y(N8163), .A(N8554), .B(N7987));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1751 (.Y(N7771), .A(N8307), .B(N8716));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1752 (.Y(N7891), .A(N8648), .B(N8115));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1753 (.Y(N7778), .A(N8050), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1754 (.Y(N8034), .A(N8606), .B(N7800));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1755 (.Y(N7862), .A(N8236), .B(N8110));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1757 (.Y(N7896), .A(N7778), .B(N7771));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1758 (.Y(N8123), .A(N8034), .B(N8163));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28233 (.Y(N8607), .A(N7676), .B(N8253), .C(N7862), .D(N7891));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1761 (.Y(N8708), .A(N7962), .B(N7670), .C(N8607));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1762 (.Y(N8439), .A(N7896), .B(N8123));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I10072 (.Y(N7851), .A(N7931), .B(N7989), .C(N8025), .D(N8439));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1765 (.Y(N8185), .A(N8176), .B(N8329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1766 (.Y(N8354), .A(N8526), .B(N8769));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1767 (.Y(N7798), .A(N8629), .B(N8354));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1768 (.Y(N8314), .A(N8727), .B(N8195));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1769 (.Y(N8566), .A(N8236), .B(N8506));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1770 (.Y(N8767), .A(N8043), .B(N8501));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1771 (.Y(N7716), .A(N7754), .B(N8716));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1772 (.Y(N8625), .A(N8115), .B(N8250));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1773 (.Y(N8242), .A(N7931), .B(N8185));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1774 (.Y(N8490), .A(N8714), .B(N7716));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1775 (.Y(N8729), .A(N8625), .B(N8767));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1776 (.Y(N7871), .A(N8314), .B(N8034));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1777 (.Y(N7709), .A(N7833), .B(N8408), .C(N7871));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1778 (.Y(N7968), .A(N8242), .B(N7798));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1779 (.Y(N8299), .AN(N8291), .BN(N8721), .C(N8566), .D(N7670));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1780 (.Y(N8069), .AN(N8490), .BN(N8729), .C(N7968), .D(N7709));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1782 (.Y(N8650), .A(N7720), .B(N8777));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1783 (.Y(N7770), .A(N8721), .B(N8057));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1784 (.Y(N8139), .A(N8195), .B(N8236));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1785 (.Y(N8263), .A(N8506), .B(N8043));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1786 (.Y(N8509), .A(N8373), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1787 (.Y(N8746), .A(N8215), .B(N8531));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1789 (.Y(N8355), .A(N8638), .B(N7933));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1790 (.Y(N7875), .A(N8201), .B(N8554));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1791 (.Y(N7918), .A(N8106), .B(N7848));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1792 (.Y(N8082), .A(N8509), .B(N7918));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I28236 (.Y(N7946), .A(N8110), .B(N8383), .C(N8524), .D(N8350));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1795 (.Y(N8700), .A(N7821), .B(N7875));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1796 (.Y(N7843), .A(N8263), .B(N8746));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1797 (.Y(N7975), .A(N8716), .B(N7677));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1798 (.Y(N8565), .A(N8355), .B(N7975));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1799 (.Y(N7683), .A(N8650), .B(N8139));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1800 (.Y(N8178), .A(N7946), .B(N7770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1801 (.Y(N8422), .A(N8700), .B(N7843));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1802 (.Y(N8276), .A(N8565), .B(N7683));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1803 (.Y(N8558), .A(N8488), .B(N8737), .C(N8082));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1804 (.Y(N8762), .A(N8422), .B(N8558));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1805 (.Y(N8527), .A(N8276), .B(N8178));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1807 (.Y(N8020), .A(N8091), .B(N8660));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1808 (.Y(N8334), .A(N8615), .B(N8458));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1809 (.Y(N8584), .A(N8727), .B(N8506));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1810 (.Y(N7705), .A(N8215), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1811 (.Y(N8267), .A(N7876), .B(N7780));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1812 (.Y(N8778), .A(N8649), .B(N8267));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1813 (.Y(N7925), .A(N8157));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1814 (.Y(N8152), .AN(N8334), .B(N8050), .C(N7925));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1815 (.Y(N8039), .A(N8524), .B(N8245));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1816 (.Y(N8401), .A(N7771), .B(N8039));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1817 (.Y(N8643), .A(N8584), .B(N7705));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1818 (.Y(N7764), .A(N7767), .B(N8126));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1819 (.Y(N8740), .A(N8643), .B(N7764));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1820 (.Y(N7994), .A(N8020), .B(N7933), .C(N8331));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1821 (.Y(N8351), .A(N8740), .B(N7994));
NAND4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1822 (.Y(N770), .AN(N8152), .B(N8401), .C(N8351), .D(N8778));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1823 (.Y(N8692), .A(N8171), .B(N8526));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1824 (.Y(N8560), .A(N8415), .B(N8291), .C(N8435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1825 (.Y(N7678), .A(N8478), .B(N8458));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1826 (.Y(N7940), .A(N8777), .B(N8236));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1827 (.Y(N8172), .A(N8215), .B(N8350));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1828 (.Y(N8044), .A(N8067), .B(N7754));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1829 (.Y(N7727), .A(N8716), .B(N8648));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1830 (.Y(N8217), .A(N8666), .B(N8050));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1831 (.Y(N8616), .A(N8250), .B(N7800));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1832 (.Y(N7903), .A(N8041), .B(N8518));
NOR3X1 inst_cellmath__195__80__2WWMM_2WWMM_I1833 (.Y(N8479), .A(N8044), .B(N8217), .C(N7727));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1834 (.Y(N7860), .AN(N8408), .B(N7864), .C(N7678), .D(N7940));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1835 (.Y(N8325), .A(N8245), .B(N8378));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1836 (.Y(N8093), .A(N8172), .B(N8325));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1837 (.Y(N8436), .A(N8692), .B(N7903), .C(N7806));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1838 (.Y(N7701), .A(N8364), .B(N8090), .C(N8616), .D(N8560));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1839 (.Y(N7805), .A(N8093), .B(N8479));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1840 (.Y(N8676), .A(N8436), .B(N7805));
NAND3X1 inst_cellmath__195__80__2WWMM_2WWMM_I1841 (.Y(N771), .A(N7701), .B(N7860), .C(N8676));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1842 (.Y(N8393), .A(N8640), .B(N8578));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1843 (.Y(N7761), .A(N7740), .B(N8312));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1844 (.Y(N8252), .A(N8371), .B(N8478));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1845 (.Y(N8348), .A(N7687), .B(N8526), .C(N7933));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1846 (.Y(N8698), .A(N8593), .B(N8554));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1847 (.Y(N7718), .A(N7987), .B(N7780));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1848 (.Y(N8079), .A(N8606), .B(N8456));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1849 (.Y(N8207), .A(N7800));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1850 (.Y(N7829), .A(N7761), .B(N8393), .C(N8079));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1851 (.Y(N8385), .A(N8223), .B(N8392));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1852 (.Y(N8303), .A(N8376), .B(N8385));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1853 (.Y(N8038), .A(N8348), .B(N8157), .C(N8698));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1854 (.Y(N8659), .A(N7829), .B(N8303));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1855 (.Y(N7781), .A(N8207), .B(N8252), .C(N7718), .D(N8659));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1857 (.Y(N7737), .A(N8435), .B(N8442));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1858 (.Y(N7993), .A(N8176), .B(N8526));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1859 (.Y(N7854), .A(N8688), .B(N7737));
NAND3X1 inst_cellmath__195__80__2WWMM_2WWMM_I1860 (.Y(N8322), .A(N8415), .B(N8578), .C(N8371));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1861 (.Y(N8573), .A(N7720), .B(N8774));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1862 (.Y(N7694), .A(N8727), .B(N8236));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1863 (.Y(N8188), .A(N8378), .B(N7902));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1864 (.Y(N8429), .A(N7985));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1865 (.Y(N8054), .A(N8363), .B(N7933), .C(N8110));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1866 (.Y(N8564), .A(N8307), .B(N8648));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1867 (.Y(N7913), .A(N8456));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1868 (.Y(N8144), .A(N7913), .B(N8188));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1869 (.Y(N8247), .A(N7993), .B(N8564));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1870 (.Y(N7877), .A(N8115), .B(N7977));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1872 (.Y(N8591), .A(N8640), .B(N7692), .C(N8144));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I28258 (.Y(N8344), .AN(N7854), .B(N7877), .C(N8054), .D(N8698));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1874 (.Y(N8107), .A(N8322), .B(N8573), .C(N8429));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1876 (.Y(N8287), .A(N8247), .B(N7694), .C(N8107));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1877 (.Y(N7972), .A(N8591), .B(N8287));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1879 (.Y(N7669), .A(N8435), .B(N8106));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1880 (.Y(N7934), .A(N7687), .B(N8769));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1881 (.Y(N7986), .AN(N8674), .B(N8177), .C(N8089));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1882 (.Y(N7777), .A(N8458), .B(N8774));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1883 (.Y(N8032), .A(N8768), .B(N8721));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1884 (.Y(N7849), .A(N8164), .B(N8067));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1885 (.Y(N8284), .A(N7876), .B(N8716));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1886 (.Y(N8605), .A(N8119), .B(N8217));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1887 (.Y(N7733), .A(N7669), .B(N7934));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1888 (.Y(N8457), .A(N8043), .B(N8350));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1889 (.Y(N8472), .A(N7777), .B(N8457));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1890 (.Y(N8705), .A(N8284), .B(N8032));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1891 (.Y(N8571), .A(N7692), .B(N8615), .C(N8472));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1892 (.Y(N7688), .A(N8605), .B(N8705));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1893 (.Y(N8182), .A(N7986), .B(N7891), .C(N7688));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1894 (.Y(N7936), .A(N7849), .B(N7733));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1895 (.Y(N8424), .A(N8571), .B(N7936));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1897 (.Y(N8717), .A(N7848), .B(N8502));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1898 (.Y(N7753), .A(N8478), .B(N8633));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1899 (.Y(N8083), .A(N8458), .B(N7937));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1900 (.Y(N8317), .A(N8083));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1901 (.Y(N7820), .A(N8110), .B(N8245));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1902 (.Y(N7947), .A(N8606), .B(N7677));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1903 (.Y(N8339), .A(N7800), .B(N7826));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1904 (.Y(N8449), .A(N8364), .B(N8717));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1905 (.Y(N7964), .A(N7947), .B(N8267));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1906 (.Y(N8549), .A(N8716), .B(N8050), .C(N8449));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1907 (.Y(N7928), .AN(N8057), .BN(N8043), .C(N8339), .D(N7820));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1908 (.Y(N8297), .AN(N7753), .B(N8083), .C(N7964));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1909 (.Y(N8783), .A(N8549), .B(N8297));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1911 (.Y(N7769), .AN(N8128), .B(N8488));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1912 (.Y(N8116), .A(N7848), .B(N8312));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1913 (.Y(N8216), .A(N7833), .B(N8378));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1914 (.Y(N8467), .A(N8392), .B(N7902));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1915 (.Y(N8313), .A(N8037), .B(N8593));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1916 (.Y(N8563), .A(N7977), .B(N7876));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1917 (.Y(N8759), .A(N8405), .B(N7952));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1918 (.Y(N8419), .AN(N8633), .BN(N7937), .C(N8313), .D(N8563));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1919 (.Y(N7791), .AN(N8578), .BN(N8442), .C(N8216), .D(N8116));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1920 (.Y(N8046), .A(N8032), .B(N8467));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1921 (.Y(N8525), .A(N8231), .B(N7769), .C(N7767));
NAND4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1922 (.Y(N8618), .A(N7933), .B(N8363), .C(N8501), .D(N8759));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1923 (.Y(N8131), .A(N8046), .B(N8419));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1924 (.Y(N7747), .A(N8618), .B(N8131));
NAND3X1 inst_cellmath__195__80__2WWMM_2WWMM_I1925 (.Y(N776), .A(N7791), .B(N8525), .C(N7747));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1927 (.Y(N8443), .A(N7687), .B(N7897));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1928 (.Y(N7814), .A(N8373), .B(N8057));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1929 (.Y(N8061), .A(N8501), .B(N8378));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1930 (.Y(N8292), .A(N7902), .B(N8383));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1934 (.Y(N8400), .A(N7987), .B(N8648));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I28263 (.Y(N8257), .AN(N8638), .B(N7870), .C(N8400), .D(N8431));
NAND2BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1932 (.Y(N7923), .AN(N7814), .B(N7933));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1933 (.Y(N8111), .A(N8164), .B(N7754));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1935 (.Y(N8639), .A(N7704), .B(N8666));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I1937 (.Y(N7721), .AN(N8061), .BN(N8292), .C(N7692), .D(N8458));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1938 (.Y(N7834), .AN(N8250), .B(N8443), .C(N7923), .D(N8639));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1939 (.Y(N8517), .A(N8111), .B(N8257));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1940 (.Y(N8690), .A(N7721), .B(N8517));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1942 (.Y(N8757), .A(N8145), .B(N7900));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1943 (.Y(N7951), .A(N7720), .B(N8458));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1944 (.Y(N7741), .A(N8638), .B(N8531), .C(N8057), .D(N8757));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1945 (.Y(N7997), .A(N7933), .B(N8554));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1946 (.Y(N7954), .A(N7727), .B(N7951), .C(N7741));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1947 (.Y(N8191), .A(N7997), .B(N8625), .C(N8785), .D(N8649));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1949 (.Y(N8390), .A(N8737), .B(N8514));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1950 (.Y(N8634), .A(N8057), .B(N8408));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1951 (.Y(N8118), .A(N8666), .B(N8250));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1952 (.Y(N7881), .A(N8456), .B(N8518));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1953 (.Y(N8685), .AN(N7891), .B(N8331), .C(N8554));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1954 (.Y(N8459), .A(N8390), .B(N8292), .C(N8634));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1955 (.Y(N7827), .A(N7881), .B(N7716), .C(N8118), .D(N8685));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10074 (.Y(N7792), .A(N8638), .B(N8331));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1958 (.Y(N8752), .A(N8201), .B(N7876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1959 (.Y(N8125), .A(N8115), .B(N7704));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1960 (.Y(N8609), .A(N7977), .B(N7677));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1961 (.Y(N8225), .A(N8217), .B(N8564));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1962 (.Y(N8710), .AN(N7740), .BN(N8373), .C(N8125), .D(N8609));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I1963 (.Y(N780), .AN(N8752), .BN(N7792), .C(N8225), .D(N8710));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1964 (.Y(N8536), .A(N7985), .B(N8067));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1965 (.Y(N8140), .A(N8307), .B(N7704));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10075 (.Y(N8047), .A(N7977), .B(N8250));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1969 (.Y(N7755), .A(N7775), .B(N8518));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1970 (.Y(N8244), .A(N8140), .B(N8047));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1971 (.Y(N8492), .A(N8079), .B(N7755));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1972 (.Y(N7969), .AN(N8383), .BN(N8408), .C(N7875), .D(N8450));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1973 (.Y(N8341), .A(N8244), .B(N8492));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1974 (.Y(N7712), .A(N8536), .B(N7814), .C(N8341));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I9890 (.Y(N22540), .A(N7712), .B(N7969));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1976 (.Y(N8702), .A(N8502), .B(N8721));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1977 (.Y(N7846), .A(N8195), .B(N8043));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1978 (.Y(N7685), .A(N8383), .B(N7985));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1979 (.Y(N8278), .A(N8041));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1980 (.Y(N8529), .A(N8278), .B(N7846));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1981 (.Y(N8136), .A(N8716), .B(N7800), .C(N8392), .D(N8378));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1982 (.Y(N7749), .A(N8111), .B(N8529));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1983 (.Y(N8473), .A(N8781), .B(N7692), .C(N8728));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1984 (.Y(N8183), .A(N8638), .B(N8435), .C(N8176));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1985 (.Y(N8724), .A(N8702), .B(N7967), .C(N8765), .D(N8183));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1986 (.Y(N8335), .AN(N8724), .B(N8473), .C(N8136));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1988 (.Y(N8294), .A(N8415), .B(N8712));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1989 (.Y(N8528), .A(N8737), .B(N8442));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1990 (.Y(N7926), .A(N8312), .B(N7720));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1991 (.Y(N8403), .A(N8285), .B(N8294));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1992 (.Y(N8644), .A(N8727), .B(N8057));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1993 (.Y(N8696), .A(N7700), .B(N8506));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1994 (.Y(N8743), .A(N7704), .B(N8456));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I1995 (.Y(N7979), .AN(N8743), .B(N7949), .C(N8403), .D(N8331));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I1996 (.Y(N8562), .AN(N8696), .BN(N8692), .C(N8392), .D(N8531));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1997 (.Y(N8076), .A(N7926), .B(N8528), .C(N7931), .D(N8644));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1998 (.Y(N8533), .A(N8164), .B(N8201));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2001 (.Y(N8233), .A(N8524), .B(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2002 (.Y(N8480), .A(N7902), .B(N8638));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2003 (.Y(N8008), .A(N8712), .B(N8578));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2004 (.Y(N8582), .A(N8023), .B(N8008));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2005 (.Y(N7958), .A(N8106), .B(N7677), .C(N8514), .D(N8582));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2006 (.Y(N8440), .AN(N8727), .BN(N8215), .C(N8462), .D(N8150));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2007 (.Y(N7810), .AN(N8307), .BN(N8250), .C(N8233), .D(N8480));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2010 (.Y(N8254), .A(N8578), .B(N7687));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2011 (.Y(N7885), .A(N8777), .B(N8768));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2012 (.Y(N7908), .A(N7775), .B(N7826));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2013 (.Y(N7830), .AN(N8254), .B(N8350), .C(N8378));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2014 (.Y(N7783), .AN(N8554), .BN(N8456), .C(N7908), .D(N8025));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2016 (.Y(N8661), .AN(N8363), .BN(N8097), .C(N8467), .D(N7885));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2017 (.Y(N8519), .AN(N7830), .B(N7803), .C(N8661), .D(N8312));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2019 (.Y(N8230), .A(N8089), .B(N8106));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2020 (.Y(N8773), .A(N8769), .B(N7848));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2021 (.Y(N8575), .A(N8506), .B(N8215));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2022 (.Y(N8146), .A(N8524), .B(N8110));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2023 (.Y(N8374), .A(N7800), .B(N8041));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2024 (.Y(N7915), .A(N8349), .B(N7900), .C(N8773));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2025 (.Y(N8388), .A(N8197), .B(N8146), .C(N8374));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I2026 (.Y(N7757), .AN(N8230), .BN(N8140), .C(N8593), .D(N8716));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2027 (.Y(N8735), .A(N8575), .B(N8216));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2028 (.Y(N8494), .A(N7915), .B(N8388));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2030 (.Y(N7715), .AN(N8777), .BN(N8721), .C(N8644), .D(N7757));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2033 (.Y(N8555), .A(N8488), .B(N8712));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2034 (.Y(N8035), .A(N8223), .B(N8245));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2035 (.Y(N8272), .A(N7833), .B(N8392));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2036 (.Y(N7690), .A(N7803), .B(N7933), .C(N8435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2037 (.Y(N7734), .A(N8067), .B(N7780));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2038 (.Y(N8361), .A(N8666), .B(N8606));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2039 (.Y(N7991), .A(N8577), .B(N7734), .C(N8555));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2040 (.Y(N8709), .AN(N8777), .BN(N8097), .C(N8564), .D(N8361));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2041 (.Y(N7852), .A(N7777), .B(N8272));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2042 (.Y(N8321), .A(N7772), .B(N8035), .C(N7991));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2043 (.Y(inst_cellmath__197[5]), .A(N7690), .B(N7852), .C(N8709), .D(N8321));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2044 (.Y(N8381), .A(N8781), .B(N8435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2045 (.Y(N8626), .A(N7692), .B(N8312));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2046 (.Y(N8731), .A(N8245), .B(N7985));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2047 (.Y(N8452), .A(N8638), .B(N8716));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2048 (.Y(N7930), .AN(N8050), .BN(N8606), .C(N8381), .D(N8452));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2049 (.Y(N8068), .A(N7931), .B(N7821), .C(N8731));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2050 (.Y(N8552), .AN(N8615), .BN(N8633), .C(N8742), .D(N8146));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2051 (.Y(N8787), .A(N8626), .B(N8317));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2052 (.Y(inst_cellmath__197[6]), .A(N8552), .B(N8068), .C(N7930), .D(N8787));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2053 (.Y(N7728), .A(N8171), .B(N8769));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2054 (.Y(N7844), .A(N7833), .B(N7949));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2055 (.Y(N8081), .A(N8408), .B(N8037));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2056 (.Y(N8316), .A(N8554), .B(N7876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2057 (.Y(N8567), .A(N7987), .B(N8050));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2059 (.Y(N8589), .A(N7700), .B(N8363));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2060 (.Y(N8421), .A(N8567), .B(N8589));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2065 (.Y(N8262), .A(N8089), .B(N8435), .C(N8421));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I28266 (.Y(N8237), .AN(N7925), .B(N7913), .C(N8262), .D(N8081));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2062 (.Y(N8133), .AN(N8215), .BN(N8524), .C(N7728), .D(N8047));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2063 (.Y(N8550), .A(N7740), .B(N8371), .C(N8316));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2068 (.Y(N8002), .A(N8721), .B(N8195));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2069 (.Y(N7766), .A(N8501), .B(N8350));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2070 (.Y(N7924), .A(N7933), .B(N7876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2071 (.Y(N8154), .A(N8648), .B(N7704));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2072 (.Y(N8642), .A(N8616), .B(N8154));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2073 (.Y(N8019), .AN(N8509), .B(N8578), .C(N7766), .D(N8488));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2074 (.Y(N8503), .A(N7687), .B(N8633), .C(N8642));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2075 (.Y(N7723), .A(N8480), .B(N7967));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2076 (.Y(N8113), .A(N8317), .B(N8019));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2077 (.Y(N8602), .AN(N8378), .BN(N8408), .C(N8002), .D(N8503));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2078 (.Y(inst_cellmath__197[8]), .A(N7924), .B(N7723), .C(N8602), .D(N8113));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2079 (.Y(N8445), .A(N8176), .B(N8514));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2080 (.Y(N8416), .A(N8329), .B(N8526));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I2081 (.Y(N7788), .AN(N7769), .B(N7692));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2082 (.Y(N8094), .A(N8097), .B(N8223));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2084 (.Y(N7955), .A(N8392), .B(N8383));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2085 (.Y(N8232), .A(N8041), .B(N8456), .C(N8067), .D(N7677));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2086 (.Y(N7982), .A(N8363), .B(N8768), .C(N8445));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2087 (.Y(N8437), .A(N8094), .B(N7982));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2088 (.Y(N8581), .A(N8371), .B(N7720), .C(N8777), .D(N7937));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2089 (.Y(N8315), .A(N7955), .B(N8581));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2090 (.Y(N8058), .A(N8717), .B(N8232), .C(N7788), .D(N8315));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2092 (.Y(N8251), .A(N7803), .B(N8502));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2093 (.Y(N7883), .A(N8245), .B(N8408));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2094 (.Y(N8304), .A(N8716), .B(N7704));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2095 (.Y(N8206), .A(N8050), .B(N7677), .C(N7775), .D(N8250));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2096 (.Y(N8461), .A(N8528), .B(N7718));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2097 (.Y(N8167), .AN(N8171), .BN(N7897), .C(N8251), .D(N7883));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2098 (.Y(N8275), .A(N8435), .B(N8728), .C(N8206));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2100 (.Y(N7782), .AN(N8304), .BN(N8461), .C(N7753), .D(N8575));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2102 (.Y(N8611), .A(N8728), .B(N8712));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2103 (.Y(N8227), .A(N8329), .B(N7740));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2104 (.Y(N8713), .A(N8478), .B(N8774));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2105 (.Y(N8323), .A(N8598), .B(N8611));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2106 (.Y(N8430), .A(N8392), .B(N8331));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2107 (.Y(N8055), .A(N8361), .B(N8713));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2108 (.Y(N8537), .AN(N8089), .BN(N8737), .C(N7769), .D(N8227));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2109 (.Y(N8771), .A(N7846), .B(N8251));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2111 (.Y(N8143), .A(N8771), .B(N8537));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2112 (.Y(N8003), .A(N7833), .B(N8106), .C(N8442));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2113 (.Y(N8246), .A(N8430), .B(N8003));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2115 (.Y(N7703), .A(N8164), .B(N7876), .C(N8246));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2116 (.Y(N8012), .A(N8765), .B(N7703));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2118 (.Y(N8200), .A(N8442), .B(N7848));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2119 (.Y(N8160), .AN(N8383), .BN(N8331), .C(N8286), .D(N8611));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I2120 (.Y(N8655), .AN(N8200), .B(N7933));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2121 (.Y(N8269), .A(N7677), .B(N7826));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2122 (.Y(N8062), .A(N8307), .B(N8666));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2123 (.Y(N7894), .A(N8269), .B(N8062));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2124 (.Y(N7732), .A(N8188), .B(N8172));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2125 (.Y(N8706), .AN(N7732), .B(N7734), .C(N7820), .D(N8713));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2127 (.Y(N7797), .A(N7937), .B(N8721));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2128 (.Y(N8532), .A(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2129 (.Y(N8380), .A(N7985), .B(N8638));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2130 (.Y(N7752), .A(N7704), .B(N7977));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2131 (.Y(N8587), .A(N8456), .B(N7800));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2132 (.Y(N8641), .A(N7740), .B(N8478));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2133 (.Y(N7966), .A(N8380), .B(N8641));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2134 (.Y(N8102), .A(N7752), .B(N8090), .C(N8532), .D(N8785));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2135 (.Y(N7708), .AN(N8587), .B(N7876), .C(N7797), .D(N8307));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2136 (.Y(N8681), .AN(N8696), .B(N8501), .C(N7925), .D(N8373));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2137 (.Y(N8601), .A(N7833), .B(N8176), .C(N8712));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2138 (.Y(N8782), .A(N7708), .B(N8601));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2140 (.Y(N8260), .A(N8640), .B(N8177));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2141 (.Y(N7725), .A(N8502), .B(N8338));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2142 (.Y(N8697), .A(N8501), .B(N8110));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2143 (.Y(N7841), .A(N8331));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2144 (.Y(N8078), .AN(N8236), .B(N7841), .C(N8260), .D(N8431));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2145 (.Y(N8614), .A(N8201), .B(N8593));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2146 (.Y(N8483), .A(N7754), .B(N7987));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2147 (.Y(N8667), .A(N7719), .B(N8483));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2148 (.Y(N8372), .AN(N8106), .BN(N8329), .C(N8697), .D(N7725));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2149 (.Y(N8308), .A(N7937), .B(N7700), .C(N8078));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2150 (.Y(N8132), .A(N8746), .B(N8308));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I2151 (.Y(N8235), .AN(N8614), .BN(N8773), .C(N8667), .D(N8372));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2152 (.Y(N8001), .A(N8781), .B(N7933), .C(N8171), .D(N8132));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2154 (.Y(N8677), .A(N8329), .B(N7937));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2155 (.Y(N7815), .A(N8195), .B(N8373));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2156 (.Y(N8018), .A(N7987), .B(N8307));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2157 (.Y(N8399), .A(N8666), .B(N7677));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2158 (.Y(N7762), .A(N8278), .B(N8399));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2159 (.Y(N8042), .A(N8383), .B(N8018), .C(N7762));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2160 (.Y(N7887), .A(N8254), .B(N8042));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2161 (.Y(N7976), .AN(N8392), .BN(N8501), .C(N7815), .D(N8677));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2162 (.Y(N8212), .A(N7976), .B(N7924));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2164 (.Y(N7742), .A(N8606), .B(N8518));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2165 (.Y(N8092), .AN(N8201), .BN(N8307), .C(N7742), .D(N8639));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2166 (.Y(N7858), .AN(N7937), .BN(N8373), .C(N7841), .D(N8380));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2167 (.Y(N8579), .A(N8215), .B(N7933), .C(N8408), .D(N7720));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2168 (.Y(inst_cellmath__197[16]), .A(N8435), .B(N8092), .C(N7858), .D(N8579));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2169 (.Y(N8391), .A(N8383), .B(N8638));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2170 (.Y(N7760), .A(N7754), .B(N7876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2171 (.Y(N8738), .A(N7800), .B(N7677));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2172 (.Y(N8594), .AN(N8738), .B(N8223), .C(N8408));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2173 (.Y(N8684), .A(N7821), .B(N8391));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2174 (.Y(N7974), .A(N7816), .B(N7760));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2175 (.Y(N8460), .AN(N8217), .B(N7937), .C(N8514));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2177 (.Y(N8556), .AN(N7931), .B(N8331), .C(N7974), .D(N8593));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2179 (.Y(N8165), .AN(N8373), .BN(N8215), .C(N8460), .D(N8594));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2181 (.Y(N8608), .A(N8215), .B(N8373), .C(N8728), .D(N8057));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2182 (.Y(N7736), .A(N8223), .B(N8638));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2183 (.Y(N7992), .A(N8331), .B(N8201));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2184 (.Y(N8224), .A(N8593), .B(N7754));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2185 (.Y(N7950), .A(N8738), .B(N7821));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2186 (.Y(N7802), .A(N8140));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2187 (.Y(N8053), .A(N7802), .B(N7950));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2188 (.Y(N8141), .A(N8284), .B(N7736), .C(N8047));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2189 (.Y(N7910), .A(N7992), .B(N8217), .C(N8224), .D(N8053));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2191 (.Y(N8367), .A(N8312), .B(N8057));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2192 (.Y(N8788), .A(N8154), .B(N8367));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2194 (.Y(N8652), .AN(N8025), .B(N8373), .C(N8788), .D(N8408));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2195 (.Y(N8512), .A(N7685), .B(N7755), .C(N8079), .D(N8047));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2198 (.Y(N7845), .A(N8615), .B(N7937));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2199 (.Y(N8569), .A(N8408));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2200 (.Y(N8669), .A(N8429), .B(N8528));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2201 (.Y(N8048), .AN(N8569), .B(N7949), .C(N8223), .D(N8435));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2202 (.Y(N8016), .A(N7933), .B(N8067));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2203 (.Y(N8135), .A(N8105), .B(N8047));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2204 (.Y(N8621), .A(N7802), .B(N8135));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2205 (.Y(N8486), .AN(N7902), .B(N8354), .C(N8048));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2206 (.Y(N8586), .AN(N8371), .BN(N8633), .C(N7845), .D(N8621));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2207 (.Y(N7961), .AN(N8669), .B(N8777), .C(N8486), .D(N8531));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2208 (.Y(inst_cellmath__195[0]), .AN(N7961), .B(N8016), .C(N8586));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2209 (.Y(N8547), .A(N8106), .B(N7687));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2210 (.Y(N8645), .A(N8350), .B(N8408));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2211 (.Y(N8352), .A(N8354), .B(N7908));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2212 (.Y(N8464), .A(N8307), .B(N8506), .C(N8115), .D(N8524));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2213 (.Y(N8694), .AN(N8645), .B(N8041), .C(N8352), .D(N7704));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2214 (.Y(N7680), .A(N8450), .B(N8025), .C(N8224), .D(N8694));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I2215 (.Y(N7943), .AN(N7804), .BN(N8547), .C(N7770), .D(N7680));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2216 (.Y(inst_cellmath__195[1]), .AN(N7943), .B(N7897), .C(N8464), .D(N7937));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2217 (.Y(N7859), .A(N7949), .B(N7985));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2218 (.Y(N8719), .A(N7841), .B(N7859));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2219 (.Y(N8192), .A(N8606), .B(N8041));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2220 (.Y(N7812), .A(N8627), .B(N8192));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2221 (.Y(N8059), .A(N7812), .B(N7694));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2222 (.Y(N8542), .AN(N7692), .BN(N8777), .C(N7813), .D(N7870));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2223 (.Y(N7920), .AN(N7780), .BN(N8115), .C(N8399), .D(N7831));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2224 (.Y(N8395), .AN(N8059), .B(N8526), .C(N8719), .D(N8737));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2225 (.Y(inst_cellmath__195[2]), .AN(N8395), .B(N8542), .C(N8016), .D(N7920));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2226 (.Y(N7995), .A(N7700), .B(N8236));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2227 (.Y(N7675), .A(N8050), .B(N7977));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2228 (.Y(N8434), .A(N8201), .B(N7987));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2229 (.Y(N8413), .A(N8391), .B(N8434));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2230 (.Y(N8662), .A(N7742), .B(N7995));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2231 (.Y(N7785), .A(N8239), .B(N8617));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2232 (.Y(N8040), .AN(N7675), .B(N8331), .C(N8413), .D(N8037));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2233 (.Y(N8755), .A(N8040), .B(N8035));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2234 (.Y(N8612), .AN(N8317), .B(N7785), .C(N8755), .D(N8662));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2235 (.Y(inst_cellmath__195[3]), .A(N8157), .B(N8126), .C(N8626), .D(N8612));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2236 (.Y(N7697), .A(N8177), .B(N8712));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2237 (.Y(N7916), .A(N8250), .B(N8041));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28267 (.Y(N8734), .A(N7916), .B(N7725), .C(N8764), .D(N8747));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2246 (.Y(N8301), .A(N8106), .B(N8526));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2248 (.Y(N7865), .A(N8531), .B(N8350));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2249 (.Y(N7917), .A(N8110), .B(N7985));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2250 (.Y(N8360), .A(N7865), .B(N7917));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2251 (.Y(N7990), .AN(N8050), .BN(N7800), .C(N8263), .D(N7908));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2253 (.Y(N7882), .A(N7987), .B(N8666), .C(N7990));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2256 (.Y(N7872), .A(N8043), .B(N8524));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2257 (.Y(N8205), .A(N8312), .B(N8768));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2258 (.Y(N8282), .A(N8611), .B(N8205));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2259 (.Y(N8009), .A(N8224), .B(N7675));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2260 (.Y(N8730), .A(N7995), .B(N7952));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2261 (.Y(N8104), .A(N7872), .B(N8009));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2262 (.Y(N7710), .AN(N7947), .B(N7803), .C(N8730), .D(N8514));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2263 (.Y(N8453), .A(N8035), .B(N7710));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2264 (.Y(N8166), .A(N7876), .B(N8648), .C(N8282));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2265 (.Y(N8070), .A(N8467), .B(N8166));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2266 (.Y(N7823), .AN(N8453), .B(N7792), .C(N8104), .D(N8785));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2267 (.Y(inst_cellmath__195[6]), .A(N8070), .B(N7823));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2268 (.Y(N8026), .A(N8435), .B(N7740));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2269 (.Y(N8264), .A(N8312), .B(N8291));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2270 (.Y(N8510), .A(N8633), .B(N8768));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2271 (.Y(N7773), .A(N8043), .B(N8373));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2272 (.Y(N7729), .A(N8532), .B(N7773));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2273 (.Y(N7794), .A(N8567), .B(N8269), .C(N8566));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2274 (.Y(N8180), .A(N8002), .B(N7804), .C(N8264));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2275 (.Y(N8277), .AN(N8363), .BN(N8350), .C(N8026), .D(N8510));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2276 (.Y(N8763), .A(N8180), .B(N7729), .C(N7933), .D(N7794));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2277 (.Y(inst_cellmath__195[7]), .A(N8277), .B(N7955), .C(N8763));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2278 (.Y(N8722), .A(N8145), .B(N8462));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2279 (.Y(N8678), .A(N8445), .B(N8722));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2280 (.Y(N8063), .A(N8037), .B(N8716));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2281 (.Y(N8153), .A(N8737), .B(N8502), .C(N8106), .D(N8312));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2282 (.Y(N8402), .A(N8236), .B(N8195), .C(N8768), .D(N8043));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2283 (.Y(N7765), .AN(N8648), .BN(N8250), .C(N7931), .D(N8678));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2284 (.Y(N8021), .AN(N8063), .B(N8531), .C(N8153), .D(N8408));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2285 (.Y(N8741), .A(N8649), .B(N8021));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2286 (.Y(N7888), .A(N7765), .B(N8741));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2287 (.Y(inst_cellmath__195[8]), .AN(N7888), .B(N8291), .C(N8402), .D(N8633));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2288 (.Y(N8273), .A(N8253), .B(N8651), .C(N8660));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2289 (.Y(N8553), .A(N8593), .B(N7780));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2290 (.Y(N8129), .A(N8115), .B(N8050));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2292 (.Y(N7999), .A(N8079), .B(N8553));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2294 (.Y(N7899), .A(N7902), .B(N8442), .C(N8728));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I28268 (.Y(N7861), .AN(N8273), .B(N8105), .C(N7899), .D(N8129));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2296 (.Y(N8330), .AN(N7999), .B(N8502), .C(N7861), .D(N8727));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2297 (.Y(inst_cellmath__195[9]), .AN(N8330), .B(N7872), .C(N7933));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2298 (.Y(N8498), .A(N8228), .B(N8200));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2299 (.Y(N7884), .A(N7704), .B(N7677));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2300 (.Y(N8226), .A(N8615), .B(N8721));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2301 (.Y(N8208), .A(N8584), .B(N8226));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2302 (.Y(N8686), .AN(N8089), .BN(N8633), .C(N7926), .D(N7773));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2303 (.Y(N8557), .AN(N8208), .B(N8374), .C(N7884), .D(N7865));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2304 (.Y(N7673), .A(N8557), .B(N8498));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2305 (.Y(inst_cellmath__195[10]), .AN(N7673), .B(N8392), .C(N8686), .D(N7780));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2306 (.Y(N8365), .A(N8777), .B(N8195));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2307 (.Y(N7738), .A(N8363), .B(N7833));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2308 (.Y(N8324), .A(N8239), .B(N8443));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2309 (.Y(N7695), .A(N8283), .B(N8081), .C(N8163));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2310 (.Y(N8189), .AN(N8478), .BN(N7720), .C(N8047), .D(N8365));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2311 (.Y(N8673), .AN(N7738), .B(N8236), .C(N8324), .D(N8373));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2312 (.Y(inst_cellmath__195[11]), .AN(N8673), .B(N8189), .C(N7695));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2313 (.Y(N8011), .A(N8502), .B(N8478));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2314 (.Y(N8345), .A(N8408), .B(N8164));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2315 (.Y(N7824), .A(N7727), .B(N7737));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2316 (.Y(N7693), .A(N8089), .B(N8777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2317 (.Y(N7935), .A(N8002), .B(N7693));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2318 (.Y(N8161), .AN(N8345), .B(N8171), .C(N7824), .D(N7803));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2319 (.Y(N8033), .AN(N8011), .B(N8666), .C(N7935), .D(N8456));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2320 (.Y(N8656), .A(N8197), .B(N8553), .C(N8192), .D(N8161));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28269 (.Y(inst_cellmath__195[12]), .A(N8272), .B(N8033), .C(N7705), .D(N8656));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2324 (.Y(N8086), .A(N7692), .B(N8291));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2325 (.Y(N8280), .A(N8250), .B(N8456));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2326 (.Y(N8624), .A(N8105), .B(N7752));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2327 (.Y(N8379), .A(N7897), .B(N7775), .C(N8606), .D(N8769));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2328 (.Y(N8006), .A(N8086), .B(N8298));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2329 (.Y(N8340), .AN(N8280), .B(N8593), .C(N8379), .D(N7876));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2330 (.Y(N8103), .A(N8415), .B(N7902), .C(N8728), .D(N8006));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2331 (.Y(N8770), .A(N8768), .B(N8506), .C(N8624));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2332 (.Y(N8196), .A(N8340), .B(N8770));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2333 (.Y(N7965), .A(N7921), .B(N8185), .C(N7753), .D(N8103));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2334 (.Y(inst_cellmath__195[13]), .A(N8196), .B(N7965));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2335 (.Y(N8784), .A(N8769), .B(N7692));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2336 (.Y(N8507), .A(N8185), .B(N8433));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2337 (.Y(N7726), .A(N8314), .B(N8405));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2338 (.Y(N8468), .A(N7931), .B(N8374), .C(N8784));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2339 (.Y(N7945), .AN(N8291), .BN(N8615), .C(N7865), .D(N8696));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2340 (.Y(N7682), .AN(N8317), .B(N8774), .C(N8468), .D(N8721));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2341 (.Y(N8420), .AN(N7876), .BN(N8050), .C(N7726), .D(N7682));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2342 (.Y(N7793), .A(N8392), .B(N8164), .C(N8420));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2343 (.Y(inst_cellmath__195[14]), .AN(N7793), .B(N8507), .C(N7945));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2344 (.Y(N8234), .A(N8043), .B(N8531));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2345 (.Y(N8010), .A(N7687), .B(N8329));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2346 (.Y(N8293), .A(N8252), .B(N8010));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2347 (.Y(N8545), .A(N8450), .B(N7727));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2348 (.Y(N7763), .A(N8146), .B(N8264));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2349 (.Y(N8151), .AN(N7704), .BN(N8050), .C(N8374), .D(N8234));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2350 (.Y(N8112), .A(N8089), .B(N8415), .C(N7692), .D(N7763));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2351 (.Y(N8258), .A(N8197), .B(N8044), .C(N7816), .D(N8317));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2352 (.Y(N7971), .A(N8383), .B(N8164), .C(N8293));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2353 (.Y(N8599), .A(N8258), .B(N7971));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2354 (.Y(inst_cellmath__195[15]), .AN(N8112), .B(N8545), .C(N8599), .D(N8151));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2355 (.Y(N7835), .A(N8781), .B(N8640));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2356 (.Y(N8109), .A(N8223), .B(N8110));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2357 (.Y(N8300), .A(N8578), .B(N8176));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2358 (.Y(N8522), .A(N8109), .B(N8300));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2359 (.Y(N7743), .A(N7870), .B(N7835), .C(N8614));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2360 (.Y(N7998), .AN(N7792), .B(N8373), .C(N8522), .D(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2361 (.Y(N7776), .A(N8329), .B(N7692));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2362 (.Y(N8477), .A(N8314), .B(N7776));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2363 (.Y(N7857), .AN(N7743), .B(N7780), .C(N8477), .D(N8307));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2364 (.Y(N8328), .A(N7967), .B(N7998), .C(N7857));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2365 (.Y(inst_cellmath__195[16]), .A(N7933), .B(N7848), .C(N7720), .D(N8328));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2366 (.Y(N8540), .A(N8721), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2367 (.Y(N8775), .A(N8110), .B(N7949));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2368 (.Y(N7717), .AN(N8089), .BN(N8526), .C(N7957), .D(N8129));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2369 (.Y(N8204), .AN(N7977), .BN(N8606), .C(N8540), .D(N8775));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2370 (.Y(N8072), .A(N8614), .B(N8163), .C(N8292), .D(N7727));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2371 (.Y(inst_cellmath__195[17]), .A(N8204), .B(N7717), .C(N8072));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2372 (.Y(N8358), .A(N8442), .B(N7740));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2373 (.Y(N8753), .A(N8555), .B(N8358));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2374 (.Y(N7898), .A(N8392), .B(N7985));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2375 (.Y(N8428), .A(N8596), .B(N7865));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2376 (.Y(N8610), .A(N7803), .B(N7933), .C(N8478));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2377 (.Y(N8711), .A(N8456), .B(N7677));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2378 (.Y(N8319), .A(N8037), .B(N8554), .C(N8753));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2379 (.Y(N7691), .A(N8207), .B(N8319));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2380 (.Y(N8187), .A(N7951), .B(N7891), .C(N8711));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2381 (.Y(N7911), .AN(N8187), .B(N8639), .C(N8610), .D(N7760));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2382 (.Y(inst_cellmath__195[18]), .AN(N7898), .B(N8428), .C(N7911), .D(N7691));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2384 (.Y(N7970), .A(N8531), .B(N8524));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2385 (.Y(N8671), .A(N8338), .B(N7720));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2386 (.Y(N8455), .A(N8228), .B(N8671));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28270 (.Y(N8653), .A(N8285), .B(N8105), .C(N8090), .D(N7884));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2389 (.Y(N8029), .AN(N8442), .BN(N8312), .C(N8569), .D(N7773));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2390 (.Y(N8511), .A(N8011), .B(N7970), .C(N8267));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2391 (.Y(N8120), .AN(N8653), .B(N8721), .C(N8455), .D(N8506));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2392 (.Y(N8138), .A(N7933), .B(N8593));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2393 (.Y(N7730), .A(N8120), .B(N8138));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2394 (.Y(inst_cellmath__195[19]), .AN(N8126), .B(N8511), .C(N7730), .D(N8029));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2395 (.Y(N7750), .A(N8569), .B(N8764));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2396 (.Y(N8622), .A(N8128), .B(N7870), .C(N8376));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2397 (.Y(N8725), .A(N8037), .B(N8067));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2398 (.Y(N8065), .A(N8354), .B(N8254), .C(N7962));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2399 (.Y(N8447), .A(N7931), .B(N8216), .C(N8725), .D(N8587));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2400 (.Y(N8295), .A(N8065), .B(N8447));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2401 (.Y(N8779), .AN(N7750), .BN(N7766), .C(N8622), .D(N8295));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2402 (.Y(inst_cellmath__195[20]), .A(N7933), .B(N8371), .C(N8312), .D(N8779));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2403 (.Y(N8101), .A(N8378), .B(N7933), .C(N7985));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2405 (.Y(N7839), .A(N8666), .B(N7977));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2406 (.Y(N8175), .A(N8207), .B(N8698), .C(N7839));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2407 (.Y(N8664), .AN(N7849), .B(N8711), .C(N8154));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2408 (.Y(N8523), .AN(N8298), .B(N8727), .C(N8664), .D(N7720));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2409 (.Y(N7819), .A(N7803), .B(N7692), .C(N8175));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28271 (.Y(inst_cellmath__195[21]), .A(N8629), .B(N8101), .C(N7819), .D(N8523));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2412 (.Y(N8543), .A(N7800), .B(N7775));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2413 (.Y(N7919), .A(N8125), .B(N7892));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2414 (.Y(N8396), .A(N8564), .B(N7814), .C(N8532));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2415 (.Y(N8255), .AN(N8524), .BN(N8501), .C(N7900), .D(N8543));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I2416 (.Y(N7886), .AN(N8025), .BN(N8528), .C(N7987), .D(N8396));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2417 (.Y(N8597), .A(N8245), .B(N8164), .C(N8255));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2418 (.Y(N8210), .AN(N8721), .BN(N8633), .C(N8298), .D(N8597));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2419 (.Y(inst_cellmath__195[22]), .AN(N7886), .B(N7679), .C(N8210), .D(N7919));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2420 (.Y(N7786), .A(N8110), .B(N7833));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2421 (.Y(N8127), .A(N8391), .B(N7697));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2422 (.Y(N8474), .AN(N8227), .B(N8115), .C(N8127), .D(N8606));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2423 (.Y(N7855), .A(N8767), .B(N7845));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2424 (.Y(N8326), .AN(N8176), .BN(N8737), .C(N8400), .D(N7786));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2425 (.Y(N7953), .A(N8725), .B(N8543), .C(N7995), .D(N8474));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2426 (.Y(N7698), .AN(N8375), .B(N8774), .C(N7855), .D(N8777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2427 (.Y(N8190), .A(N7953), .B(N7698));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2428 (.Y(inst_cellmath__195[23]), .A(N8326), .B(N8190));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2429 (.Y(N8302), .AN(N8176), .BN(N8769), .C(N7932), .D(N8109));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2430 (.Y(N8647), .A(N8171), .B(N7687), .C(N7933));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2431 (.Y(N8036), .AN(N8435), .B(N8647), .C(N7835));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2432 (.Y(N7890), .A(N8245), .B(N7902));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2433 (.Y(N7672), .A(N8298), .B(N7890));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2434 (.Y(N8658), .A(N8339), .B(N8002), .C(N7865), .D(N7884));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I2435 (.Y(N8410), .AN(N8264), .BN(N8334), .C(N7672), .D(N8302));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2436 (.Y(N7779), .A(N8658), .B(N8410));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2437 (.Y(inst_cellmath__195[24]), .A(N8036), .B(N7779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2438 (.Y(N8124), .A(N8640), .B(N8712));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2439 (.Y(N8362), .A(N8435), .B(N8526));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2440 (.Y(N7735), .A(N8312), .B(N7937));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2441 (.Y(N8088), .A(N7754), .B(N8050));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2442 (.Y(N8426), .A(N8047), .B(N8738));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2443 (.Y(N7799), .AN(N8088), .B(N8223), .C(N8362), .D(N8593));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2444 (.Y(N7873), .A(N7696), .B(N7908), .C(N8124), .D(N7970));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2445 (.Y(N8243), .AN(N7679), .BN(N8426), .C(N8263), .D(N7735));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I2446 (.Y(inst_cellmath__195[25]), .AN(N8139), .BN(N7799), .C(N7873), .D(N8243));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2447 (.Y(N8071), .A(N8195), .B(N8215));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2448 (.Y(N8466), .A(N8041), .B(N7775));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2449 (.Y(N8027), .A(N8483), .B(N8466));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2450 (.Y(N8356), .AN(N8118), .B(N8329), .C(N8721));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2451 (.Y(N8469), .AN(N8071), .B(N8378), .C(N8027), .D(N8593));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2452 (.Y(N8218), .A(N8094), .B(N8124), .C(N8356));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2453 (.Y(N8701), .A(N8785), .B(N7771), .C(N8587), .D(N8469));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2454 (.Y(inst_cellmath__195[26]), .A(N8218), .B(N8701));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2455 (.Y(N8723), .A(N8483), .B(N8698));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2456 (.Y(N8098), .A(N7675), .B(N8380));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2457 (.Y(N8238), .A(N7947), .B(N7900));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2458 (.Y(N8484), .A(N8785), .B(N8374));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2459 (.Y(N7867), .A(N8371), .B(N8777), .C(N8723));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2460 (.Y(N8444), .AN(N8238), .BN(N8484), .C(N7771), .D(N8098));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2461 (.Y(inst_cellmath__195[27]), .AN(N7867), .B(N8195), .C(N8444), .D(N8223));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2462 (.Y(N8463), .AN(N7992), .B(N8338), .C(N8057));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2465 (.Y(N8417), .A(N7716), .B(N7900), .C(N7892));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I28272 (.Y(N7941), .A(N8785), .B(N7891), .C(N8217), .D(N8463));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2467 (.Y(N8173), .A(N7736), .B(N8698), .C(N8374), .D(N7941));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2468 (.Y(inst_cellmath__195[28]), .A(N8417), .B(N8173));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2469 (.Y(N7904), .A(N7692), .B(N8223));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2470 (.Y(N7956), .A(N7908), .B(N8747));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I2471 (.Y(N8438), .AN(N8593), .BN(N8067), .C(N8483), .D(N8374));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I10077 (.Y(N7809), .A(N7685), .B(N7792), .C(N7904));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2473 (.Y(N8288), .A(N7778), .B(N7727), .C(N7947));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2474 (.Y(inst_cellmath__195[29]), .A(N7956), .B(N8438), .C(N8288), .D(N7809));
INVX3 inst_cellmath__198_0_I2475 (.Y(N10506), .A(inst_cellmath__61[1]));
INVXL inst_cellmath__198_0_I9934 (.Y(N22556), .A(N10506));
INVXL inst_cellmath__198_0_I9939 (.Y(N22561), .A(N22556));
XNOR2X1 inst_cellmath__198_0_I28273 (.Y(N9963), .A(N7631), .B(N736));
NOR2XL node_cs_const1_cs_A_I10767 (.Y(N22635), .A(N7131), .B(N7352));
XNOR2X1 node_cs_const1_cs_A_I10768 (.Y(N10287), .A(N7631), .B(N22635));
INVX3 inst_cellmath__198_0_I2485 (.Y(N10490), .A(inst_cellmath__61[5]));
XNOR2X1 inst_cellmath__198_0_I10081 (.Y(N10458), .A(N7631), .B(N740));
NOR2XL node_cs_const1_cs_A_I10769 (.Y(N22642), .A(N7131), .B(N7371));
XNOR2X1 node_cs_const1_cs_A_I10770 (.Y(N10433), .A(N7631), .B(N22642));
INVX3 inst_cellmath__198_0_I2492 (.Y(N10472), .A(inst_cellmath__61[11]));
INVX3 inst_cellmath__198_0_I2495 (.Y(N10039), .A(inst_cellmath__61[12]));
INVX3 inst_cellmath__198_0_I2498 (.Y(N10515), .A(inst_cellmath__61[13]));
INVX2 inst_cellmath__198_0_I2501 (.Y(N10016), .A(inst_cellmath__61[14]));
INVX2 inst_cellmath__198_0_I2503 (.Y(N10204), .A(inst_cellmath__61[15]));
INVX2 inst_cellmath__198_0_I2504 (.Y(N10486), .A(inst_cellmath__115__W1[0]));
XNOR2X1 inst_cellmath__198_0_I9988 (.Y(N10181), .A(N7631), .B(N733));
INVX2 inst_cellmath__198_0_I9944 (.Y(N22566), .A(N10181));
INVXL inst_cellmath__198_0_I9952 (.Y(N22574), .A(N22566));
INVX1 inst_cellmath__198_0_I9951 (.Y(N22573), .A(N22566));
INVXL inst_cellmath__198_0_I9950 (.Y(N22572), .A(N22566));
INVX1 inst_cellmath__198_0_I9946 (.Y(N22568), .A(N22566));
INVX2 inst_cellmath__198_0_I9945 (.Y(N22567), .A(N22566));
NOR2XL inst_cellmath__198_0_I2510 (.Y(N9981), .A(N22574), .B(N9963));
NOR2XL inst_cellmath__198_0_I2511 (.Y(N10246), .A(N10287), .B(N22573));
NOR2BX1 inst_cellmath__198_0_I2512 (.Y(N10535), .AN(inst_cellmath__61[5]), .B(N22573));
NOR2BXL inst_cellmath__198_0_I2513 (.Y(N10171), .AN(inst_cellmath__61[6]), .B(N10181));
NOR2XL inst_cellmath__198_0_I2514 (.Y(N10443), .A(N10458), .B(N22567));
NOR2XL inst_cellmath__198_0_I2515 (.Y(N10093), .A(N3665), .B(N22567));
NOR2XL inst_cellmath__198_0_I2516 (.Y(N10359), .A(N10433), .B(N22567));
NOR2BX1 inst_cellmath__198_0_I2517 (.Y(N10015), .AN(inst_cellmath__61[10]), .B(N22573));
NOR2XL inst_cellmath__198_0_I2518 (.Y(N10280), .A(N22573), .B(N10472));
NOR2BXL inst_cellmath__198_0_I2519 (.Y(N9933), .AN(inst_cellmath__61[12]), .B(N22573));
NOR2XL inst_cellmath__198_0_I2520 (.Y(N10203), .A(N22572), .B(N10515));
NOR2X2 inst_cellmath__198_0_I2521 (.Y(N10483), .A(N10016), .B(N22567));
NOR2BX2 inst_cellmath__198_0_I2522 (.Y(N10126), .AN(inst_cellmath__61[15]), .B(N22568));
OR2XL inst_cellmath__198_0_I2523 (.Y(N10168), .A(N10486), .B(N22568));
NOR2XL inst_cellmath__198_0_I2524 (.Y(N10084), .A(N10506), .B(N3661));
NOR2XL inst_cellmath__198_0_I2525 (.Y(N10347), .A(N10506), .B(N9963));
NOR2XL inst_cellmath__198_0_I2526 (.Y(N9999), .A(N10506), .B(N10287));
NOR2XL inst_cellmath__198_0_I2527 (.Y(N10267), .A(N10506), .B(N10490));
NOR2XL inst_cellmath__198_0_I2528 (.Y(N9920), .A(N10506), .B(N3659));
NOR2XL inst_cellmath__198_0_I2529 (.Y(N10189), .A(N10506), .B(N10458));
NOR2XL inst_cellmath__198_0_I2530 (.Y(N10469), .A(N10506), .B(N3665));
NOR2XL inst_cellmath__198_0_I2531 (.Y(N10111), .A(N10506), .B(N10433));
NOR2XL inst_cellmath__198_0_I2532 (.Y(N10380), .A(N10506), .B(N3657));
NOR2XL inst_cellmath__198_0_I2533 (.Y(N10036), .A(N10506), .B(N10472));
NOR2XL inst_cellmath__198_0_I2534 (.Y(N10304), .A(N10506), .B(N10039));
NOR2X1 inst_cellmath__198_0_I2535 (.Y(N9953), .A(N10506), .B(N10515));
NOR2X1 inst_cellmath__198_0_I2536 (.Y(N10223), .A(N10506), .B(N10016));
NOR2XL inst_cellmath__198_0_I2537 (.Y(N10508), .A(N10506), .B(N10204));
NOR2X2 inst_cellmath__198_0_I9980 (.Y(N22602), .A(N10486), .B(N10506));
INVX1 inst_cellmath__198_0_I9981 (.Y(N10305), .A(N22602));
NOR2XL inst_cellmath__198_0_I2540 (.Y(N10448), .A(N3661), .B(N9963));
NOR2XL inst_cellmath__198_0_I2541 (.Y(N10098), .A(N3661), .B(N10287));
NOR2XL inst_cellmath__198_0_I2542 (.Y(N10365), .A(N3661), .B(N10490));
NOR2XL inst_cellmath__198_0_I2543 (.Y(N10021), .A(N3661), .B(N3659));
NOR2XL inst_cellmath__198_0_I2544 (.Y(N10290), .A(N3661), .B(N10458));
NOR2XL inst_cellmath__198_0_I2545 (.Y(N9939), .A(N3661), .B(N3665));
NOR2XL inst_cellmath__198_0_I2546 (.Y(N10211), .A(N3661), .B(N10433));
NOR2XL inst_cellmath__198_0_I2547 (.Y(N10494), .A(N3661), .B(N3657));
NOR2XL inst_cellmath__198_0_I2548 (.Y(N10130), .A(N3661), .B(N10472));
NOR2XL inst_cellmath__198_0_I2549 (.Y(N10401), .A(N3661), .B(N10039));
NOR2X2 inst_cellmath__198_0_I2550 (.Y(N10054), .A(N3661), .B(N10515));
NOR2XL inst_cellmath__198_0_I2551 (.Y(N10324), .A(N3661), .B(N10016));
NOR2XL inst_cellmath__198_0_I2552 (.Y(N9975), .A(N3661), .B(N10204));
OR2XL inst_cellmath__198_0_I2553 (.Y(N10439), .A(N10486), .B(N3661));
INVXL inst_cellmath__198_0_I2554 (.Y(N10008), .A(N9963));
NOR2XL inst_cellmath__198_0_I2555 (.Y(N9927), .A(N10287), .B(N9963));
NOR2XL inst_cellmath__198_0_I2556 (.Y(N10195), .A(N10490), .B(N9963));
NOR2XL inst_cellmath__198_0_I2557 (.Y(N10476), .A(N3659), .B(N9963));
NOR2XL inst_cellmath__198_0_I2558 (.Y(N10118), .A(N10458), .B(N9963));
NOR2XL inst_cellmath__198_0_I2559 (.Y(N10388), .A(N3665), .B(N9963));
NOR2XL inst_cellmath__198_0_I2560 (.Y(N10041), .A(N10433), .B(N9963));
NOR2XL inst_cellmath__198_0_I2561 (.Y(N10311), .A(N3657), .B(N9963));
NOR2XL inst_cellmath__198_0_I2562 (.Y(N9964), .A(N10472), .B(N9963));
NOR2XL inst_cellmath__198_0_I2563 (.Y(N10230), .A(N9963), .B(N10039));
NOR2X1 inst_cellmath__198_0_I2564 (.Y(N10518), .A(N9963), .B(N10515));
NOR2X1 inst_cellmath__198_0_I2565 (.Y(N10154), .A(N10016), .B(N9963));
NOR2XL inst_cellmath__198_0_I2566 (.Y(N10421), .A(N10204), .B(N9963));
OR2XL inst_cellmath__198_0_I2567 (.Y(N9955), .A(N10486), .B(N9963));
INVXL inst_cellmath__198_0_I2568 (.Y(N10459), .A(N10287));
NOR2XL inst_cellmath__198_0_I2569 (.Y(N10373), .A(N10287), .B(N10490));
NOR2XL inst_cellmath__198_0_I2570 (.Y(N10031), .A(N10287), .B(N3659));
NOR2XL inst_cellmath__198_0_I2571 (.Y(N10298), .A(N10458), .B(N10287));
NOR2XL inst_cellmath__198_0_I2572 (.Y(N9947), .A(N3665), .B(N10287));
NOR2XL inst_cellmath__198_0_I2573 (.Y(N10219), .A(N10433), .B(N10287));
NOR2XL inst_cellmath__198_0_I2574 (.Y(N10502), .A(N3657), .B(N10287));
NOR2XL inst_cellmath__198_0_I2575 (.Y(N10137), .A(N10287), .B(N10472));
NOR2XL inst_cellmath__198_0_I2576 (.Y(N10409), .A(N10287), .B(N10039));
NOR2XL inst_cellmath__198_0_I2577 (.Y(N10062), .A(N10287), .B(N10515));
NOR2XL inst_cellmath__198_0_I2578 (.Y(N10329), .A(N10016), .B(N10287));
NOR2XL inst_cellmath__198_0_I2579 (.Y(N9982), .A(N10204), .B(N10287));
OR2XL inst_cellmath__198_0_I2580 (.Y(N10091), .A(N10486), .B(N10287));
INVXL inst_cellmath__198_0_I2581 (.Y(N10017), .A(N10490));
NOR2XL inst_cellmath__198_0_I2582 (.Y(N9934), .A(N10490), .B(N3659));
NOR2XL inst_cellmath__198_0_I2583 (.Y(N10205), .A(N10490), .B(N10458));
NOR2XL inst_cellmath__198_0_I2584 (.Y(N10487), .A(N10490), .B(N3665));
NOR2XL inst_cellmath__198_0_I2585 (.Y(N10127), .A(N10490), .B(N10433));
NOR2X2 inst_cellmath__198_0_I2586 (.Y(N10396), .A(N3657), .B(N10490));
NOR2X2 inst_cellmath__198_0_I2587 (.Y(N10049), .A(N10472), .B(N10490));
NOR2X2 inst_cellmath__198_0_I2588 (.Y(N10319), .A(N10039), .B(N10490));
NOR2XL inst_cellmath__198_0_I2589 (.Y(N9970), .A(N10515), .B(N10490));
NOR2XL inst_cellmath__198_0_I2590 (.Y(N10237), .A(N10490), .B(N10016));
NOR2XL inst_cellmath__198_0_I2591 (.Y(N10526), .A(N10204), .B(N10490));
OR2XL inst_cellmath__198_0_I2592 (.Y(N10224), .A(N10490), .B(N10486));
NOR2XL inst_cellmath__198_0_I2594 (.Y(N10470), .A(N3659), .B(N10458));
NOR2XL inst_cellmath__198_0_I2595 (.Y(N10112), .A(N3659), .B(N3665));
NOR2XL inst_cellmath__198_0_I2596 (.Y(N10382), .A(N3659), .B(N10433));
NOR2X1 inst_cellmath__198_0_I2597 (.Y(N10037), .A(N3657), .B(N3659));
NOR2X2 inst_cellmath__198_0_I2598 (.Y(N10306), .A(N10472), .B(N3659));
NOR2XL inst_cellmath__198_0_I2599 (.Y(N9958), .A(N3659), .B(N10039));
NOR2XL inst_cellmath__198_0_I2600 (.Y(N10226), .A(N3659), .B(N10515));
NOR2XL inst_cellmath__198_0_I2601 (.Y(N10511), .A(N3659), .B(N10016));
NOR2XL inst_cellmath__198_0_I2602 (.Y(N10149), .A(N10204), .B(N3659));
OR2XL inst_cellmath__198_0_I2603 (.Y(N10356), .A(N10486), .B(N3659));
INVXL inst_cellmath__198_0_I2604 (.Y(N10179), .A(N10458));
NOR2XL inst_cellmath__198_0_I2605 (.Y(N10102), .A(N3665), .B(N10458));
NOR2XL inst_cellmath__198_0_I2606 (.Y(N10368), .A(N10458), .B(N10433));
NOR2X1 inst_cellmath__198_0_I2607 (.Y(N10024), .A(N10458), .B(N3657));
NOR2XL inst_cellmath__198_0_I2608 (.Y(N10294), .A(N10458), .B(N10472));
NOR2XL inst_cellmath__198_0_I2609 (.Y(N9942), .A(N10039), .B(N10458));
NOR2XL inst_cellmath__198_0_I2610 (.Y(N10214), .A(N10458), .B(N10515));
NOR2XL inst_cellmath__198_0_I2611 (.Y(N10498), .A(N10458), .B(N10016));
NOR2XL inst_cellmath__198_0_I2612 (.Y(N10133), .A(N10204), .B(N10458));
OR2XL inst_cellmath__198_0_I2613 (.Y(N10509), .A(N10486), .B(N10458));
NOR2XL inst_cellmath__198_0_I2615 (.Y(N10090), .A(N3665), .B(N10433));
NOR2XL inst_cellmath__198_0_I2616 (.Y(N10353), .A(N3665), .B(N3657));
NOR2XL inst_cellmath__198_0_I2617 (.Y(N10011), .A(N3665), .B(N10472));
NOR2XL inst_cellmath__198_0_I2618 (.Y(N10276), .A(N3665), .B(N10039));
NOR2XL inst_cellmath__198_0_I2619 (.Y(N9929), .A(N3665), .B(N10515));
NOR2XL inst_cellmath__198_0_I2620 (.Y(N10198), .A(N3665), .B(N10016));
NOR2XL inst_cellmath__198_0_I2621 (.Y(N10478), .A(N3665), .B(N10204));
OR2XL inst_cellmath__198_0_I2622 (.Y(N10012), .A(N10486), .B(N3665));
INVX1 inst_cellmath__198_0_I2623 (.Y(N10521), .A(N10433));
NOR2XL inst_cellmath__198_0_I2624 (.Y(N10423), .A(N3657), .B(N10433));
NOR2XL inst_cellmath__198_0_I2625 (.Y(N10078), .A(N10472), .B(N10433));
NOR2XL inst_cellmath__198_0_I2626 (.Y(N10342), .A(N10039), .B(N10433));
NOR2XL inst_cellmath__198_0_I2627 (.Y(N9995), .A(N10433), .B(N10515));
NOR2XL inst_cellmath__198_0_I2628 (.Y(N10263), .A(N10433), .B(N10016));
NOR2XL inst_cellmath__198_0_I2629 (.Y(N9914), .A(N10204), .B(N10433));
OR2XL inst_cellmath__198_0_I2630 (.Y(N10147), .A(N10486), .B(N10433));
NOR2XL inst_cellmath__198_0_I2632 (.Y(N10505), .A(N3657), .B(N10472));
NOR2XL inst_cellmath__198_0_I2633 (.Y(N10140), .A(N10039), .B(N3657));
NOR2XL inst_cellmath__198_0_I2634 (.Y(N10413), .A(N3657), .B(N10515));
NOR2XL inst_cellmath__198_0_I2635 (.Y(N10066), .A(N3657), .B(N10016));
NOR2XL inst_cellmath__198_0_I2636 (.Y(N10334), .A(N10204), .B(N3657));
OR2XL inst_cellmath__198_0_I2637 (.Y(N10278), .A(N10486), .B(N3657));
INVXL inst_cellmath__198_0_I2638 (.Y(N10362), .A(N10472));
NOR2XL inst_cellmath__198_0_I2639 (.Y(N10286), .A(N10472), .B(N10039));
NOR2XL inst_cellmath__198_0_I2640 (.Y(N9937), .A(N10472), .B(N10515));
NOR2XL inst_cellmath__198_0_I2641 (.Y(N10208), .A(N10472), .B(N10016));
NOR2XL inst_cellmath__198_0_I2642 (.Y(N10489), .A(N10472), .B(N10204));
OR2XL inst_cellmath__198_0_I2643 (.Y(N10416), .A(N10472), .B(N10486));
INVXL inst_cellmath__198_0_I2644 (.Y(N10528), .A(N10039));
NOR2XL inst_cellmath__198_0_I2645 (.Y(N10432), .A(N10039), .B(N10515));
NOR2XL inst_cellmath__198_0_I2646 (.Y(N10086), .A(N10039), .B(N10016));
NOR2XL inst_cellmath__198_0_I2647 (.Y(N10349), .A(N10039), .B(N10204));
OR2XL inst_cellmath__198_0_I2648 (.Y(N9930), .A(N10039), .B(N10486));
INVXL inst_cellmath__198_0_I2649 (.Y(N10384), .A(N10515));
NOR2XL inst_cellmath__198_0_I2650 (.Y(N10308), .A(N10016), .B(N10515));
NOR2XL inst_cellmath__198_0_I2651 (.Y(N9960), .A(N10204), .B(N10515));
OR2XL inst_cellmath__198_0_I2652 (.Y(N10070), .A(N10486), .B(N10515));
INVXL inst_cellmath__198_0_I2653 (.Y(N9992), .A(N10016));
NOR2XL inst_cellmath__198_0_I2654 (.Y(N9909), .A(N10204), .B(N10016));
OR2XL inst_cellmath__198_0_I2655 (.Y(N10200), .A(N10486), .B(N10016));
INVXL inst_cellmath__198_0_I2656 (.Y(N9945), .A(N10204));
ADDHX1 inst_cellmath__198_0_I2657 (.CO(N10481), .S(N10336), .A(N3662), .B(N10084));
ADDHXL inst_cellmath__198_0_I2658 (.CO(N10122), .S(N9989), .A(N10246), .B(N10347));
ADDHX1 inst_cellmath__198_0_I2659 (.CO(N10393), .S(N10254), .A(N10535), .B(N10448));
ADDFX1 inst_cellmath__198_0_I2660 (.CO(N10043), .S(N9906), .A(N9999), .B(N10008), .CI(N10122));
ADDHX1 inst_cellmath__198_0_I2661 (.CO(N10316), .S(N10177), .A(N10171), .B(N10267));
ADDFXL inst_cellmath__198_0_I2662 (.CO(N9967), .S(N10449), .A(N10098), .B(N10393), .CI(N10177));
ADDHX1 inst_cellmath__198_0_I2663 (.CO(N10232), .S(N10100), .A(N10365), .B(N10443));
ADDFX1 inst_cellmath__198_0_I2664 (.CO(N10523), .S(N10367), .A(N9927), .B(N9920), .CI(N10459));
ADDFXL inst_cellmath__198_0_I2665 (.CO(N10157), .S(N10022), .A(N10100), .B(N10316), .CI(N9967));
ADDHX1 inst_cellmath__198_0_I2666 (.CO(N10425), .S(N10292), .A(N10021), .B(N10189));
ADDFX1 inst_cellmath__198_0_I2667 (.CO(N10081), .S(N9941), .A(N10093), .B(N10195), .CI(N10232));
ADDFX1 inst_cellmath__198_0_I2668 (.CO(N10344), .S(N10212), .A(N10523), .B(N10292), .CI(N9941));
ADDHX1 inst_cellmath__198_0_I2669 (.CO(N9997), .S(N10496), .A(N10017), .B(N10290));
ADDFX1 inst_cellmath__198_0_I2670 (.CO(N10265), .S(N10132), .A(N10476), .B(N10359), .CI(N10373));
ADDFX1 inst_cellmath__198_0_I2671 (.CO(N9916), .S(N10402), .A(N10425), .B(N10469), .CI(N10496));
ADDFX1 inst_cellmath__198_0_I2672 (.CO(N10187), .S(N10056), .A(N10132), .B(N10081), .CI(N10402));
ADDHX1 inst_cellmath__198_0_I2673 (.CO(N10466), .S(N10326), .A(N10015), .B(N10118));
ADDFX1 inst_cellmath__198_0_I2674 (.CO(N10109), .S(N9976), .A(N9939), .B(N10111), .CI(N10031));
ADDFX1 inst_cellmath__198_0_I2675 (.CO(N10376), .S(N10242), .A(N10326), .B(N9997), .CI(N10265));
ADDFX1 inst_cellmath__198_0_I2676 (.CO(N10034), .S(N10532), .A(N9976), .B(N9916), .CI(N10242));
ADDHX1 inst_cellmath__198_0_I2677 (.CO(N10301), .S(N10164), .A(N3660), .B(N9934));
ADDFXL inst_cellmath__198_0_I2678 (.CO(N9951), .S(N10436), .A(N10211), .B(N10380), .CI(N10280));
ADDFX1 inst_cellmath__198_0_I2679 (.CO(N10221), .S(N10089), .A(N10298), .B(N10388), .CI(N10164));
ADDFXL inst_cellmath__198_0_I2680 (.CO(N10507), .S(N10351), .A(N10109), .B(N10466), .CI(N10436));
ADDFXL inst_cellmath__198_0_I2681 (.CO(N10143), .S(N10009), .A(N10376), .B(N10089), .CI(N10351));
ADDHX1 inst_cellmath__198_0_I2682 (.CO(N10414), .S(N10275), .A(N10494), .B(N10205));
ADDFX1 inst_cellmath__198_0_I2683 (.CO(N10068), .S(N9928), .A(N10036), .B(N10041), .CI(N9933));
ADDFX1 inst_cellmath__198_0_I2684 (.CO(N10335), .S(N10196), .A(N10301), .B(N9947), .CI(N10275));
ADDFX1 inst_cellmath__198_0_I2685 (.CO(N9986), .S(N10477), .A(N9928), .B(N9951), .CI(N10221));
ADDFX1 inst_cellmath__198_0_I2686 (.CO(N10252), .S(N10119), .A(N10507), .B(N10196), .CI(N10477));
ADDHXL inst_cellmath__198_0_I2687 (.CO(N9903), .S(N10389), .A(N10130), .B(N10179));
ADDFX1 inst_cellmath__198_0_I2688 (.CO(N10173), .S(N10042), .A(N10304), .B(N10470), .CI(N10203));
ADDFX1 inst_cellmath__198_0_I2689 (.CO(N10447), .S(N10312), .A(N10311), .B(N10219), .CI(N10487));
ADDFX1 inst_cellmath__198_0_I2690 (.CO(N10097), .S(N9965), .A(N10389), .B(N10414), .CI(N10068));
ADDFX1 inst_cellmath__198_0_I2691 (.CO(N10363), .S(N10231), .A(N10335), .B(N10042), .CI(N10312));
ADDFX1 inst_cellmath__198_0_I2692 (.CO(N10020), .S(N10519), .A(N9986), .B(N9965), .CI(N10231));
ADDHX1 inst_cellmath__198_0_I2693 (.CO(N10288), .S(N10155), .A(N9953), .B(N10483));
ADDFX1 inst_cellmath__198_0_I2694 (.CO(N9938), .S(N10422), .A(N9964), .B(N10401), .CI(N10502));
ADDFX1 inst_cellmath__198_0_I2695 (.CO(N10209), .S(N10077), .A(N10127), .B(N10112), .CI(N9903));
ADDFX1 inst_cellmath__198_0_I2696 (.CO(N10491), .S(N10341), .A(N10447), .B(N10155), .CI(N10173));
ADDFX1 inst_cellmath__198_0_I2697 (.CO(N10129), .S(N9994), .A(N10422), .B(N10077), .CI(N10097));
ADDFXL inst_cellmath__198_0_I2698 (.CO(N10399), .S(N10261), .A(N10363), .B(N10341), .CI(N9994));
ADDHXL inst_cellmath__198_0_I2699 (.CO(N10052), .S(N9912), .A(N10054), .B(N10396));
ADDFXL inst_cellmath__198_0_I2700 (.CO(N10322), .S(N10185), .A(N10223), .B(N10126), .CI(N10230));
ADDFX1 inst_cellmath__198_0_I2701 (.CO(N9973), .S(N10460), .A(N10102), .B(N10382), .CI(N10137));
ADDFHXL inst_cellmath__198_0_I2702 (.CO(N10239), .S(N10106), .A(N10288), .B(N3666), .CI(N9912));
ADDFX1 inst_cellmath__198_0_I2703 (.CO(N10529), .S(N10374), .A(N10185), .B(N9938), .CI(N10209));
ADDFX1 inst_cellmath__198_0_I2704 (.CO(N10162), .S(N10032), .A(N10460), .B(N10106), .CI(N10491));
ADDFX1 inst_cellmath__198_0_I2705 (.CO(N10434), .S(N10299), .A(N10129), .B(N10374), .CI(N10032));
XNOR2X1 inst_cellmath__198_0_I2706 (.Y(N9948), .A(N10037), .B(N10508));
OR2XL inst_cellmath__198_0_I2707 (.Y(N10087), .A(N10508), .B(N10037));
ADDFXL inst_cellmath__198_0_I2708 (.CO(N10004), .S(N10503), .A(N10049), .B(N10518), .CI(N10324));
ADDFX1 inst_cellmath__198_0_I2709 (.CO(N10271), .S(N10138), .A(N10409), .B(N10368), .CI(N10168));
ADDFHXL inst_cellmath__198_0_I2710 (.CO(N9923), .S(N10410), .A(N9948), .B(N10052), .CI(N10322));
ADDFHXL inst_cellmath__198_0_I2711 (.CO(N10192), .S(N10063), .A(N10503), .B(N9973), .CI(N10239));
ADDFXL inst_cellmath__198_0_I2712 (.CO(N10473), .S(N10331), .A(N10410), .B(N10138), .CI(N10529));
ADDFHXL inst_cellmath__198_0_I2713 (.CO(N10115), .S(N9983), .A(N10162), .B(N10063), .CI(N10331));
ADDFX1 inst_cellmath__198_0_I2714 (.CO(N10386), .S(N10247), .A(N10306), .B(N10319), .CI(N9975));
ADDFXL inst_cellmath__198_0_I2715 (.CO(N10040), .S(N10538), .A(N10024), .B(N10154), .CI(N10090));
ADDFHXL inst_cellmath__198_0_I2716 (.CO(N10310), .S(N10172), .A(N10521), .B(N10305), .CI(N10062));
ADDFXL inst_cellmath__198_0_I2717 (.CO(N9961), .S(N10445), .A(N10004), .B(N10087), .CI(N10271));
ADDFX1 inst_cellmath__198_0_I2718 (.CO(N10228), .S(N10096), .A(N10172), .B(N10538), .CI(N10247));
ADDFHXL inst_cellmath__198_0_I2719 (.CO(N10516), .S(N10361), .A(N9923), .B(N10192), .CI(N10445));
ADDFHXL inst_cellmath__198_0_I2720 (.CO(N10151), .S(N10018), .A(N10096), .B(N10473), .CI(N10361));
ADDFXL inst_cellmath__198_0_I2721 (.CO(N10419), .S(N10284), .A(N10294), .B(N9958), .CI(N9970));
ADDFX1 inst_cellmath__198_0_I2722 (.CO(N10075), .S(N9935), .A(N10439), .B(N10421), .CI(N10329));
ADDFHXL inst_cellmath__198_0_I2723 (.CO(N10339), .S(N10206), .A(N10386), .B(N10353), .CI(N10310));
ADDFX1 inst_cellmath__198_0_I2724 (.CO(N9993), .S(N10488), .A(N10284), .B(N10040), .CI(N9935));
ADDFHXL inst_cellmath__198_0_I2725 (.CO(N10260), .S(N10128), .A(N9961), .B(N10206), .CI(N10228));
ADDFHXL inst_cellmath__198_0_I2726 (.CO(N9911), .S(N10397), .A(N10516), .B(N10488), .CI(N10128));
ADDFXL inst_cellmath__198_0_I2727 (.CO(N10182), .S(N10050), .A(N3658), .B(N10226), .CI(N10237));
ADDFXL inst_cellmath__198_0_I2728 (.CO(N10456), .S(N10321), .A(N10423), .B(N9942), .CI(N10011));
ADDFXL inst_cellmath__198_0_I2729 (.CO(N10104), .S(N9971), .A(N9955), .B(N9982), .CI(N10419));
ADDFX1 inst_cellmath__198_0_I2730 (.CO(N10371), .S(N10238), .A(N10075), .B(N10050), .CI(N10321));
ADDFXL inst_cellmath__198_0_I2731 (.CO(N10029), .S(N10527), .A(N9971), .B(N10339), .CI(N9993));
ADDFXL inst_cellmath__198_0_I2732 (.CO(N10296), .S(N10161), .A(N10260), .B(N10238), .CI(N10527));
ADDFXL inst_cellmath__198_0_I2733 (.CO(N9946), .S(N10431), .A(N10511), .B(N10214), .CI(N10526));
ADDFX1 inst_cellmath__198_0_I2734 (.CO(N10218), .S(N10085), .A(N10276), .B(N10078), .CI(N10091));
ADDFX1 inst_cellmath__198_0_I2735 (.CO(N10500), .S(N10348), .A(N10456), .B(N10182), .CI(N10431));
ADDFHXL inst_cellmath__198_0_I2736 (.CO(N10136), .S(N10002), .A(N10104), .B(N10085), .CI(N10371));
ADDFHXL inst_cellmath__198_0_I2737 (.CO(N10408), .S(N10269), .A(N10029), .B(N10348), .CI(N10002));
ADDFX1 inst_cellmath__198_0_I2738 (.CO(N10059), .S(N9922), .A(N10362), .B(N10149), .CI(N10505));
ADDFX1 inst_cellmath__198_0_I2739 (.CO(N10328), .S(N10191), .A(N10224), .B(N10498), .CI(N9929));
ADDFX1 inst_cellmath__198_0_I2740 (.CO(N9980), .S(N10471), .A(N9946), .B(N10342), .CI(N9922));
ADDFHXL inst_cellmath__198_0_I2741 (.CO(N10245), .S(N10113), .A(N10218), .B(N10191), .CI(N10500));
ADDFXL inst_cellmath__198_0_I2742 (.CO(N10536), .S(N10383), .A(N10136), .B(N10471), .CI(N10113));
ADDFX1 inst_cellmath__198_0_I2743 (.CO(N10170), .S(N10038), .A(N10133), .B(N10140), .CI(N10356));
ADDFXL inst_cellmath__198_0_I2744 (.CO(N10442), .S(N10307), .A(N10198), .B(N9995), .CI(N10059));
ADDFXL inst_cellmath__198_0_I2745 (.CO(N10094), .S(N9959), .A(N10038), .B(N10328), .CI(N10307));
ADDFXL inst_cellmath__198_0_I2746 (.CO(N10358), .S(N10227), .A(N9980), .B(N10245), .CI(N9959));
ADDFX1 inst_cellmath__198_0_I2747 (.CO(N10014), .S(N10512), .A(N10528), .B(N10413), .CI(N10286));
ADDFX1 inst_cellmath__198_0_I2748 (.CO(N10281), .S(N10150), .A(N10509), .B(N10263), .CI(N10478));
ADDFXL inst_cellmath__198_0_I2749 (.CO(N9932), .S(N10418), .A(N10512), .B(N10170), .CI(N10442));
ADDFXL inst_cellmath__198_0_I2750 (.CO(N10202), .S(N10073), .A(N10418), .B(N10150), .CI(N10094));
ADDFX1 inst_cellmath__198_0_I2751 (.CO(N10484), .S(N10338), .A(N10066), .B(N9937), .CI(N9914));
ADDFX1 inst_cellmath__198_0_I2752 (.CO(N10125), .S(N9991), .A(N10014), .B(N10012), .CI(N10281));
ADDFX1 inst_cellmath__198_0_I2753 (.CO(N10395), .S(N10257), .A(N9932), .B(N10338), .CI(N9991));
ADDFX1 inst_cellmath__198_0_I2754 (.CO(N10046), .S(N9908), .A(N10334), .B(N10384), .CI(N10432));
ADDFX1 inst_cellmath__198_0_I2755 (.CO(N10318), .S(N10180), .A(N10147), .B(N10208), .CI(N10484));
ADDFX1 inst_cellmath__198_0_I2756 (.CO(N9969), .S(N10451), .A(N10125), .B(N9908), .CI(N10180));
ADDFX1 inst_cellmath__198_0_I2757 (.CO(N10234), .S(N10103), .A(N10086), .B(N10489), .CI(N10278));
ADDFX1 inst_cellmath__198_0_I2758 (.CO(N10525), .S(N10370), .A(N10103), .B(N10046), .CI(N10318));
ADDFX1 inst_cellmath__198_0_I2759 (.CO(N10159), .S(N10025), .A(N10349), .B(N9992), .CI(N10308));
ADDFX1 inst_cellmath__198_0_I2760 (.CO(N10427), .S(N10295), .A(N10234), .B(N10416), .CI(N10025));
ADDFX1 inst_cellmath__198_0_I2761 (.CO(N10083), .S(N9944), .A(N9930), .B(N9960), .CI(N10159));
ADDFX1 inst_cellmath__198_0_I2762 (.CO(N10346), .S(N10215), .A(N9909), .B(N9945), .CI(N10070));
OR2XL inst_cellmath__198_0_I2764 (.Y(N10134), .A(N9981), .B(N10336));
AND2XL inst_cellmath__198_0_I2765 (.Y(N10266), .A(N9981), .B(N10336));
NOR2XL inst_cellmath__198_0_I2766 (.Y(N10404), .A(N10481), .B(N9989));
NAND2XL inst_cellmath__198_0_I2767 (.Y(N9919), .A(N10481), .B(N9989));
OR2XL inst_cellmath__198_0_I2768 (.Y(N10058), .A(N10254), .B(N9906));
AND2XL inst_cellmath__198_0_I2769 (.Y(N10188), .A(N10254), .B(N9906));
NOR2XL inst_cellmath__198_0_I2770 (.Y(N10327), .A(N10043), .B(N10449));
NAND2XL inst_cellmath__198_0_I2771 (.Y(N10468), .A(N10043), .B(N10449));
OR2XL inst_cellmath__198_0_I2772 (.Y(N9978), .A(N10367), .B(N10022));
AND2XL inst_cellmath__198_0_I2773 (.Y(N10110), .A(N10367), .B(N10022));
NOR2XL inst_cellmath__198_0_I2774 (.Y(N10244), .A(N10157), .B(N10212));
NAND2XL inst_cellmath__198_0_I2775 (.Y(N10379), .A(N10157), .B(N10212));
OR2XL inst_cellmath__198_0_I2776 (.Y(N10534), .A(N10344), .B(N10056));
AND2XL inst_cellmath__198_0_I2777 (.Y(N10035), .A(N10344), .B(N10056));
NOR2XL inst_cellmath__198_0_I2778 (.Y(N10166), .A(N10187), .B(N10532));
NAND2XL inst_cellmath__198_0_I2779 (.Y(N10303), .A(N10187), .B(N10532));
NOR2XL inst_cellmath__198_0_I2780 (.Y(N10438), .A(N10034), .B(N10009));
NAND2X1 inst_cellmath__198_0_I2781 (.Y(N9952), .A(N10034), .B(N10009));
NOR4BX1 inst_cellmath__198_0_I10615 (.Y(N10354), .AN(inst_cellmath__61[2]), .B(N22574), .C(N22567), .D(N10506));
OAI21XL inst_cellmath__198_0_I2785 (.Y(N10480), .A0(N10266), .A1(N10354), .B0(N10134));
AOI21XL inst_cellmath__198_0_I2786 (.Y(N10314), .A0(N9919), .A1(N10480), .B0(N10404));
OAI21XL inst_cellmath__198_0_I2789 (.Y(N10079), .A0(N10188), .A1(N10314), .B0(N10058));
AOI21X1 inst_cellmath__198_0_I2790 (.Y(N10464), .A0(N10468), .A1(N10079), .B0(N10327));
OAI21X1 inst_cellmath__198_0_I2793 (.Y(N10142), .A0(N10110), .A1(N10464), .B0(N9978));
AOI21X1 inst_cellmath__198_0_I2794 (.Y(N10446), .A0(N10379), .A1(N10142), .B0(N10244));
OAI21X2 inst_cellmath__198_0_I2797 (.Y(N10051), .A0(N10035), .A1(N10446), .B0(N10534));
AOI21X1 inst_cellmath__198_0_I2798 (.Y(N9972), .A0(N10166), .A1(N9952), .B0(N10438));
INVX1 inst_cellmath__198_0_I2799 (.Y(N10123), .A(N9972));
CLKAND2X2 inst_cellmath__198_0_I2800 (.Y(N10255), .A(N10303), .B(N9952));
AOI21X2 inst_cellmath__198_0_I2802 (.Y(N10385), .A0(N10051), .A1(N10255), .B0(N10123));
INVX1 inst_cellmath__198_0_I2823 (.Y(N10169), .A(N10385));
NOR2XL inst_cellmath__198_0_I2824 (.Y(N10440), .A(N10143), .B(N10119));
NAND2X1 inst_cellmath__198_0_I2825 (.Y(N9957), .A(N10143), .B(N10119));
NOR2XL inst_cellmath__198_0_I2826 (.Y(N10092), .A(N10252), .B(N10519));
NOR2XL inst_cellmath__198_0_I2828 (.Y(N10357), .A(N10020), .B(N10261));
NAND2X1 inst_cellmath__198_0_I2829 (.Y(N10510), .A(N10020), .B(N10261));
NOR2X1 inst_cellmath__198_0_I2830 (.Y(N10013), .A(N10399), .B(N10299));
NAND2X1 inst_cellmath__198_0_I2831 (.Y(N10148), .A(N10399), .B(N10299));
NOR2XL inst_cellmath__198_0_I2832 (.Y(N10279), .A(N10434), .B(N9983));
NAND2X2 inst_cellmath__198_0_I2833 (.Y(N10417), .A(N10434), .B(N9983));
NOR2X1 inst_cellmath__198_0_I2834 (.Y(N9931), .A(N10115), .B(N10018));
NAND2X1 inst_cellmath__198_0_I2835 (.Y(N10071), .A(N10115), .B(N10018));
NOR2XL inst_cellmath__198_0_I2836 (.Y(N10201), .A(N10151), .B(N10397));
NAND2X2 inst_cellmath__198_0_I2837 (.Y(N10337), .A(N10151), .B(N10397));
NOR2XL inst_cellmath__198_0_I2840 (.Y(N10124), .A(N10296), .B(N10269));
NAND2X2 inst_cellmath__198_0_I2841 (.Y(N10256), .A(N10296), .B(N10269));
NOR2XL inst_cellmath__198_0_I2844 (.Y(N10044), .A(N10536), .B(N10227));
NAND2X1 inst_cellmath__198_0_I2845 (.Y(N10178), .A(N10536), .B(N10227));
NOR2X1 inst_cellmath__198_0_I2846 (.Y(N10317), .A(N10358), .B(N10073));
NAND2X1 inst_cellmath__198_0_I2847 (.Y(N10450), .A(N10358), .B(N10073));
NOR2XL inst_cellmath__198_0_I2848 (.Y(N9968), .A(N10202), .B(N10257));
NAND2X1 inst_cellmath__198_0_I2849 (.Y(N10101), .A(N10202), .B(N10257));
NOR2XL inst_cellmath__198_0_I2850 (.Y(N10233), .A(N10395), .B(N10451));
NAND2XL inst_cellmath__198_0_I2851 (.Y(N10369), .A(N10395), .B(N10451));
NOR2XL inst_cellmath__198_0_I2852 (.Y(N10524), .A(N9969), .B(N10370));
NAND2XL inst_cellmath__198_0_I2853 (.Y(N10023), .A(N9969), .B(N10370));
NOR2XL inst_cellmath__198_0_I2854 (.Y(N10158), .A(N10525), .B(N10295));
NAND2XL inst_cellmath__198_0_I2855 (.Y(N10293), .A(N10525), .B(N10295));
NOR2XL inst_cellmath__198_0_I2856 (.Y(N10426), .A(N9944), .B(N10427));
NAND2XL inst_cellmath__198_0_I2857 (.Y(N9943), .A(N9944), .B(N10427));
NOR2XL inst_cellmath__198_0_I2858 (.Y(N10082), .A(N10215), .B(N10083));
NAND2XL inst_cellmath__198_0_I2859 (.Y(N10213), .A(N10215), .B(N10083));
NOR2XL inst_cellmath__198_0_I2860 (.Y(N10345), .A(N10200), .B(N10346));
NAND2XL inst_cellmath__198_0_I2861 (.Y(N10497), .A(N10200), .B(N10346));
AOI21X2 inst_cellmath__198_0_I2862 (.Y(N9918), .A0(N9957), .A1(N10169), .B0(N10440));
AOI21X1 inst_cellmath__198_0_I2863 (.Y(N10467), .A0(N10510), .A1(N10092), .B0(N10357));
OAI2BB1X1 inst_cellmath__198_0_I10095 (.Y(N9977), .A0N(N10252), .A1N(N10519), .B0(N10510));
AOI21X2 inst_cellmath__198_0_I2865 (.Y(N10378), .A0(N10417), .A1(N10013), .B0(N10279));
NAND2X1 inst_cellmath__198_0_I2866 (.Y(N10533), .A(N10148), .B(N10417));
AOI21X2 inst_cellmath__198_0_I2867 (.Y(N10302), .A0(N10337), .A1(N9931), .B0(N10201));
NAND2X1 inst_cellmath__198_0_I2868 (.Y(N10437), .A(N10337), .B(N10071));
NOR2X1 inst_cellmath__203_0_I28082 (.Y(N10482), .A(N9911), .B(N10161));
AOI21X2 inst_cellmath__198_0_I2869 (.Y(N10222), .A0(N10482), .A1(N10256), .B0(N10124));
NAND2X1 inst_cellmath__203_0_I28083 (.Y(N9990), .A(N9911), .B(N10161));
NAND2X2 inst_cellmath__198_0_I2870 (.Y(N10352), .A(N10256), .B(N9990));
NOR2XL inst_cellmath__203_0_I28084 (.Y(N10394), .A(N10408), .B(N10383));
AOI21X1 inst_cellmath__198_0_I2871 (.Y(N10145), .A0(N10394), .A1(N10178), .B0(N10044));
NAND2X1 inst_cellmath__203_0_I28085 (.Y(N9907), .A(N10408), .B(N10383));
NAND2X2 inst_cellmath__198_0_I2872 (.Y(N10277), .A(N9907), .B(N10178));
AOI21X1 inst_cellmath__198_0_I2873 (.Y(N10069), .A0(N10101), .A1(N10317), .B0(N9968));
NAND2X1 inst_cellmath__198_0_I2874 (.Y(N10197), .A(N10101), .B(N10450));
INVXL inst_cellmath__198_0_I2875 (.Y(N10403), .A(N10233));
INVXL inst_cellmath__198_0_I2876 (.Y(N9917), .A(N10369));
AOI21XL inst_cellmath__198_0_I2877 (.Y(N9988), .A0(N10023), .A1(N10233), .B0(N10524));
NAND2XL inst_cellmath__198_0_I2878 (.Y(N10121), .A(N10023), .B(N10369));
OAI21XL inst_cellmath__198_0_I2879 (.Y(N10174), .A0(N9917), .A1(N10069), .B0(N10403));
NOR2XL inst_cellmath__198_0_I2880 (.Y(N10313), .A(N9917), .B(N10197));
AOI21XL inst_cellmath__198_0_I2881 (.Y(N10364), .A0(N9943), .A1(N10158), .B0(N10426));
NAND2XL inst_cellmath__198_0_I2882 (.Y(N10520), .A(N9943), .B(N10293));
INVXL inst_cellmath__198_0_I2883 (.Y(N10243), .A(N10082));
INVXL inst_cellmath__198_0_I2884 (.Y(N10377), .A(N10213));
AOI21XL inst_cellmath__198_0_I2885 (.Y(N10289), .A0(N10497), .A1(N10082), .B0(N10345));
NAND2XL inst_cellmath__198_0_I2886 (.Y(N10424), .A(N10497), .B(N10213));
OAI21XL inst_cellmath__198_0_I2887 (.Y(N10492), .A0(N10377), .A1(N10364), .B0(N10243));
NOR2XL inst_cellmath__198_0_I2888 (.Y(N9996), .A(N10377), .B(N10520));
OA21X1 inst_cellmath__198_0_I2889 (.Y(N10010), .A0(N10121), .A1(N10069), .B0(N9988));
OR2XL inst_cellmath__198_0_I2890 (.Y(N10144), .A(N10121), .B(N10197));
OA21X1 inst_cellmath__198_0_I2891 (.Y(N10479), .A0(N10424), .A1(N10364), .B0(N10289));
OR2XL inst_cellmath__198_0_I2892 (.Y(N9987), .A(N10424), .B(N10520));
INVXL inst_cellmath__198_0_I2893 (.Y(N10120), .A(N9918));
OAI21X1 inst_cellmath__198_0_I2895 (.Y(N10273), .A0(N10533), .A1(N10467), .B0(N10378));
NOR2XL inst_cellmath__198_0_I2896 (.Y(N10412), .A(N9977), .B(N10533));
OAI21X1 inst_cellmath__198_0_I2899 (.Y(N10194), .A0(N10352), .A1(N10302), .B0(N10222));
NOR2XL inst_cellmath__198_0_I2900 (.Y(N10333), .A(N10352), .B(N10437));
OAI21X2 inst_cellmath__198_0_I2901 (.Y(N10475), .A0(N10277), .A1(N10222), .B0(N10145));
NOR2X1 inst_cellmath__198_0_I2902 (.Y(N9985), .A(N10277), .B(N10352));
OAI21XL inst_cellmath__198_0_I2903 (.Y(N10117), .A0(N10144), .A1(N10145), .B0(N10010));
NOR2X1 inst_cellmath__198_0_I2904 (.Y(N10249), .A(N10144), .B(N10277));
OAI21XL inst_cellmath__198_0_I2905 (.Y(N10387), .A0(N9987), .A1(N10010), .B0(N10479));
NOR2XL inst_cellmath__198_0_I2906 (.Y(N10539), .A(N9987), .B(N10144));
OAI21X1 inst_cellmath__203_0_I28086 (.Y(N10006), .A0(N9977), .A1(N9918), .B0(N10467));
INVXL inst_cellmath__198_0_I2908 (.Y(N10390), .A(N10006));
AOI21X1 inst_cellmath__198_0_I2909 (.Y(N9962), .A0(N10412), .A1(N10120), .B0(N10273));
OAI21X1 inst_cellmath__203_0_I28087 (.Y(N9925), .A0(N10437), .A1(N10378), .B0(N10302));
AOI21X1 inst_cellmath__198_0_I2913 (.Y(N10152), .A0(N9985), .A1(N9925), .B0(N10475));
NOR2XL inst_cellmath__203_0_I28088 (.Y(N10065), .A(N10533), .B(N10437));
NAND2X1 inst_cellmath__198_0_I2914 (.Y(N10285), .A(N9985), .B(N10065));
AOI21XL inst_cellmath__198_0_I2915 (.Y(N10420), .A0(N10249), .A1(N10194), .B0(N10117));
NAND2XL inst_cellmath__198_0_I2916 (.Y(N9936), .A(N10249), .B(N10333));
AOI21XL inst_cellmath__198_0_I2917 (.Y(N10076), .A0(N10539), .A1(N10475), .B0(N10387));
NAND2XL inst_cellmath__198_0_I2918 (.Y(N10207), .A(N10539), .B(N9985));
OAI21X2 inst_cellmath__198_0_I2920 (.Y(N10457), .A0(N10285), .A1(N10390), .B0(N10152));
OAI21X2 inst_cellmath__198_0_I2921 (.Y(N10105), .A0(N9936), .A1(N9962), .B0(N10420));
AOI21X1 inst_cellmath__203_0_I28090 (.Y(N10229), .A0(N10006), .A1(N10065), .B0(N9925));
OAI21XL inst_cellmath__198_0_I2922 (.Y(N10372), .A0(N10207), .A1(N10229), .B0(N10076));
INVXL inst_cellmath__198_0_I2923 (.Y(N10210), .A(N10069));
INVXL inst_cellmath__198_0_I2924 (.Y(N10400), .A(N10364));
NAND2BXL inst_cellmath__198_0_I2929 (.Y(N10258), .AN(N10279), .B(N10417));
NAND2BXL inst_cellmath__198_0_I2930 (.Y(N10047), .AN(N9931), .B(N10071));
NAND2BXL inst_cellmath__198_0_I2931 (.Y(N10452), .AN(N10201), .B(N10337));
NAND2BXL inst_cellmath__198_0_I2932 (.Y(N10235), .AN(N10482), .B(N9990));
NAND2BXL inst_cellmath__198_0_I2935 (.Y(N10216), .AN(N10044), .B(N10178));
NAND2BXL inst_cellmath__198_0_I2936 (.Y(N10000), .AN(N10317), .B(N10450));
NAND2BXL inst_cellmath__198_0_I2937 (.Y(N10405), .AN(N9968), .B(N10101));
NAND2BXL inst_cellmath__198_0_I2938 (.Y(N10190), .AN(N10233), .B(N10369));
NAND2BXL inst_cellmath__198_0_I2939 (.Y(N9979), .AN(N10524), .B(N10023));
NAND2BXL inst_cellmath__198_0_I2940 (.Y(N10381), .AN(N10158), .B(N10293));
NAND2BXL inst_cellmath__198_0_I2941 (.Y(N10167), .AN(N10426), .B(N9943));
NAND2BXL inst_cellmath__198_0_I2942 (.Y(N9954), .AN(N10082), .B(N10213));
NAND2BXL inst_cellmath__198_0_I2943 (.Y(N10355), .AN(N10345), .B(N10497));
NOR2BX1 inst_cellmath__198_0_I2944 (.Y(N10146), .AN(N10204), .B(N10486));
XNOR2X1 inst_cellmath__198_0_I2948 (.Y(inst_cellmath__198[18]), .A(N9962), .B(N10047));
XNOR2XL inst_cellmath__198_0_I2949 (.Y(inst_cellmath__198[20]), .A(N10229), .B(N10235));
XNOR2XL inst_cellmath__198_0_I2952 (.Y(inst_cellmath__198[28]), .A(N10381), .B(N10105));
XOR2XL inst_cellmath__198_0_I2953 (.Y(inst_cellmath__198[32]), .A(N10372), .B(N10146));
XNOR2XL inst_cellmath__198_0_I2957 (.Y(N10176), .A(N10258), .B(N10148));
XNOR2XL inst_cellmath__198_0_I2958 (.Y(N10315), .A(N10258), .B(N10013));
XNOR2X1 inst_cellmath__198_0_I2960 (.Y(N9966), .A(N10071), .B(N10452));
XNOR2X1 inst_cellmath__198_0_I2961 (.Y(N10099), .A(N9931), .B(N10452));
MXI2X1 inst_cellmath__198_0_I2962 (.Y(inst_cellmath__198[19]), .A(N9966), .B(N10099), .S0(N9962));
XNOR2X1 inst_cellmath__198_0_I2966 (.Y(N10156), .A(N10216), .B(N9907));
XNOR2X1 inst_cellmath__198_0_I2967 (.Y(N10291), .A(N10394), .B(N10216));
XNOR2X1 inst_cellmath__198_0_I2969 (.Y(N9940), .A(N10405), .B(N10450));
XNOR2X1 inst_cellmath__198_0_I2970 (.Y(N10080), .A(N10405), .B(N10317));
MX2X1 inst_cellmath__198_0_I2971 (.Y(inst_cellmath__198[25]), .A(N10080), .B(N9940), .S0(N10457));
XNOR2X1 inst_cellmath__198_0_I2972 (.Y(N10343), .A(N10190), .B(N10210));
NOR2BX1 inst_cellmath__198_0_I2973 (.Y(N10199), .AN(N10197), .B(N10210));
XOR2XL inst_cellmath__198_0_I2974 (.Y(N10495), .A(N10190), .B(N10199));
MX2XL inst_cellmath__198_0_I2975 (.Y(inst_cellmath__198[26]), .A(N10343), .B(N10495), .S0(N10457));
XNOR2X1 inst_cellmath__198_0_I2976 (.Y(N10131), .A(N9979), .B(N10174));
NOR2XL inst_cellmath__198_0_I2977 (.Y(N10175), .A(N10313), .B(N10174));
XOR2XL inst_cellmath__198_0_I2978 (.Y(N10264), .A(N9979), .B(N10175));
MX2XL inst_cellmath__198_0_I2979 (.Y(inst_cellmath__198[27]), .A(N10131), .B(N10264), .S0(N10457));
XNOR2X1 inst_cellmath__198_0_I2980 (.Y(N9915), .A(N10167), .B(N10293));
XNOR2X1 inst_cellmath__198_0_I2981 (.Y(N10055), .A(N10167), .B(N10158));
MXI2XL inst_cellmath__198_0_I2982 (.Y(inst_cellmath__198[29]), .A(N10055), .B(N9915), .S0(N10105));
XNOR2X1 inst_cellmath__198_0_I2983 (.Y(N10325), .A(N9954), .B(N10400));
NOR2BX1 inst_cellmath__198_0_I2984 (.Y(N10493), .AN(N10520), .B(N10400));
XOR2XL inst_cellmath__198_0_I2985 (.Y(N10465), .A(N9954), .B(N10493));
MXI2XL inst_cellmath__198_0_I2986 (.Y(inst_cellmath__198[30]), .A(N10325), .B(N10465), .S0(N10105));
XNOR2X1 inst_cellmath__198_0_I2987 (.Y(N10108), .A(N10355), .B(N10492));
NOR2XL inst_cellmath__198_0_I2988 (.Y(N10463), .A(N9996), .B(N10492));
XOR2XL inst_cellmath__198_0_I2989 (.Y(N10241), .A(N10355), .B(N10463));
MXI2XL inst_cellmath__198_0_I2990 (.Y(inst_cellmath__198[31]), .A(N10108), .B(N10241), .S0(N10105));
NOR4BBX1 inst_cellmath__203_0_I10096 (.Y(N11288), .AN(N7933), .BN(N8335), .C(N7685), .D(N7749));
NOR4BX1 inst_cellmath__203_0_I10222 (.Y(N12219), .AN(N8076), .B(N8562), .C(N7979), .D(N8533));
NAND4XL hyperpropagate_4_1_A_I28289 (.Y(N22651), .A(N8164), .B(N8440), .C(N7780), .D(N7810));
NOR2XL hyperpropagate_4_1_A_I10772 (.Y(N12579), .A(N7958), .B(N22651));
NOR4BX1 inst_cellmath__203_0_I10223 (.Y(N11223), .AN(N7783), .B(N7777), .C(N8519), .D(N8584));
NAND3XL hyperpropagate_4_1_A_I10773 (.Y(N22659), .A(N8735), .B(N7849), .C(N7715));
NOR2X1 hyperpropagate_4_1_A_I10774 (.Y(N11600), .A(N22659), .B(N8494));
INVX1 inst_cellmath__203_0_I2996 (.Y(N11999), .A(inst_cellmath__197[5]));
INVX1 inst_cellmath__203_0_I2997 (.Y(N12373), .A(inst_cellmath__197[6]));
NOR4BBX1 inst_cellmath__203_0_I10225 (.Y(N12720), .AN(N8133), .BN(N8237), .C(N8550), .D(N7844));
INVXL inst_cellmath__203_0_I2999 (.Y(N11377), .A(inst_cellmath__197[8]));
NOR4BBX1 inst_cellmath__203_0_I10226 (.Y(N11761), .AN(N8437), .BN(N8058), .C(N7787), .D(N8416));
NOR4BBX1 inst_cellmath__203_0_I10227 (.Y(N12154), .AN(N8167), .BN(N7782), .C(N8649), .D(N8275));
NAND3XL hyperpropagate_4_1_A_I28624 (.Y(N44079), .A(N8055), .B(N8323), .C(N8012));
NOR2XL hyperpropagate_4_1_A_I28625 (.Y(N12523), .A(N8143), .B(N44079));
NAND3XL hyperpropagate_4_1_A_I28626 (.Y(N44087), .A(N7894), .B(N8160), .C(N8706));
NOR2XL hyperpropagate_4_1_A_I28627 (.Y(N12874), .A(N8655), .B(N44087));
NAND3XL hyperpropagate_4_1_A_I28628 (.Y(N44095), .A(N7966), .B(N8782), .C(N8102));
NOR2XL hyperpropagate_4_1_A_I28629 (.Y(N11540), .A(N8681), .B(N44095));
NOR2XL inst_cellmath__203_0_I10107 (.Y(N11930), .A(N8001), .B(N8235));
NAND3XL hyperpropagate_4_1_A_I28630 (.Y(N44103), .A(N8363), .B(N8215), .C(N7887));
NOR2XL hyperpropagate_4_1_A_I28631 (.Y(N12313), .A(N8212), .B(N44103));
INVX1 inst_cellmath__203_0_I3007 (.Y(N12667), .A(inst_cellmath__197[16]));
NAND3XL hyperpropagate_4_1_A_I10783 (.Y(N22699), .A(N8684), .B(N8304), .C(N8165));
NOR2X1 hyperpropagate_4_1_A_I10784 (.Y(N11318), .A(N8556), .B(N22699));
NAND2XL hyperpropagate_3_1_A_I10785 (.Y(N22705), .A(N8141), .B(N7910));
NOR2X1 hyperpropagate_3_1_A_I10786 (.Y(N11691), .A(N22705), .B(N8608));
NAND3XL hyperpropagate_4_1_A_I10787 (.Y(N22714), .A(N8316), .B(N8512), .C(N8018));
NOR2X1 hyperpropagate_4_1_A_I10788 (.Y(N12093), .A(N8652), .B(N22714));
CLKMX2X2 inst_cellmath__203_0_I10112 (.Y(N11631), .A(N10176), .B(N10315), .S0(N10390));
NOR2XL inst_cellmath__203_0_I3017 (.Y(N12835), .A(N11631), .B(N12219));
NOR2XL inst_cellmath__203_0_I3018 (.Y(N11889), .A(N11631), .B(N12579));
NOR2XL inst_cellmath__203_0_I3019 (.Y(N12628), .A(N11631), .B(N11223));
NOR2XL inst_cellmath__203_0_I3020 (.Y(N11653), .A(N11631), .B(N11600));
NOR2XL inst_cellmath__203_0_I3021 (.Y(N12422), .A(N11631), .B(N11999));
NOR2XL inst_cellmath__203_0_I3022 (.Y(N11435), .A(N11631), .B(N12373));
NOR2XL inst_cellmath__203_0_I3023 (.Y(N12208), .A(N11631), .B(N12720));
NOR2XL inst_cellmath__203_0_I3024 (.Y(N11209), .A(N11631), .B(N11377));
NOR2X1 inst_cellmath__203_0_I3025 (.Y(N11986), .A(N11761), .B(N11631));
NOR2XL inst_cellmath__203_0_I3026 (.Y(N12709), .A(N11631), .B(N12154));
NOR2XL inst_cellmath__203_0_I3027 (.Y(N11749), .A(N11631), .B(N12523));
NOR2XL inst_cellmath__203_0_I3028 (.Y(N12509), .A(N11631), .B(N12874));
NOR2XL inst_cellmath__203_0_I3029 (.Y(N11528), .A(N11631), .B(N11540));
NOR2XL inst_cellmath__203_0_I3030 (.Y(N12301), .A(N11631), .B(N11930));
NOR2XL inst_cellmath__203_0_I3031 (.Y(N11305), .A(N11631), .B(N12313));
NOR2XL inst_cellmath__203_0_I3032 (.Y(N12081), .A(N11631), .B(N12667));
NOR2X1 inst_cellmath__203_0_I3033 (.Y(N12800), .A(N11318), .B(N11631));
NOR2XL inst_cellmath__203_0_I3034 (.Y(N11853), .A(N11631), .B(N11691));
NOR2XL inst_cellmath__203_0_I3035 (.Y(N12595), .A(N11631), .B(N12093));
INVX2 inst_cellmath__203_0_I3037 (.Y(N11183), .A(inst_cellmath__198[18]));
NAND2BX2 inst_cellmath__203_0_I10113 (.Y(N12488), .AN(inst_cellmath__198[19]), .B(inst_cellmath__198[18]));
INVXL inst_cellmath__203_0_I3040 (.Y(N12839), .A(inst_cellmath__198[19]));
NOR2XL inst_cellmath__203_0_I3041 (.Y(N12032), .A(N11288), .B(N11183));
MXI2XL inst_cellmath__203_0_I3042 (.Y(inst_cellmath__203__W0[1]), .A(N12839), .B(N12488), .S0(N12032));
MXI2XL inst_cellmath__203_0_I3043 (.Y(N11965), .A(N12219), .B(N11288), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3044 (.Y(N11504), .A(N12839), .B(N12488), .S0(N11965));
MXI2XL inst_cellmath__203_0_I3046 (.Y(N11899), .A(N12579), .B(N12219), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3047 (.Y(N12324), .A(N12839), .B(N12488), .S0(N11899));
MXI2XL inst_cellmath__203_0_I3048 (.Y(N11829), .A(N11223), .B(N12579), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3049 (.Y(N12680), .A(N12839), .B(N12488), .S0(N11829));
MXI2XL inst_cellmath__203_0_I3050 (.Y(N11760), .A(N11600), .B(N11223), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3051 (.Y(N11332), .A(N12839), .B(N12488), .S0(N11760));
MXI2XL inst_cellmath__203_0_I3052 (.Y(N11690), .A(N11999), .B(N11600), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3053 (.Y(N11711), .A(N12839), .B(N12488), .S0(N11690));
MXI2XL inst_cellmath__203_0_I3054 (.Y(N11630), .A(N12373), .B(N11999), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3055 (.Y(N12109), .A(N12839), .B(N12488), .S0(N11630));
MXI2XL inst_cellmath__203_0_I3056 (.Y(N11565), .A(N12720), .B(N12373), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3057 (.Y(N12473), .A(N12839), .B(N12488), .S0(N11565));
MXI2XL inst_cellmath__203_0_I3058 (.Y(N11503), .A(N11377), .B(N12720), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3059 (.Y(N12826), .A(N12839), .B(N12488), .S0(N11503));
MXI2XL inst_cellmath__203_0_I3060 (.Y(N11437), .A(N11761), .B(N11377), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3061 (.Y(N11494), .A(N12839), .B(N12488), .S0(N11437));
MXI2XL inst_cellmath__203_0_I3062 (.Y(N11365), .A(N12154), .B(N11761), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3063 (.Y(N11879), .A(N12839), .B(N12488), .S0(N11365));
MXI2XL inst_cellmath__203_0_I3064 (.Y(N11308), .A(N12523), .B(N12154), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3065 (.Y(N12263), .A(N12839), .B(N12488), .S0(N11308));
MXI2XL inst_cellmath__203_0_I3066 (.Y(N11241), .A(N12874), .B(N12523), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3067 (.Y(N12621), .A(N12839), .B(N12488), .S0(N11241));
MXI2XL inst_cellmath__203_0_I3068 (.Y(N11175), .A(N11540), .B(N12874), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3069 (.Y(N11267), .A(N12839), .B(N12488), .S0(N11175));
MXI2XL inst_cellmath__203_0_I3070 (.Y(N12828), .A(N11930), .B(N11540), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3071 (.Y(N11648), .A(N12839), .B(N12488), .S0(N12828));
MXI2XL inst_cellmath__203_0_I3072 (.Y(N12767), .A(N12313), .B(N11930), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3073 (.Y(N12045), .A(N12839), .B(N12488), .S0(N12767));
MXI2XL inst_cellmath__203_0_I3074 (.Y(N12704), .A(N12667), .B(N12313), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3075 (.Y(N12414), .A(N12839), .B(N12488), .S0(N12704));
MXI2XL inst_cellmath__203_0_I3076 (.Y(N12652), .A(N11318), .B(N12667), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3077 (.Y(N12764), .A(N12839), .B(N12488), .S0(N12652));
MXI2XL inst_cellmath__203_0_I3078 (.Y(N12590), .A(N11691), .B(N11318), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3079 (.Y(N11429), .A(N12839), .B(N12488), .S0(N12590));
MXI2XL inst_cellmath__203_0_I3080 (.Y(N12532), .A(N12093), .B(N11691), .S0(N11183));
MXI2XL inst_cellmath__203_0_I3081 (.Y(N11811), .A(N12839), .B(N12488), .S0(N12532));
NAND2XL inst_cellmath__203_0_I3082 (.Y(N12468), .A(N12093), .B(N11183));
MXI2XL inst_cellmath__203_0_I3083 (.Y(N12200), .A(N12839), .B(N12488), .S0(N12468));
XOR2XL inst_cellmath__203_0_I3084 (.Y(N11979), .A(inst_cellmath__198[20]), .B(inst_cellmath__198[19]));
INVXL inst_cellmath__203_0_I28099 (.Y(N43769), .A(N10482));
NAND2BXL inst_cellmath__203_0_I28094 (.Y(N43761), .AN(N10124), .B(N10256));
XOR2XL inst_cellmath__203_0_I28296 (.Y(N43755), .A(N43769), .B(N43761));
XNOR2X1 inst_cellmath__203_0_I28097 (.Y(N43747), .A(N9990), .B(N43761));
INVXL inst_cellmath__203_0_I28101 (.Y(N43739), .A(N10229));
MX2X1 inst_cellmath__203_0_I28102 (.Y(inst_cellmath__198[21]), .A(N43755), .B(N43747), .S0(N43739));
AOI21XL inst_cellmath__203_0_I10530 (.Y(N12702), .A0(inst_cellmath__198[20]), .A1(inst_cellmath__198[19]), .B0(inst_cellmath__198[21]));
OA21X1 inst_cellmath__203_0_I10531 (.Y(N12350), .A0(inst_cellmath__198[20]), .A1(inst_cellmath__198[19]), .B0(inst_cellmath__198[21]));
INVX2 inst_cellmath__203_0_I3090 (.Y(N12426), .A(N11979));
INVX3 inst_cellmath__203_0_I9955 (.Y(N22577), .A(N12426));
INVX2 inst_cellmath__203_0_I9959 (.Y(N22581), .A(N22577));
INVX2 inst_cellmath__203_0_I9958 (.Y(N22580), .A(N22577));
INVX1 inst_cellmath__203_0_I9957 (.Y(N22579), .A(N22577));
INVX1 inst_cellmath__203_0_I9956 (.Y(N22578), .A(N22577));
INVX1 inst_cellmath__203_0_I3095 (.Y(N11990), .A(N12350));
INVX1 inst_cellmath__203_0_I3097 (.Y(N12362), .A(N12702));
NOR2XL inst_cellmath__203_0_I3098 (.Y(N12129), .A(N11288), .B(N22580));
MXI2XL inst_cellmath__203_0_I3099 (.Y(N12504), .A(N12362), .B(N11990), .S0(N12129));
MXI2XL inst_cellmath__203_0_I3100 (.Y(N12067), .A(N12219), .B(N11288), .S0(N22581));
MXI2XL inst_cellmath__203_0_I3101 (.Y(N12856), .A(N12362), .B(N11990), .S0(N12067));
MXI2XL inst_cellmath__203_0_I3102 (.Y(N12003), .A(N12579), .B(N12219), .S0(N22578));
MXI2XL inst_cellmath__203_0_I3103 (.Y(N11522), .A(N12362), .B(N11990), .S0(N12003));
MXI2XL inst_cellmath__203_0_I3104 (.Y(N11933), .A(N11223), .B(N12579), .S0(N22578));
MXI2X1 inst_cellmath__203_0_I3105 (.Y(N11911), .A(N12362), .B(N11990), .S0(N11933));
MXI2XL inst_cellmath__203_0_I3106 (.Y(N11864), .A(N11600), .B(N11223), .S0(N12426));
MXI2XL inst_cellmath__203_0_I3107 (.Y(N12290), .A(N12362), .B(N11990), .S0(N11864));
MXI2XL inst_cellmath__203_0_I3108 (.Y(N11794), .A(N11999), .B(N11600), .S0(N22578));
MXI2XL inst_cellmath__203_0_I3109 (.Y(N12649), .A(N12362), .B(N11990), .S0(N11794));
MXI2XL inst_cellmath__203_0_I3110 (.Y(N11724), .A(N12373), .B(N11999), .S0(N22578));
MXI2XL inst_cellmath__203_0_I3111 (.Y(N11299), .A(N12362), .B(N11990), .S0(N11724));
MXI2XL inst_cellmath__203_0_I3112 (.Y(N11658), .A(N12720), .B(N12373), .S0(N22578));
MXI2X1 inst_cellmath__203_0_I3113 (.Y(N11673), .A(N12362), .B(N11990), .S0(N11658));
MXI2XL inst_cellmath__203_0_I3114 (.Y(N11594), .A(N11377), .B(N12720), .S0(N12426));
MXI2XL inst_cellmath__203_0_I3115 (.Y(N12073), .A(N12362), .B(N11990), .S0(N11594));
MXI2XL inst_cellmath__203_0_I3116 (.Y(N11534), .A(N11761), .B(N11377), .S0(N22579));
MXI2XL inst_cellmath__203_0_I3117 (.Y(N12442), .A(N12362), .B(N11990), .S0(N11534));
MXI2XL inst_cellmath__203_0_I3118 (.Y(N11471), .A(N12154), .B(N11761), .S0(N22579));
MXI2XL inst_cellmath__203_0_I3119 (.Y(N12793), .A(N12362), .B(N11990), .S0(N11471));
MXI2XL inst_cellmath__203_0_I3120 (.Y(N11400), .A(N12523), .B(N12154), .S0(N22579));
MXI2XL inst_cellmath__203_0_I3121 (.Y(N11458), .A(N12362), .B(N11990), .S0(N11400));
MXI2XL inst_cellmath__203_0_I3122 (.Y(N11338), .A(N12874), .B(N12523), .S0(N22579));
MXI2XL inst_cellmath__203_0_I3123 (.Y(N11845), .A(N12362), .B(N11990), .S0(N11338));
MXI2XL inst_cellmath__203_0_I3124 (.Y(N11274), .A(N11540), .B(N12874), .S0(N22579));
MXI2XL inst_cellmath__203_0_I3125 (.Y(N12230), .A(N12362), .B(N11990), .S0(N11274));
MXI2XL inst_cellmath__203_0_I3126 (.Y(N11206), .A(N11930), .B(N11540), .S0(N22580));
MXI2XL inst_cellmath__203_0_I3127 (.Y(N12587), .A(N12362), .B(N11990), .S0(N11206));
MXI2XL inst_cellmath__203_0_I3128 (.Y(N12863), .A(N12313), .B(N11930), .S0(N22580));
MXI2XL inst_cellmath__203_0_I3129 (.Y(N11234), .A(N12362), .B(N11990), .S0(N12863));
MXI2X1 inst_cellmath__203_0_I3130 (.Y(N12801), .A(N12667), .B(N12313), .S0(N22580));
MXI2X1 inst_cellmath__203_0_I3131 (.Y(N11614), .A(N12362), .B(N11990), .S0(N12801));
MXI2X1 inst_cellmath__203_0_I3132 (.Y(N12739), .A(N11318), .B(N12667), .S0(N22580));
MXI2X1 inst_cellmath__203_0_I3133 (.Y(N12009), .A(N12362), .B(N11990), .S0(N12739));
MXI2XL inst_cellmath__203_0_I3134 (.Y(N12681), .A(N11691), .B(N11318), .S0(N12426));
MXI2XL inst_cellmath__203_0_I3135 (.Y(N12382), .A(N12362), .B(N11990), .S0(N12681));
MXI2X1 inst_cellmath__203_0_I3136 (.Y(N12622), .A(N12093), .B(N11691), .S0(N22581));
MXI2X1 inst_cellmath__203_0_I3137 (.Y(N12731), .A(N12362), .B(N11990), .S0(N12622));
NAND2X1 inst_cellmath__203_0_I3138 (.Y(N12562), .A(N12093), .B(N22581));
MXI2X1 inst_cellmath__203_0_I3139 (.Y(N11387), .A(N12362), .B(N11990), .S0(N12562));
NAND2BXL inst_cellmath__203_0_I28095 (.Y(N43770), .AN(N10394), .B(N9907));
NAND2XL inst_cellmath__203_0_I28092 (.Y(N43743), .A(N10412), .B(N10333));
INVXL inst_cellmath__203_0_I28089 (.Y(N43757), .A(N10120));
AOI21X1 inst_cellmath__203_0_I28091 (.Y(N43775), .A0(N10333), .A1(N10273), .B0(N10194));
OAI21X1 inst_cellmath__203_0_I28093 (.Y(N10183), .A0(N43757), .A1(N43743), .B0(N43775));
XNOR2XL inst_cellmath__203_0_I28096 (.Y(inst_cellmath__198[22]), .A(N10183), .B(N43770));
NOR2XL inst_cellmath__203_0_I3140 (.Y(N12505), .A(inst_cellmath__198[21]), .B(inst_cellmath__198[22]));
NAND2XL inst_cellmath__203_0_I3141 (.Y(N11523), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
MX2XL inst_cellmath__203_0_I27945 (.Y(inst_cellmath__198[23]), .A(N10291), .B(N10156), .S0(N10183));
NOR2XL inst_cellmath__203_0_I3142 (.Y(N11938), .A(N12505), .B(inst_cellmath__198[23]));
CLKXOR2X1 inst_cellmath__203_0_I28103 (.Y(N12713), .A(inst_cellmath__198[21]), .B(inst_cellmath__198[22]));
INVX2 inst_cellmath__203_0_I3144 (.Y(N12514), .A(N12713));
CLKINVX4 inst_cellmath__203_0_I9960 (.Y(N22582), .A(N12514));
CLKINVX12 inst_cellmath__203_0_I9961 (.Y(N22583), .A(N22582));
NAND2X2 inst_cellmath__203_0_I3148 (.Y(N12451), .A(N11523), .B(inst_cellmath__198[23]));
INVX1 inst_cellmath__203_0_I3149 (.Y(N12804), .A(N11938));
NOR2XL inst_cellmath__203_0_I3150 (.Y(N12227), .A(N11288), .B(N22583));
MXI2X1 inst_cellmath__203_0_I3151 (.Y(N11701), .A(N12804), .B(N12451), .S0(N12227));
MXI2XL inst_cellmath__203_0_I3152 (.Y(N12163), .A(N11288), .B(N12219), .S0(N12713));
MXI2XL inst_cellmath__203_0_I3153 (.Y(N12101), .A(N12804), .B(N12451), .S0(N12163));
MXI2XL inst_cellmath__203_0_I3154 (.Y(N12102), .A(N12579), .B(N12219), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3155 (.Y(N12465), .A(N12804), .B(N12451), .S0(N12102));
MXI2XL inst_cellmath__203_0_I3156 (.Y(N12037), .A(N11223), .B(N12579), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3157 (.Y(N12820), .A(N12804), .B(N12451), .S0(N12037));
MXI2XL inst_cellmath__203_0_I3158 (.Y(N11970), .A(N11600), .B(N11223), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3159 (.Y(N11486), .A(N12804), .B(N12451), .S0(N11970));
MXI2XL inst_cellmath__203_0_I3160 (.Y(N11902), .A(N11999), .B(N11600), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3161 (.Y(N11869), .A(N12804), .B(N12451), .S0(N11902));
MXI2XL inst_cellmath__203_0_I3162 (.Y(N11835), .A(N12373), .B(N11999), .S0(N12514));
MXI2XL inst_cellmath__203_0_I3163 (.Y(N12255), .A(N12804), .B(N12451), .S0(N11835));
MXI2XL inst_cellmath__203_0_I3164 (.Y(N11764), .A(N12720), .B(N12373), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3165 (.Y(N12615), .A(N12804), .B(N12451), .S0(N11764));
MXI2XL inst_cellmath__203_0_I3166 (.Y(N11694), .A(N11377), .B(N12720), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3167 (.Y(N11260), .A(N12804), .B(N12451), .S0(N11694));
MXI2XL inst_cellmath__203_0_I3168 (.Y(N11633), .A(N11761), .B(N11377), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3169 (.Y(N11639), .A(N12804), .B(N12451), .S0(N11633));
MXI2XL inst_cellmath__203_0_I3170 (.Y(N11567), .A(N12154), .B(N11761), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3171 (.Y(N12036), .A(N12804), .B(N12451), .S0(N11567));
MXI2XL inst_cellmath__203_0_I3172 (.Y(N11505), .A(N12523), .B(N12154), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3173 (.Y(N12406), .A(N12804), .B(N12451), .S0(N11505));
MXI2XL inst_cellmath__203_0_I3174 (.Y(N11440), .A(N12874), .B(N12523), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3175 (.Y(N12757), .A(N12804), .B(N12451), .S0(N11440));
MXI2XL inst_cellmath__203_0_I3176 (.Y(N11369), .A(N11540), .B(N12874), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3177 (.Y(N11419), .A(N12804), .B(N12451), .S0(N11369));
MXI2XL inst_cellmath__203_0_I3178 (.Y(N11311), .A(N11930), .B(N11540), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3179 (.Y(N11801), .A(N12804), .B(N12451), .S0(N11311));
MXI2XL inst_cellmath__203_0_I3180 (.Y(N11245), .A(N12313), .B(N11930), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3181 (.Y(N12191), .A(N12804), .B(N12451), .S0(N11245));
MXI2X1 inst_cellmath__203_0_I3182 (.Y(N11179), .A(N12667), .B(N12313), .S0(N22583));
MXI2X1 inst_cellmath__203_0_I3183 (.Y(N12557), .A(N12804), .B(N12451), .S0(N11179));
MXI2XL inst_cellmath__203_0_I3184 (.Y(N12832), .A(N11318), .B(N12667), .S0(N12514));
MXI2XL inst_cellmath__203_0_I3185 (.Y(N11193), .A(N12804), .B(N12451), .S0(N12832));
MXI2XL inst_cellmath__203_0_I3186 (.Y(N12771), .A(N11691), .B(N11318), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3187 (.Y(N11576), .A(N12804), .B(N12451), .S0(N12771));
MXI2XL inst_cellmath__203_0_I3188 (.Y(N12707), .A(N12093), .B(N11691), .S0(N22583));
MXI2XL inst_cellmath__203_0_I3189 (.Y(N11969), .A(N12804), .B(N12451), .S0(N12707));
NAND2XL inst_cellmath__203_0_I3190 (.Y(N12655), .A(N12093), .B(N22583));
MXI2XL inst_cellmath__203_0_I3191 (.Y(N12344), .A(N12804), .B(N12451), .S0(N12655));
XNOR2XL inst_cellmath__203_0_I27944 (.Y(inst_cellmath__198[24]), .A(N10000), .B(N10457));
NOR2XL inst_cellmath__203_0_I3193 (.Y(N12593), .A(inst_cellmath__198[23]), .B(inst_cellmath__198[24]));
NAND2XL inst_cellmath__203_0_I3194 (.Y(N11620), .A(inst_cellmath__198[24]), .B(inst_cellmath__198[23]));
NOR2XL inst_cellmath__203_0_I3195 (.Y(N12848), .A(N12593), .B(inst_cellmath__198[25]));
XOR2XL inst_cellmath__203_0_I27946 (.Y(N43395), .A(inst_cellmath__198[24]), .B(inst_cellmath__198[23]));
INVX2 inst_cellmath__203_0_I27947 (.Y(N43396), .A(N43395));
CLKINVX4 inst_cellmath__203_0_I27948 (.Y(N22584), .A(N43396));
INVXL buf1_A_I28632 (.Y(N44110), .A(N43396));
INVXL buf1_A_I28633 (.Y(N11622), .A(N44110));
INVXL inst_cellmath__203_0_I9966 (.Y(N22588), .A(N22584));
CLKINVX4 inst_cellmath__203_0_I9965 (.Y(N22587), .A(N22584));
INVX2 inst_cellmath__203_0_I9964 (.Y(N22586), .A(N22584));
INVXL inst_cellmath__203_0_I9963 (.Y(N22585), .A(N22584));
NAND2X2 inst_cellmath__203_0_I3202 (.Y(N11177), .A(N11620), .B(inst_cellmath__198[25]));
INVX1 inst_cellmath__203_0_I3203 (.Y(N12478), .A(N12848));
NOR2XL inst_cellmath__203_0_I3205 (.Y(N12322), .A(N11288), .B(N11622));
MXI2XL inst_cellmath__203_0_I3206 (.Y(N12641), .A(N12478), .B(N11177), .S0(N12322));
MXI2XL inst_cellmath__203_0_I3207 (.Y(N12261), .A(N12219), .B(N11288), .S0(N22588));
MXI2XL inst_cellmath__203_0_I3208 (.Y(N11290), .A(N12478), .B(N11177), .S0(N12261));
MXI2X1 inst_cellmath__203_0_I3209 (.Y(N12198), .A(N12579), .B(N12219), .S0(N22585));
MXI2X1 inst_cellmath__203_0_I3210 (.Y(N11663), .A(N12478), .B(N11177), .S0(N12198));
MXI2XL inst_cellmath__203_0_I3211 (.Y(N12133), .A(N11223), .B(N12579), .S0(N22585));
MXI2XL inst_cellmath__203_0_I3212 (.Y(N12064), .A(N12478), .B(N11177), .S0(N12133));
MXI2XL inst_cellmath__203_0_I3213 (.Y(N12070), .A(N11600), .B(N11223), .S0(N11622));
MXI2XL inst_cellmath__203_0_I3214 (.Y(N12436), .A(N12478), .B(N11177), .S0(N12070));
MXI2XL inst_cellmath__203_0_I3215 (.Y(N12007), .A(N11999), .B(N11600), .S0(N22585));
MXI2XL inst_cellmath__203_0_I3216 (.Y(N12784), .A(N12478), .B(N11177), .S0(N12007));
MXI2XL inst_cellmath__203_0_I3217 (.Y(N11936), .A(N12373), .B(N11999), .S0(N22585));
MXI2XL inst_cellmath__203_0_I3218 (.Y(N11448), .A(N12478), .B(N11177), .S0(N11936));
MXI2XL inst_cellmath__203_0_I3219 (.Y(N11867), .A(N12720), .B(N12373), .S0(N22585));
MXI2XL inst_cellmath__203_0_I3220 (.Y(N11834), .A(N12478), .B(N11177), .S0(N11867));
MXI2XL inst_cellmath__203_0_I3221 (.Y(N11799), .A(N11377), .B(N12720), .S0(N22586));
MXI2XL inst_cellmath__203_0_I3222 (.Y(N12220), .A(N12478), .B(N11177), .S0(N11799));
MXI2XL inst_cellmath__203_0_I3223 (.Y(N11727), .A(N11761), .B(N11377), .S0(N22586));
MXI2XL inst_cellmath__203_0_I3224 (.Y(N12580), .A(N12478), .B(N11177), .S0(N11727));
MXI2X1 inst_cellmath__203_0_I3225 (.Y(N11662), .A(N12154), .B(N11761), .S0(N22586));
MXI2X1 inst_cellmath__203_0_I3226 (.Y(N11225), .A(N12478), .B(N11177), .S0(N11662));
MXI2X1 inst_cellmath__203_0_I3227 (.Y(N11598), .A(N12523), .B(N12154), .S0(N22586));
MXI2X1 inst_cellmath__203_0_I3228 (.Y(N11601), .A(N12478), .B(N11177), .S0(N11598));
MXI2X1 inst_cellmath__203_0_I3229 (.Y(N11539), .A(N12874), .B(N12523), .S0(N22586));
MXI2X1 inst_cellmath__203_0_I3230 (.Y(N12000), .A(N12478), .B(N11177), .S0(N11539));
MXI2XL inst_cellmath__203_0_I3231 (.Y(N11474), .A(N11540), .B(N12874), .S0(N22587));
MXI2XL inst_cellmath__203_0_I3232 (.Y(N12374), .A(N12478), .B(N11177), .S0(N11474));
MXI2X1 inst_cellmath__203_0_I3233 (.Y(N11405), .A(N11930), .B(N11540), .S0(N22587));
MXI2X1 inst_cellmath__203_0_I3234 (.Y(N12721), .A(N12478), .B(N11177), .S0(N11405));
MXI2X1 inst_cellmath__203_0_I3235 (.Y(N11341), .A(N12313), .B(N11930), .S0(N22587));
MXI2X1 inst_cellmath__203_0_I3236 (.Y(N11378), .A(N12478), .B(N11177), .S0(N11341));
MXI2XL inst_cellmath__203_0_I3237 (.Y(N11278), .A(N12667), .B(N12313), .S0(N22587));
MXI2XL inst_cellmath__203_0_I3238 (.Y(N11763), .A(N12478), .B(N11177), .S0(N11278));
MXI2XL inst_cellmath__203_0_I3239 (.Y(N11212), .A(N11318), .B(N12667), .S0(N22587));
MXI2XL inst_cellmath__203_0_I3240 (.Y(N12155), .A(N12478), .B(N11177), .S0(N11212));
MXI2XL inst_cellmath__203_0_I3241 (.Y(N12865), .A(N11691), .B(N11318), .S0(N22588));
MXI2XL inst_cellmath__203_0_I3242 (.Y(N12525), .A(N12478), .B(N11177), .S0(N12865));
MXI2XL inst_cellmath__203_0_I3243 (.Y(N12803), .A(N12093), .B(N11691), .S0(N22588));
MXI2XL inst_cellmath__203_0_I3244 (.Y(N11161), .A(N12478), .B(N11177), .S0(N12803));
NAND2XL inst_cellmath__203_0_I3245 (.Y(N12741), .A(N12093), .B(N22588));
MXI2XL inst_cellmath__203_0_I3246 (.Y(N11541), .A(N12478), .B(N11177), .S0(N12741));
NOR2XL inst_cellmath__203_0_I3247 (.Y(N12683), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
NAND2XL inst_cellmath__203_0_I3248 (.Y(N11715), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
NOR2X1 inst_cellmath__203_0_I3249 (.Y(N12095), .A(N12683), .B(inst_cellmath__198[27]));
XOR2X1 inst_cellmath__203_0_I3251 (.Y(N12830), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
CLKINVX6 inst_cellmath__203_0_I3252 (.Y(N11497), .A(N12830));
NAND2X2 inst_cellmath__203_0_I10123 (.Y(N12769), .A(N11715), .B(inst_cellmath__198[27]));
INVX2 inst_cellmath__203_0_I3255 (.Y(N11432), .A(N12095));
NOR2XL inst_cellmath__203_0_I3256 (.Y(N12419), .A(N11288), .B(N11497));
MXI2XL inst_cellmath__203_0_I3257 (.Y(N11861), .A(N11432), .B(N12769), .S0(N12419));
MXI2XL inst_cellmath__203_0_I3258 (.Y(N12353), .A(N12219), .B(N11288), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3259 (.Y(N12250), .A(N11432), .B(N12769), .S0(N12353));
MXI2XL inst_cellmath__203_0_I3260 (.Y(N12294), .A(N12579), .B(N12219), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3261 (.Y(N12608), .A(N11432), .B(N12769), .S0(N12294));
MXI2XL inst_cellmath__203_0_I3262 (.Y(N12233), .A(N11223), .B(N12579), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3263 (.Y(N11253), .A(N11432), .B(N12769), .S0(N12233));
MXI2XL inst_cellmath__203_0_I3264 (.Y(N12165), .A(N11600), .B(N11223), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3265 (.Y(N11632), .A(N11432), .B(N12769), .S0(N12165));
MXI2XL inst_cellmath__203_0_I3266 (.Y(N12103), .A(N11999), .B(N11600), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3267 (.Y(N12028), .A(N11432), .B(N12769), .S0(N12103));
MXI2XL inst_cellmath__203_0_I3268 (.Y(N12039), .A(N12373), .B(N11999), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3269 (.Y(N12400), .A(N11432), .B(N12769), .S0(N12039));
MXI2XL inst_cellmath__203_0_I3270 (.Y(N11972), .A(N12720), .B(N12373), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3271 (.Y(N12750), .A(N11432), .B(N12769), .S0(N11972));
MXI2XL inst_cellmath__203_0_I3272 (.Y(N11905), .A(N11377), .B(N12720), .S0(N11497));
MXI2X1 inst_cellmath__203_0_I3273 (.Y(N11408), .A(N11432), .B(N12769), .S0(N11905));
MXI2XL inst_cellmath__203_0_I3274 (.Y(N11839), .A(N11761), .B(N11377), .S0(N11497));
MXI2X1 inst_cellmath__203_0_I3275 (.Y(N11791), .A(N11432), .B(N12769), .S0(N11839));
MXI2X1 inst_cellmath__203_0_I3276 (.Y(N11767), .A(N12154), .B(N11761), .S0(N11497));
MXI2X1 inst_cellmath__203_0_I3277 (.Y(N12183), .A(N11432), .B(N12769), .S0(N11767));
MXI2X1 inst_cellmath__203_0_I3278 (.Y(N11697), .A(N12523), .B(N12154), .S0(N11497));
MXI2X1 inst_cellmath__203_0_I3279 (.Y(N12548), .A(N11432), .B(N12769), .S0(N11697));
MXI2XL inst_cellmath__203_0_I3280 (.Y(N11635), .A(N12874), .B(N12523), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3281 (.Y(N11184), .A(N11432), .B(N12769), .S0(N11635));
MXI2X1 inst_cellmath__203_0_I3282 (.Y(N11571), .A(N11540), .B(N12874), .S0(N11497));
MXI2X1 inst_cellmath__203_0_I3283 (.Y(N11566), .A(N11432), .B(N12769), .S0(N11571));
MXI2XL inst_cellmath__203_0_I3284 (.Y(N11507), .A(N11930), .B(N11540), .S0(N11497));
MXI2X1 inst_cellmath__203_0_I3285 (.Y(N11960), .A(N11432), .B(N12769), .S0(N11507));
MXI2XL inst_cellmath__203_0_I3286 (.Y(N11443), .A(N12313), .B(N11930), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3287 (.Y(N12338), .A(N11432), .B(N12769), .S0(N11443));
MXI2XL inst_cellmath__203_0_I3288 (.Y(N11372), .A(N12667), .B(N12313), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3289 (.Y(N12690), .A(N11432), .B(N12769), .S0(N11372));
MXI2XL inst_cellmath__203_0_I3290 (.Y(N11313), .A(N11318), .B(N12667), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3291 (.Y(N11344), .A(N11432), .B(N12769), .S0(N11313));
MXI2XL inst_cellmath__203_0_I3292 (.Y(N11248), .A(N11691), .B(N11318), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3293 (.Y(N11723), .A(N11432), .B(N12769), .S0(N11248));
MXI2XL inst_cellmath__203_0_I3294 (.Y(N11181), .A(N12093), .B(N11691), .S0(N11497));
MXI2XL inst_cellmath__203_0_I3295 (.Y(N12122), .A(N11432), .B(N12769), .S0(N11181));
NAND2XL inst_cellmath__203_0_I3296 (.Y(N12836), .A(N12093), .B(N11497));
MXI2XL inst_cellmath__203_0_I3297 (.Y(N12491), .A(N11432), .B(N12769), .S0(N12836));
CLKXOR2X1 inst_cellmath__203_0_I3298 (.Y(N12279), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
OA21X1 inst_cellmath__203_0_I10540 (.Y(N11281), .A0(inst_cellmath__198[27]), .A1(inst_cellmath__198[28]), .B0(inst_cellmath__198[29]));
INVX3 inst_cellmath__203_0_I3304 (.Y(N12354), .A(N12279));
INVX3 inst_cellmath__203_0_I9967 (.Y(N22589), .A(N12354));
INVXL inst_cellmath__203_0_I9971 (.Y(N22593), .A(N22589));
CLKINVX4 inst_cellmath__203_0_I9970 (.Y(N22592), .A(N22589));
INVX2 inst_cellmath__203_0_I9968 (.Y(N22590), .A(N22589));
AO21X1 inst_cellmath__203_0_I10542 (.Y(N11915), .A0(inst_cellmath__198[27]), .A1(inst_cellmath__198[28]), .B0(inst_cellmath__198[29]));
INVX1 inst_cellmath__203_0_I3310 (.Y(N12295), .A(N11281));
NOR2XL inst_cellmath__203_0_I3311 (.Y(N12510), .A(N11288), .B(N12354));
MXI2XL inst_cellmath__203_0_I3312 (.Y(N12776), .A(N12295), .B(N11915), .S0(N12510));
MXI2XL inst_cellmath__203_0_I3313 (.Y(N12447), .A(N12219), .B(N11288), .S0(N22593));
MXI2XL inst_cellmath__203_0_I3314 (.Y(N11439), .A(N12295), .B(N11915), .S0(N12447));
MXI2XL inst_cellmath__203_0_I3315 (.Y(N12387), .A(N12579), .B(N12219), .S0(N22590));
MXI2XL inst_cellmath__203_0_I3316 (.Y(N11825), .A(N12295), .B(N11915), .S0(N12387));
MXI2XL inst_cellmath__203_0_I3317 (.Y(N12325), .A(N11223), .B(N12579), .S0(N22590));
MXI2XL inst_cellmath__203_0_I3318 (.Y(N12213), .A(N12295), .B(N11915), .S0(N12325));
MXI2XL inst_cellmath__203_0_I3319 (.Y(N12264), .A(N11600), .B(N11223), .S0(N22590));
MXI2XL inst_cellmath__203_0_I3320 (.Y(N12570), .A(N12295), .B(N11915), .S0(N12264));
MXI2XL inst_cellmath__203_0_I3321 (.Y(N12201), .A(N11999), .B(N11600), .S0(N22590));
MXI2XL inst_cellmath__203_0_I3322 (.Y(N11215), .A(N12295), .B(N11915), .S0(N12201));
MXI2XL inst_cellmath__203_0_I3323 (.Y(N12135), .A(N12373), .B(N11999), .S0(N12354));
MXI2XL inst_cellmath__203_0_I3324 (.Y(N11592), .A(N12295), .B(N11915), .S0(N12135));
MXI2XL inst_cellmath__203_0_I3325 (.Y(N12074), .A(N12720), .B(N12373), .S0(N12354));
MXI2XL inst_cellmath__203_0_I3326 (.Y(N11992), .A(N12295), .B(N11915), .S0(N12074));
MXI2XL inst_cellmath__203_0_I3327 (.Y(N12010), .A(N11377), .B(N12720), .S0(N12354));
MXI2XL inst_cellmath__203_0_I3328 (.Y(N12365), .A(N12295), .B(N11915), .S0(N12010));
MXI2XL inst_cellmath__203_0_I3329 (.Y(N11941), .A(N11761), .B(N11377), .S0(N22592));
MXI2X1 inst_cellmath__203_0_I3330 (.Y(N12714), .A(N12295), .B(N11915), .S0(N11941));
MXI2X1 inst_cellmath__203_0_I3331 (.Y(N11872), .A(N12154), .B(N11761), .S0(N22592));
MXI2X1 inst_cellmath__203_0_I3332 (.Y(N11368), .A(N12295), .B(N11915), .S0(N11872));
MXI2XL inst_cellmath__203_0_I3333 (.Y(N11804), .A(N12523), .B(N12154), .S0(N22592));
MXI2XL inst_cellmath__203_0_I3334 (.Y(N11754), .A(N12295), .B(N11915), .S0(N11804));
MXI2XL inst_cellmath__203_0_I3335 (.Y(N11731), .A(N12874), .B(N12523), .S0(N22592));
MXI2XL inst_cellmath__203_0_I3336 (.Y(N12148), .A(N12295), .B(N11915), .S0(N11731));
MXI2XL inst_cellmath__203_0_I3337 (.Y(N11665), .A(N11540), .B(N12874), .S0(N22592));
MXI2X1 inst_cellmath__203_0_I3338 (.Y(N12515), .A(N12295), .B(N11915), .S0(N11665));
MXI2XL inst_cellmath__203_0_I3339 (.Y(N11603), .A(N11930), .B(N11540), .S0(N22593));
MXI2XL inst_cellmath__203_0_I3340 (.Y(N12868), .A(N12295), .B(N11915), .S0(N11603));
MXI2XL inst_cellmath__203_0_I3341 (.Y(N11543), .A(N12313), .B(N11930), .S0(N22592));
MXI2X1 inst_cellmath__203_0_I3342 (.Y(N11531), .A(N12295), .B(N11915), .S0(N11543));
MXI2XL inst_cellmath__203_0_I3343 (.Y(N11477), .A(N12667), .B(N12313), .S0(N22592));
MXI2XL inst_cellmath__203_0_I3344 (.Y(N11924), .A(N12295), .B(N11915), .S0(N11477));
MXI2XL inst_cellmath__203_0_I3345 (.Y(N11409), .A(N11318), .B(N12667), .S0(N22592));
MXI2XL inst_cellmath__203_0_I3346 (.Y(N12306), .A(N12295), .B(N11915), .S0(N11409));
MXI2XL inst_cellmath__203_0_I3347 (.Y(N11345), .A(N11691), .B(N11318), .S0(N22590));
MXI2XL inst_cellmath__203_0_I3348 (.Y(N12660), .A(N12295), .B(N11915), .S0(N11345));
MXI2XL inst_cellmath__203_0_I3349 (.Y(N11282), .A(N12093), .B(N11691), .S0(N22592));
MXI2XL inst_cellmath__203_0_I3350 (.Y(N11310), .A(N12295), .B(N11915), .S0(N11282));
NAND2XL inst_cellmath__203_0_I3351 (.Y(N11216), .A(N12093), .B(N22592));
MXI2XL inst_cellmath__203_0_I3352 (.Y(N11685), .A(N12295), .B(N11915), .S0(N11216));
NAND2XL inst_cellmath__203_0_I3353 (.Y(N12869), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
NOR2XL inst_cellmath__203_0_I3354 (.Y(N11925), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
AND2XL inst_cellmath__203_0_I3355 (.Y(N12243), .A(inst_cellmath__198[31]), .B(N12869));
XNOR2X2 inst_cellmath__203_0_I10128 (.Y(N11464), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
OR2XL inst_cellmath__203_0_I3359 (.Y(N12734), .A(N11925), .B(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I3360 (.Y(N11392), .A(N12243));
NOR2XL inst_cellmath__203_0_I3361 (.Y(N12600), .A(N11288), .B(N11464));
MXI2XL inst_cellmath__203_0_I3362 (.Y(N12022), .A(N11392), .B(N12734), .S0(N12600));
MXI2XL inst_cellmath__203_0_I3363 (.Y(N12540), .A(N12219), .B(N11288), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3364 (.Y(N12392), .A(N11392), .B(N12734), .S0(N12540));
MXI2XL inst_cellmath__203_0_I3365 (.Y(N12482), .A(N12579), .B(N12219), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3366 (.Y(N12744), .A(N11392), .B(N12734), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3367 (.Y(N12421), .A(N11223), .B(N12579), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3368 (.Y(N11397), .A(N11392), .B(N12734), .S0(N12421));
MXI2XL inst_cellmath__203_0_I3369 (.Y(N12356), .A(N11600), .B(N11223), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3370 (.Y(N11784), .A(N11392), .B(N12734), .S0(N12356));
MXI2XL inst_cellmath__203_0_I3371 (.Y(N12298), .A(N11999), .B(N11600), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3372 (.Y(N12176), .A(N11392), .B(N12734), .S0(N12298));
MXI2XL inst_cellmath__203_0_I3373 (.Y(N12235), .A(N12373), .B(N11999), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3374 (.Y(N12539), .A(N11392), .B(N12734), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3375 (.Y(N12169), .A(N12720), .B(N12373), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3376 (.Y(N11178), .A(N11392), .B(N12734), .S0(N12169));
MXI2XL inst_cellmath__203_0_I3377 (.Y(N12106), .A(N11377), .B(N12720), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3378 (.Y(N11561), .A(N11392), .B(N12734), .S0(N12106));
MXI2XL inst_cellmath__203_0_I3379 (.Y(N12042), .A(N11761), .B(N11377), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3380 (.Y(N11955), .A(N11392), .B(N12734), .S0(N12042));
MXI2XL inst_cellmath__203_0_I3381 (.Y(N11976), .A(N12154), .B(N11761), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3382 (.Y(N12329), .A(N11392), .B(N12734), .S0(N11976));
MXI2XL inst_cellmath__203_0_I3383 (.Y(N11909), .A(N12523), .B(N12154), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3384 (.Y(N12686), .A(N11392), .B(N12734), .S0(N11909));
MXI2XL inst_cellmath__203_0_I3385 (.Y(N11842), .A(N12874), .B(N12523), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3386 (.Y(N11337), .A(N11392), .B(N12734), .S0(N11842));
MXI2XL inst_cellmath__203_0_I3387 (.Y(N11770), .A(N11540), .B(N12874), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3388 (.Y(N11718), .A(N11392), .B(N12734), .S0(N11770));
MXI2XL inst_cellmath__203_0_I3389 (.Y(N11700), .A(N11930), .B(N11540), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3390 (.Y(N12115), .A(N11392), .B(N12734), .S0(N11700));
MXI2XL inst_cellmath__203_0_I3391 (.Y(N11637), .A(N12313), .B(N11930), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3392 (.Y(N12481), .A(N11392), .B(N12734), .S0(N11637));
MXI2XL inst_cellmath__203_0_I3393 (.Y(N11574), .A(N12667), .B(N12313), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3394 (.Y(N12831), .A(N11392), .B(N12734), .S0(N11574));
MXI2XL inst_cellmath__203_0_I3395 (.Y(N11511), .A(N11318), .B(N12667), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3396 (.Y(N11499), .A(N11392), .B(N12734), .S0(N11511));
MXI2XL inst_cellmath__203_0_I3397 (.Y(N11447), .A(N11691), .B(N11318), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3398 (.Y(N11888), .A(N11392), .B(N12734), .S0(N11447));
MXI2XL inst_cellmath__203_0_I3399 (.Y(N11375), .A(N12093), .B(N11691), .S0(N11464));
MXI2XL inst_cellmath__203_0_I3400 (.Y(N12269), .A(N11392), .B(N12734), .S0(N11375));
NAND2XL inst_cellmath__203_0_I3401 (.Y(N11317), .A(N12093), .B(N11464));
MXI2XL inst_cellmath__203_0_I3402 (.Y(N12626), .A(N11392), .B(N12734), .S0(N11317));
ADDHX1 inst_cellmath__203_0_I3403 (.CO(N12770), .S(N12051), .A(inst_cellmath__198[32]), .B(inst_cellmath__198[31]));
INVX2 inst_cellmath__203_0_I3404 (.Y(N11776), .A(N12051));
INVX1 inst_cellmath__203_0_I3405 (.Y(N12166), .A(N12770));
NOR2XL inst_cellmath__203_0_I3406 (.Y(N12706), .A(N11776), .B(N11288));
OAI22XL inst_cellmath__203_0_I3407 (.Y(N11746), .A0(N11288), .A1(N12166), .B0(N11776), .B1(N12219));
OAI22XL inst_cellmath__203_0_I3408 (.Y(N12507), .A0(N12219), .A1(N12166), .B0(N11776), .B1(N12579));
OAI22XL inst_cellmath__203_0_I3409 (.Y(N11526), .A0(N12579), .A1(N12166), .B0(N11776), .B1(N11223));
OAI22XL inst_cellmath__203_0_I3410 (.Y(N12297), .A0(N11223), .A1(N12166), .B0(N11776), .B1(N11600));
OAI22XL inst_cellmath__203_0_I3411 (.Y(N11303), .A0(N11600), .A1(N12166), .B0(N11776), .B1(N11999));
OAI22XL inst_cellmath__203_0_I3412 (.Y(N12078), .A0(N11999), .A1(N12166), .B0(N11776), .B1(N12373));
OAI22XL inst_cellmath__203_0_I3413 (.Y(N12797), .A0(N12373), .A1(N12166), .B0(N11776), .B1(N12720));
OAI22XL inst_cellmath__203_0_I3414 (.Y(N11850), .A0(N12720), .A1(N12166), .B0(N11776), .B1(N11377));
OAI22XL inst_cellmath__203_0_I3415 (.Y(N12592), .A0(N11377), .A1(N12166), .B0(N11776), .B1(N11761));
OAI22XL inst_cellmath__203_0_I3416 (.Y(N11619), .A0(N11761), .A1(N12166), .B0(N11776), .B1(N12154));
OAI22XL inst_cellmath__203_0_I3417 (.Y(N12386), .A0(N12154), .A1(N12166), .B0(N11776), .B1(N12523));
OAI22XL inst_cellmath__203_0_I3418 (.Y(N11393), .A0(N12523), .A1(N12166), .B0(N11776), .B1(N12874));
OAI22XL inst_cellmath__203_0_I3419 (.Y(N12168), .A0(N12874), .A1(N12166), .B0(N11776), .B1(N11540));
OAI22XL inst_cellmath__203_0_I3420 (.Y(N11172), .A0(N11540), .A1(N12166), .B0(N11776), .B1(N11930));
OAI22XL inst_cellmath__203_0_I3421 (.Y(N11945), .A0(N11930), .A1(N12166), .B0(N11776), .B1(N12313));
OAI22XL inst_cellmath__203_0_I3422 (.Y(N12677), .A0(N12313), .A1(N12166), .B0(N11776), .B1(N12667));
OAI22XL inst_cellmath__203_0_I3423 (.Y(N11708), .A0(N12667), .A1(N12166), .B0(N11776), .B1(N11318));
OAI22XL inst_cellmath__203_0_I3424 (.Y(N12471), .A0(N11318), .A1(N12166), .B0(N11776), .B1(N11691));
OAI22XL inst_cellmath__203_0_I3425 (.Y(N11492), .A0(N11691), .A1(N12166), .B0(N11776), .B1(N12093));
OAI21XL inst_cellmath__203_0_I3426 (.Y(N12260), .A0(N12166), .A1(N12093), .B0(N11776));
AND2XL inst_cellmath__203_0_I3427 (.Y(N12749), .A(N12166), .B(N11776));
AND2XL inst_cellmath__203_0_I10129 (.Y(N12534), .A(N8454), .B(N8198));
AND2X1 inst_cellmath__203_0_I10130 (.Y(N11170), .A(N8568), .B(N7684));
AND2X1 inst_cellmath__203_0_I10131 (.Y(N11553), .A(N7817), .B(N8064));
AND2X1 inst_cellmath__203_0_I10132 (.Y(N11944), .A(N8045), .B(N7790));
AND2X1 inst_cellmath__203_0_I10133 (.Y(N12320), .A(N8394), .B(N8636));
CLKAND2X2 inst_cellmath__203_0_I10134 (.Y(N12675), .A(N8754), .B(N8520));
AND2X1 inst_cellmath__203_0_I10135 (.Y(N11330), .A(N7878), .B(N8495));
CLKAND2X2 inst_cellmath__203_0_I10136 (.Y(N11705), .A(N8708), .B(N7851));
AND2X1 inst_cellmath__203_0_I10137 (.Y(N12104), .A(N8069), .B(N8299));
AND2X1 inst_cellmath__203_0_I10138 (.Y(N12470), .A(N8527), .B(N8762));
INVX1 inst_cellmath__203_0_I3438 (.Y(N12823), .A(N770));
INVX2 inst_cellmath__203_0_I3439 (.Y(N11489), .A(N771));
CLKAND2X2 inst_cellmath__203_0_I10141 (.Y(N11876), .A(N8038), .B(N7781));
AND2X1 inst_cellmath__203_0_I10142 (.Y(N12258), .A(N7972), .B(N8344));
AND2X1 inst_cellmath__203_0_I10143 (.Y(N12617), .A(N8424), .B(N8182));
AND2X1 inst_cellmath__203_0_I10144 (.Y(N11265), .A(N8783), .B(N7928));
INVX2 inst_cellmath__203_0_I3444 (.Y(N11643), .A(N776));
CLKAND2X2 inst_cellmath__203_0_I10146 (.Y(N12040), .A(N7834), .B(N8690));
AND2X1 inst_cellmath__203_0_I10147 (.Y(N12412), .A(N8191), .B(N7954));
AND2XL inst_cellmath__203_0_I10148 (.Y(N12760), .A(N8459), .B(N7827));
INVXL inst_cellmath__203_0_I3448 (.Y(N11423), .A(N780));
NOR2XL inst_cellmath__203_0_I3451 (.Y(N12137), .A(N12534), .B(N22568));
NOR2XL inst_cellmath__203_0_I3452 (.Y(N12860), .A(N11170), .B(N22568));
NOR2XL inst_cellmath__203_0_I3453 (.Y(N11914), .A(N11553), .B(N22568));
NOR2XL inst_cellmath__203_0_I3454 (.Y(N12651), .A(N22574), .B(N11944));
NOR2XL inst_cellmath__203_0_I3455 (.Y(N11676), .A(N22574), .B(N12320));
NOR2XL inst_cellmath__203_0_I3456 (.Y(N12444), .A(N22574), .B(N12675));
NOR2XL inst_cellmath__203_0_I3457 (.Y(N11462), .A(N22574), .B(N11330));
NOR2XL inst_cellmath__203_0_I3458 (.Y(N12232), .A(N22574), .B(N11705));
NOR2XL inst_cellmath__203_0_I3459 (.Y(N11237), .A(N22574), .B(N12104));
NOR2XL inst_cellmath__203_0_I3460 (.Y(N12013), .A(N22574), .B(N12470));
NOR2XL inst_cellmath__203_0_I3461 (.Y(N12733), .A(N22574), .B(N12823));
NOR2XL inst_cellmath__203_0_I3462 (.Y(N11775), .A(N22574), .B(N11489));
NOR2XL inst_cellmath__203_0_I3463 (.Y(N12531), .A(N22574), .B(N11876));
NOR2XL inst_cellmath__203_0_I3464 (.Y(N11552), .A(N22574), .B(N12258));
NOR2XL inst_cellmath__203_0_I3465 (.Y(N12319), .A(N22574), .B(N12617));
NOR2XL inst_cellmath__203_0_I3466 (.Y(N11329), .A(N22574), .B(N11265));
NOR2XL inst_cellmath__203_0_I3467 (.Y(N11743), .A(N22574), .B(N11643));
NOR2XL inst_cellmath__203_0_I3468 (.Y(N12469), .A(N22574), .B(N12040));
NOR2XL inst_cellmath__203_0_I3469 (.Y(N11874), .A(N22572), .B(N12412));
NOR2XL inst_cellmath__203_0_I3470 (.Y(N11410), .A(N22572), .B(N12760));
NOR2XL inst_cellmath__203_0_I3471 (.Y(N11373), .A(N22572), .B(N11423));
NOR2XL inst_cellmath__203_0_I3472 (.Y(N12411), .A(N22572), .B(N22540));
NAND2BXL inst_cellmath__203_0_I3474 (.Y(N11293), .AN(N3662), .B(inst_cellmath__61[1]));
INVXL inst_cellmath__203_0_I3475 (.Y(N11668), .A(N3662));
NOR2XL inst_cellmath__203_0_I3476 (.Y(N12689), .A(N12534), .B(N22561));
MXI2XL inst_cellmath__203_0_I3477 (.Y(N12696), .A(N11668), .B(N11293), .S0(N12689));
MXI2XL inst_cellmath__203_0_I3478 (.Y(N12630), .A(N11170), .B(N12534), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3479 (.Y(N11355), .A(N11668), .B(N11293), .S0(N12630));
MXI2XL inst_cellmath__203_0_I3480 (.Y(N12569), .A(N11553), .B(N11170), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3481 (.Y(N11733), .A(N11668), .B(N11293), .S0(N12569));
MXI2XL inst_cellmath__203_0_I3482 (.Y(N12513), .A(N11944), .B(N11553), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3483 (.Y(N12128), .A(N11668), .B(N11293), .S0(N12513));
MXI2XL inst_cellmath__203_0_I3484 (.Y(N12450), .A(N12320), .B(N11944), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3485 (.Y(N12498), .A(N11668), .B(N11293), .S0(N12450));
MXI2XL inst_cellmath__203_0_I3486 (.Y(N12390), .A(N12675), .B(N12320), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3487 (.Y(N12852), .A(N11668), .B(N11293), .S0(N12390));
MXI2XL inst_cellmath__203_0_I3488 (.Y(N12328), .A(N11330), .B(N12675), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3489 (.Y(N11514), .A(N11668), .B(N11293), .S0(N12328));
MXI2XL inst_cellmath__203_0_I3490 (.Y(N12268), .A(N11705), .B(N11330), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3491 (.Y(N11904), .A(N11668), .B(N11293), .S0(N12268));
MXI2XL inst_cellmath__203_0_I3492 (.Y(N12205), .A(N12104), .B(N11705), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3493 (.Y(N12286), .A(N11668), .B(N11293), .S0(N12205));
MXI2XL inst_cellmath__203_0_I3494 (.Y(N12139), .A(N12470), .B(N12104), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3495 (.Y(N12643), .A(N11668), .B(N11293), .S0(N12139));
MXI2XL inst_cellmath__203_0_I3496 (.Y(N12077), .A(N12823), .B(N12470), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3497 (.Y(N11292), .A(N11668), .B(N11293), .S0(N12077));
MXI2XL inst_cellmath__203_0_I3498 (.Y(N12015), .A(N11489), .B(N12823), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3499 (.Y(N11666), .A(N11668), .B(N11293), .S0(N12015));
MXI2X1 inst_cellmath__203_0_I3500 (.Y(N11943), .A(N11876), .B(N11489), .S0(N22561));
MXI2X1 inst_cellmath__203_0_I3501 (.Y(N12066), .A(N11668), .B(N11293), .S0(N11943));
MXI2XL inst_cellmath__203_0_I3502 (.Y(N11875), .A(N12258), .B(N11876), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3503 (.Y(N12438), .A(N11668), .B(N11293), .S0(N11875));
MXI2XL inst_cellmath__203_0_I3504 (.Y(N11806), .A(N12617), .B(N12258), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3505 (.Y(N12789), .A(N11668), .B(N11293), .S0(N11806));
MXI2XL inst_cellmath__203_0_I3506 (.Y(N11734), .A(N11265), .B(N12617), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3507 (.Y(N11451), .A(N11668), .B(N11293), .S0(N11734));
MXI2XL inst_cellmath__203_0_I3508 (.Y(N11667), .A(N11643), .B(N11265), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3509 (.Y(N11837), .A(N11668), .B(N11293), .S0(N11667));
MXI2X1 inst_cellmath__203_0_I3510 (.Y(N11607), .A(N12040), .B(N11643), .S0(N22561));
MXI2X1 inst_cellmath__203_0_I3511 (.Y(N12224), .A(N11668), .B(N11293), .S0(N11607));
MXI2XL inst_cellmath__203_0_I3512 (.Y(N11545), .A(N12412), .B(N12040), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3513 (.Y(N12582), .A(N11668), .B(N11293), .S0(N11545));
MXI2XL inst_cellmath__203_0_I3514 (.Y(N11480), .A(N12760), .B(N12412), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3515 (.Y(N11228), .A(N11668), .B(N11293), .S0(N11480));
MXI2XL inst_cellmath__203_0_I3516 (.Y(N11412), .A(N11423), .B(N12760), .S0(N22561));
MXI2XL inst_cellmath__203_0_I3517 (.Y(N11606), .A(N11668), .B(N11293), .S0(N11412));
MXI2X1 inst_cellmath__203_0_I3518 (.Y(N11347), .A(N22540), .B(N11423), .S0(N22561));
MXI2X1 inst_cellmath__203_0_I3519 (.Y(N12001), .A(N11668), .B(N11293), .S0(N11347));
NOR2BX1 inst_cellmath__203_0_I3520 (.Y(N11285), .AN(N22561), .B(N22540));
MXI2XL inst_cellmath__203_0_I3521 (.Y(N12376), .A(N11668), .B(N11293), .S0(N11285));
XNOR2X1 inst_cellmath__203_0_I3524 (.Y(N12159), .A(N10008), .B(N3662));
NAND2XL inst_cellmath__203_0_I3525 (.Y(N11218), .A(N10008), .B(N3662));
NOR2XL inst_cellmath__203_0_I3526 (.Y(N11995), .A(N10008), .B(N3662));
AND2XL inst_cellmath__203_0_I3529 (.Y(N11164), .A(N11218), .B(N10459));
OR2XL inst_cellmath__203_0_I3530 (.Y(N11481), .A(N11995), .B(N10459));
INVXL inst_cellmath__203_0_I3531 (.Y(N11413), .A(N11164));
NOR2XL inst_cellmath__203_0_I3532 (.Y(N12664), .A(N12534), .B(N12159));
MXI2XL inst_cellmath__203_0_I3533 (.Y(N12671), .A(N11413), .B(N11481), .S0(N12664));
MXI2XL inst_cellmath__203_0_I3534 (.Y(N12603), .A(N11170), .B(N12534), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3535 (.Y(N11321), .A(N11413), .B(N11481), .S0(N12603));
MXI2XL inst_cellmath__203_0_I3536 (.Y(N12543), .A(N11553), .B(N11170), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3537 (.Y(N11696), .A(N11413), .B(N11481), .S0(N12543));
MXI2XL inst_cellmath__203_0_I3538 (.Y(N12485), .A(N11944), .B(N11553), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3539 (.Y(N12097), .A(N11413), .B(N11481), .S0(N12485));
MXI2XL inst_cellmath__203_0_I3540 (.Y(N12424), .A(N12320), .B(N11944), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3541 (.Y(N12461), .A(N11413), .B(N11481), .S0(N12424));
MXI2XL inst_cellmath__203_0_I3542 (.Y(N12359), .A(N12675), .B(N12320), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3543 (.Y(N12816), .A(N11413), .B(N11481), .S0(N12359));
MXI2XL inst_cellmath__203_0_I3544 (.Y(N12302), .A(N11330), .B(N12675), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3545 (.Y(N11479), .A(N11413), .B(N11481), .S0(N12302));
MXI2XL inst_cellmath__203_0_I3546 (.Y(N12238), .A(N11705), .B(N11330), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3547 (.Y(N11863), .A(N11413), .B(N11481), .S0(N12238));
MXI2XL inst_cellmath__203_0_I3548 (.Y(N12171), .A(N12104), .B(N11705), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3549 (.Y(N12252), .A(N11413), .B(N11481), .S0(N12171));
MXI2XL inst_cellmath__203_0_I3550 (.Y(N12110), .A(N12470), .B(N12104), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3551 (.Y(N12611), .A(N11413), .B(N11481), .S0(N12110));
MXI2XL inst_cellmath__203_0_I3552 (.Y(N12046), .A(N12823), .B(N12470), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3553 (.Y(N11256), .A(N11413), .B(N11481), .S0(N12046));
MXI2XL inst_cellmath__203_0_I3554 (.Y(N11980), .A(N11489), .B(N12823), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3555 (.Y(N11634), .A(N11413), .B(N11481), .S0(N11980));
MXI2XL inst_cellmath__203_0_I3556 (.Y(N11912), .A(N11876), .B(N11489), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3557 (.Y(N12030), .A(N11413), .B(N11481), .S0(N11912));
MXI2XL inst_cellmath__203_0_I3558 (.Y(N11846), .A(N12258), .B(N11876), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3559 (.Y(N12402), .A(N11413), .B(N11481), .S0(N11846));
MXI2XL inst_cellmath__203_0_I3560 (.Y(N11773), .A(N12617), .B(N12258), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3561 (.Y(N12752), .A(N11413), .B(N11481), .S0(N11773));
MXI2XL inst_cellmath__203_0_I3562 (.Y(N11703), .A(N11265), .B(N12617), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3563 (.Y(N11411), .A(N11413), .B(N11481), .S0(N11703));
MXI2XL inst_cellmath__203_0_I3564 (.Y(N11641), .A(N11643), .B(N11265), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3565 (.Y(N11793), .A(N11413), .B(N11481), .S0(N11641));
MXI2XL inst_cellmath__203_0_I3566 (.Y(N11578), .A(N12040), .B(N11643), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3567 (.Y(N12186), .A(N11413), .B(N11481), .S0(N11578));
MXI2XL inst_cellmath__203_0_I3568 (.Y(N11513), .A(N12412), .B(N12040), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3569 (.Y(N12552), .A(N11413), .B(N11481), .S0(N11513));
MXI2XL inst_cellmath__203_0_I3570 (.Y(N11450), .A(N12760), .B(N12412), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3571 (.Y(N11188), .A(N11413), .B(N11481), .S0(N11450));
MXI2XL inst_cellmath__203_0_I3572 (.Y(N11380), .A(N11423), .B(N12760), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3573 (.Y(N11570), .A(N11413), .B(N11481), .S0(N11380));
MXI2XL inst_cellmath__203_0_I3574 (.Y(N11320), .A(N22540), .B(N11423), .S0(N12159));
MXI2XL inst_cellmath__203_0_I3575 (.Y(N11963), .A(N11413), .B(N11481), .S0(N11320));
NOR2BX1 inst_cellmath__203_0_I3576 (.Y(N11255), .AN(N12159), .B(N22540));
MXI2XL inst_cellmath__203_0_I3577 (.Y(N12341), .A(N11413), .B(N11481), .S0(N11255));
XNOR2X1 inst_cellmath__203_0_I3578 (.Y(N12123), .A(inst_cellmath__61[5]), .B(N10459));
NAND2XL inst_cellmath__203_0_I3579 (.Y(N11186), .A(inst_cellmath__61[5]), .B(N10459));
NOR2XL inst_cellmath__203_0_I3580 (.Y(N11961), .A(N10459), .B(inst_cellmath__61[5]));
AND2XL inst_cellmath__203_0_I3583 (.Y(N12843), .A(N11186), .B(N3660));
OR2XL inst_cellmath__203_0_I3584 (.Y(N12638), .A(N11961), .B(N3660));
INVXL inst_cellmath__203_0_I3585 (.Y(N12576), .A(N12843));
NOR2XL inst_cellmath__203_0_I3586 (.Y(N12635), .A(N12534), .B(N12123));
MXI2XL inst_cellmath__203_0_I3587 (.Y(N12636), .A(N12576), .B(N12638), .S0(N12635));
MXI2XL inst_cellmath__203_0_I3588 (.Y(N12572), .A(N11170), .B(N12534), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3589 (.Y(N11284), .A(N12576), .B(N12638), .S0(N12572));
MXI2XL inst_cellmath__203_0_I3590 (.Y(N12517), .A(N11553), .B(N11170), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3591 (.Y(N11660), .A(N12576), .B(N12638), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3592 (.Y(N12454), .A(N11944), .B(N11553), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3593 (.Y(N12060), .A(N12576), .B(N12638), .S0(N12454));
MXI2XL inst_cellmath__203_0_I3594 (.Y(N12393), .A(N12320), .B(N11944), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3595 (.Y(N12431), .A(N12576), .B(N12638), .S0(N12393));
MXI2XL inst_cellmath__203_0_I3596 (.Y(N12332), .A(N12675), .B(N12320), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3597 (.Y(N12780), .A(N12576), .B(N12638), .S0(N12332));
MXI2XL inst_cellmath__203_0_I3598 (.Y(N12272), .A(N11330), .B(N12675), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3599 (.Y(N11442), .A(N12576), .B(N12638), .S0(N12272));
MXI2XL inst_cellmath__203_0_I3600 (.Y(N12207), .A(N11705), .B(N11330), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3601 (.Y(N11828), .A(N12576), .B(N12638), .S0(N12207));
MXI2XL inst_cellmath__203_0_I3602 (.Y(N12141), .A(N12104), .B(N11705), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3603 (.Y(N12216), .A(N12576), .B(N12638), .S0(N12141));
MXI2XL inst_cellmath__203_0_I3604 (.Y(N12080), .A(N12470), .B(N12104), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3605 (.Y(N12573), .A(N12576), .B(N12638), .S0(N12080));
MXI2XL inst_cellmath__203_0_I3606 (.Y(N12017), .A(N12823), .B(N12470), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3607 (.Y(N11217), .A(N12576), .B(N12638), .S0(N12017));
MXI2XL inst_cellmath__203_0_I3608 (.Y(N11947), .A(N11489), .B(N12823), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3609 (.Y(N11595), .A(N12576), .B(N12638), .S0(N11947));
MXI2XL inst_cellmath__203_0_I3610 (.Y(N11878), .A(N11876), .B(N11489), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3611 (.Y(N11993), .A(N12576), .B(N12638), .S0(N11878));
MXI2XL inst_cellmath__203_0_I3612 (.Y(N11810), .A(N12258), .B(N11876), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3613 (.Y(N12368), .A(N12576), .B(N12638), .S0(N11810));
MXI2XL inst_cellmath__203_0_I3614 (.Y(N11739), .A(N12617), .B(N12258), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3615 (.Y(N12717), .A(N12576), .B(N12638), .S0(N11739));
MXI2XL inst_cellmath__203_0_I3616 (.Y(N11671), .A(N11265), .B(N12617), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3617 (.Y(N11371), .A(N12576), .B(N12638), .S0(N11671));
MXI2XL inst_cellmath__203_0_I3618 (.Y(N11611), .A(N11643), .B(N11265), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3619 (.Y(N11757), .A(N12576), .B(N12638), .S0(N11611));
MXI2XL inst_cellmath__203_0_I3620 (.Y(N11548), .A(N12040), .B(N11643), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3621 (.Y(N12151), .A(N12576), .B(N12638), .S0(N11548));
MXI2XL inst_cellmath__203_0_I3622 (.Y(N11483), .A(N12412), .B(N12040), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3623 (.Y(N12518), .A(N12576), .B(N12638), .S0(N11483));
MXI2XL inst_cellmath__203_0_I3624 (.Y(N11416), .A(N12760), .B(N12412), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3625 (.Y(N12871), .A(N12576), .B(N12638), .S0(N11416));
MXI2XL inst_cellmath__203_0_I3626 (.Y(N11350), .A(N11423), .B(N12760), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3627 (.Y(N11536), .A(N12576), .B(N12638), .S0(N11350));
MXI2XL inst_cellmath__203_0_I3628 (.Y(N11287), .A(N22540), .B(N11423), .S0(N12123));
MXI2XL inst_cellmath__203_0_I3629 (.Y(N11926), .A(N12576), .B(N12638), .S0(N11287));
NOR2BX1 inst_cellmath__203_0_I3630 (.Y(N11222), .AN(N12123), .B(N22540));
MXI2XL inst_cellmath__203_0_I3631 (.Y(N12309), .A(N12576), .B(N12638), .S0(N11222));
XNOR2X1 inst_cellmath__203_0_I3634 (.Y(N12090), .A(N10179), .B(N3660));
NAND2XL inst_cellmath__203_0_I3635 (.Y(N12875), .A(N10179), .B(N3660));
NOR2XL inst_cellmath__203_0_I3636 (.Y(N11931), .A(N10179), .B(N3660));
AND2XL inst_cellmath__203_0_I3639 (.Y(N12808), .A(N12875), .B(N3666));
OR2XL inst_cellmath__203_0_I3640 (.Y(N12809), .A(N11931), .B(N3666));
INVXL inst_cellmath__203_0_I3641 (.Y(N12747), .A(N12808));
NOR2XL inst_cellmath__203_0_I3642 (.Y(N12606), .A(N12534), .B(N12090));
MXI2XL inst_cellmath__203_0_I3643 (.Y(N12602), .A(N12747), .B(N12809), .S0(N12606));
MXI2XL inst_cellmath__203_0_I3644 (.Y(N12546), .A(N11170), .B(N12534), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3645 (.Y(N11247), .A(N12747), .B(N12809), .S0(N12546));
MXI2XL inst_cellmath__203_0_I3646 (.Y(N12487), .A(N11553), .B(N11170), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3647 (.Y(N11627), .A(N12747), .B(N12809), .S0(N12487));
MXI2XL inst_cellmath__203_0_I3648 (.Y(N12425), .A(N11944), .B(N11553), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3649 (.Y(N12025), .A(N12747), .B(N12809), .S0(N12425));
MXI2XL inst_cellmath__203_0_I3650 (.Y(N12361), .A(N12320), .B(N11944), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3651 (.Y(N12394), .A(N12747), .B(N12809), .S0(N12361));
MXI2XL inst_cellmath__203_0_I3652 (.Y(N12304), .A(N12675), .B(N12320), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3653 (.Y(N12746), .A(N12747), .B(N12809), .S0(N12304));
MXI2XL inst_cellmath__203_0_I3654 (.Y(N12240), .A(N11330), .B(N12675), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3655 (.Y(N11402), .A(N12747), .B(N12809), .S0(N12240));
MXI2XL inst_cellmath__203_0_I3656 (.Y(N12173), .A(N11705), .B(N11330), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3657 (.Y(N11786), .A(N12747), .B(N12809), .S0(N12173));
MXI2XL inst_cellmath__203_0_I3658 (.Y(N12113), .A(N12104), .B(N11705), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3659 (.Y(N12179), .A(N12747), .B(N12809), .S0(N12113));
MXI2XL inst_cellmath__203_0_I3660 (.Y(N12050), .A(N12470), .B(N12104), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3661 (.Y(N12542), .A(N12747), .B(N12809), .S0(N12050));
MXI2XL inst_cellmath__203_0_I3662 (.Y(N11982), .A(N12823), .B(N12470), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3663 (.Y(N11180), .A(N12747), .B(N12809), .S0(N11982));
MXI2XL inst_cellmath__203_0_I3664 (.Y(N11916), .A(N11489), .B(N12823), .S0(N12090));
MXI2X1 inst_cellmath__203_0_I3665 (.Y(N11563), .A(N12747), .B(N12809), .S0(N11916));
MXI2XL inst_cellmath__203_0_I3666 (.Y(N11848), .A(N11876), .B(N11489), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3667 (.Y(N11957), .A(N12747), .B(N12809), .S0(N11848));
MXI2XL inst_cellmath__203_0_I3668 (.Y(N11777), .A(N12258), .B(N11876), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3669 (.Y(N12333), .A(N12747), .B(N12809), .S0(N11777));
MXI2XL inst_cellmath__203_0_I3670 (.Y(N11706), .A(N12617), .B(N12258), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3671 (.Y(N12687), .A(N12747), .B(N12809), .S0(N11706));
MXI2XL inst_cellmath__203_0_I3672 (.Y(N11644), .A(N11265), .B(N12617), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3673 (.Y(N11339), .A(N12747), .B(N12809), .S0(N11644));
MXI2XL inst_cellmath__203_0_I3674 (.Y(N11580), .A(N11643), .B(N11265), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3675 (.Y(N11720), .A(N12747), .B(N12809), .S0(N11580));
MXI2XL inst_cellmath__203_0_I3676 (.Y(N11516), .A(N12040), .B(N11643), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3677 (.Y(N12119), .A(N12747), .B(N12809), .S0(N11516));
MXI2XL inst_cellmath__203_0_I3678 (.Y(N11454), .A(N12412), .B(N12040), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3679 (.Y(N12484), .A(N12747), .B(N12809), .S0(N11454));
MXI2XL inst_cellmath__203_0_I3680 (.Y(N11383), .A(N12760), .B(N12412), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3681 (.Y(N12834), .A(N12747), .B(N12809), .S0(N11383));
MXI2XL inst_cellmath__203_0_I3682 (.Y(N11323), .A(N11423), .B(N12760), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3683 (.Y(N11501), .A(N12747), .B(N12809), .S0(N11323));
MXI2XL inst_cellmath__203_0_I3684 (.Y(N11257), .A(N22540), .B(N11423), .S0(N12090));
MXI2XL inst_cellmath__203_0_I3685 (.Y(N11891), .A(N12747), .B(N12809), .S0(N11257));
NOR2BX1 inst_cellmath__203_0_I3686 (.Y(N11189), .AN(N12090), .B(N22540));
MXI2XL inst_cellmath__203_0_I3687 (.Y(N12273), .A(N12747), .B(N12809), .S0(N11189));
XNOR2X1 inst_cellmath__203_0_I3690 (.Y(N12054), .A(N10521), .B(N3666));
NAND2XL inst_cellmath__203_0_I3691 (.Y(N12844), .A(N10521), .B(N3666));
NOR2XL inst_cellmath__203_0_I3692 (.Y(N11897), .A(N10521), .B(N3666));
INVXL buf1_A_I10789 (.Y(N22721), .A(N3658));
INVXL buf1_A_I10790 (.Y(N12544), .A(N22721));
AND2XL inst_cellmath__203_0_I3695 (.Y(N12773), .A(N12844), .B(N12544));
OR2XL inst_cellmath__203_0_I3696 (.Y(N11276), .A(N11897), .B(N12544));
INVXL inst_cellmath__203_0_I3697 (.Y(N11210), .A(N12773));
NOR2XL inst_cellmath__203_0_I3698 (.Y(N12575), .A(N12534), .B(N12054));
MXI2XL inst_cellmath__203_0_I3699 (.Y(N12567), .A(N11210), .B(N11276), .S0(N12575));
MXI2XL inst_cellmath__203_0_I3700 (.Y(N12520), .A(N11170), .B(N12534), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3701 (.Y(N11208), .A(N11210), .B(N11276), .S0(N12520));
MXI2XL inst_cellmath__203_0_I3702 (.Y(N12456), .A(N11553), .B(N11170), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3703 (.Y(N11590), .A(N11210), .B(N11276), .S0(N12456));
MXI2XL inst_cellmath__203_0_I3704 (.Y(N12396), .A(N11944), .B(N11553), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3705 (.Y(N11985), .A(N11210), .B(N11276), .S0(N12396));
MXI2XL inst_cellmath__203_0_I3706 (.Y(N12335), .A(N12320), .B(N11944), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3707 (.Y(N12358), .A(N11210), .B(N11276), .S0(N12335));
MXI2XL inst_cellmath__203_0_I3708 (.Y(N12275), .A(N12675), .B(N12320), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3709 (.Y(N12711), .A(N11210), .B(N11276), .S0(N12275));
MXI2XL inst_cellmath__203_0_I3710 (.Y(N12210), .A(N11330), .B(N12675), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3711 (.Y(N11362), .A(N11210), .B(N11276), .S0(N12210));
MXI2XL inst_cellmath__203_0_I3712 (.Y(N12144), .A(N11705), .B(N11330), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3713 (.Y(N11748), .A(N11210), .B(N11276), .S0(N12144));
MXI2XL inst_cellmath__203_0_I3714 (.Y(N12084), .A(N12104), .B(N11705), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3715 (.Y(N12143), .A(N11210), .B(N11276), .S0(N12084));
MXI2XL inst_cellmath__203_0_I3716 (.Y(N12020), .A(N12470), .B(N12104), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3717 (.Y(N12508), .A(N11210), .B(N11276), .S0(N12020));
MXI2XL inst_cellmath__203_0_I3718 (.Y(N11950), .A(N12823), .B(N12470), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3719 (.Y(N12862), .A(N11210), .B(N11276), .S0(N11950));
MXI2XL inst_cellmath__203_0_I3720 (.Y(N11882), .A(N11489), .B(N12823), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3721 (.Y(N11529), .A(N11210), .B(N11276), .S0(N11882));
MXI2XL inst_cellmath__203_0_I3722 (.Y(N11814), .A(N11876), .B(N11489), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3723 (.Y(N11919), .A(N11210), .B(N11276), .S0(N11814));
MXI2XL inst_cellmath__203_0_I3724 (.Y(N11741), .A(N12258), .B(N11876), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3725 (.Y(N12300), .A(N11210), .B(N11276), .S0(N11741));
MXI2XL inst_cellmath__203_0_I3726 (.Y(N11674), .A(N12617), .B(N12258), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3727 (.Y(N12658), .A(N11210), .B(N11276), .S0(N11674));
MXI2XL inst_cellmath__203_0_I3728 (.Y(N11615), .A(N11265), .B(N12617), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3729 (.Y(N11304), .A(N11210), .B(N11276), .S0(N11615));
MXI2XL inst_cellmath__203_0_I3730 (.Y(N11550), .A(N11643), .B(N11265), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3731 (.Y(N11680), .A(N11210), .B(N11276), .S0(N11550));
MXI2XL inst_cellmath__203_0_I3732 (.Y(N11487), .A(N12040), .B(N11643), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3733 (.Y(N12083), .A(N11210), .B(N11276), .S0(N11487));
MXI2XL inst_cellmath__203_0_I3734 (.Y(N11420), .A(N12412), .B(N12040), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3735 (.Y(N12446), .A(N11210), .B(N11276), .S0(N11420));
MXI2XL inst_cellmath__203_0_I3736 (.Y(N11353), .A(N12760), .B(N12412), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3737 (.Y(N12799), .A(N11210), .B(N11276), .S0(N11353));
MXI2XL inst_cellmath__203_0_I3738 (.Y(N11291), .A(N11423), .B(N12760), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3739 (.Y(N11467), .A(N11210), .B(N11276), .S0(N11291));
MXI2XL inst_cellmath__203_0_I3740 (.Y(N11226), .A(N22540), .B(N11423), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3741 (.Y(N11852), .A(N11210), .B(N11276), .S0(N11226));
NOR2BX1 inst_cellmath__203_0_I3742 (.Y(N11162), .AN(N12054), .B(N22540));
MXI2XL inst_cellmath__203_0_I3743 (.Y(N12237), .A(N11210), .B(N11276), .S0(N11162));
XNOR2X1 inst_cellmath__203_0_I3744 (.Y(N12019), .A(inst_cellmath__61[11]), .B(N12544));
NAND2XL inst_cellmath__203_0_I3745 (.Y(N12814), .A(inst_cellmath__61[11]), .B(N12544));
NOR2XL inst_cellmath__203_0_I3746 (.Y(N11862), .A(N12544), .B(inst_cellmath__61[11]));
AND2XL inst_cellmath__203_0_I3747 (.Y(N12737), .A(N12814), .B(inst_cellmath__61[12]));
OR2XL inst_cellmath__203_0_I3748 (.Y(N11681), .A(N11862), .B(inst_cellmath__61[12]));
INVXL inst_cellmath__203_0_I3749 (.Y(N11240), .A(N12737));
NOR2XL inst_cellmath__203_0_I3750 (.Y(N12550), .A(N12534), .B(N12019));
MXI2XL inst_cellmath__203_0_I3751 (.Y(N12537), .A(N11240), .B(N11681), .S0(N12550));
MXI2XL inst_cellmath__203_0_I3752 (.Y(N12492), .A(N11170), .B(N12534), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3753 (.Y(N11173), .A(N11240), .B(N11681), .S0(N12492));
MXI2XL inst_cellmath__203_0_I3754 (.Y(N12429), .A(N11553), .B(N11170), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3755 (.Y(N11557), .A(N11240), .B(N11681), .S0(N12429));
MXI2XL inst_cellmath__203_0_I3756 (.Y(N12366), .A(N11944), .B(N11553), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3757 (.Y(N11949), .A(N11240), .B(N11681), .S0(N12366));
MXI2XL inst_cellmath__203_0_I3758 (.Y(N12307), .A(N12320), .B(N11944), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3759 (.Y(N12323), .A(N11240), .B(N11681), .S0(N12307));
MXI2XL inst_cellmath__203_0_I3760 (.Y(N12244), .A(N12675), .B(N12320), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3761 (.Y(N12679), .A(N11240), .B(N11681), .S0(N12244));
MXI2XL inst_cellmath__203_0_I3762 (.Y(N12177), .A(N11330), .B(N12675), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3763 (.Y(N11333), .A(N11240), .B(N11681), .S0(N12177));
MXI2XL inst_cellmath__203_0_I3764 (.Y(N12117), .A(N11705), .B(N11330), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3765 (.Y(N11710), .A(N11240), .B(N11681), .S0(N12117));
MXI2XL inst_cellmath__203_0_I3766 (.Y(N12052), .A(N12104), .B(N11705), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3767 (.Y(N12108), .A(N11240), .B(N11681), .S0(N12052));
MXI2XL inst_cellmath__203_0_I3768 (.Y(N11984), .A(N12470), .B(N12104), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3769 (.Y(N12475), .A(N11240), .B(N11681), .S0(N11984));
MXI2XL inst_cellmath__203_0_I3770 (.Y(N11918), .A(N12823), .B(N12470), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3771 (.Y(N12825), .A(N11240), .B(N11681), .S0(N11918));
MXI2XL inst_cellmath__203_0_I3772 (.Y(N11851), .A(N11489), .B(N12823), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3773 (.Y(N11493), .A(N11240), .B(N11681), .S0(N11851));
MXI2XL inst_cellmath__203_0_I3774 (.Y(N11778), .A(N11876), .B(N11489), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3775 (.Y(N11881), .A(N11240), .B(N11681), .S0(N11778));
MXI2XL inst_cellmath__203_0_I3776 (.Y(N11709), .A(N12258), .B(N11876), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3777 (.Y(N12262), .A(N11240), .B(N11681), .S0(N11709));
MXI2XL inst_cellmath__203_0_I3778 (.Y(N11646), .A(N12617), .B(N12258), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3779 (.Y(N12620), .A(N11240), .B(N11681), .S0(N11646));
MXI2XL inst_cellmath__203_0_I3780 (.Y(N11583), .A(N11265), .B(N12617), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3781 (.Y(N11269), .A(N11240), .B(N11681), .S0(N11583));
MXI2XL inst_cellmath__203_0_I3782 (.Y(N11520), .A(N11643), .B(N11265), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3783 (.Y(N11647), .A(N11240), .B(N11681), .S0(N11520));
MXI2XL inst_cellmath__203_0_I3784 (.Y(N11457), .A(N12040), .B(N11643), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3785 (.Y(N12044), .A(N11240), .B(N11681), .S0(N11457));
MXI2XL inst_cellmath__203_0_I3786 (.Y(N11386), .A(N12412), .B(N12040), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3787 (.Y(N12416), .A(N11240), .B(N11681), .S0(N11386));
MXI2XL inst_cellmath__203_0_I3788 (.Y(N11326), .A(N12760), .B(N12412), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3789 (.Y(N12763), .A(N11240), .B(N11681), .S0(N11326));
MXI2XL inst_cellmath__203_0_I3790 (.Y(N11259), .A(N11423), .B(N12760), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3791 (.Y(N11428), .A(N11240), .B(N11681), .S0(N11259));
MXI2XL inst_cellmath__203_0_I3792 (.Y(N11192), .A(N22540), .B(N11423), .S0(N12019));
MXI2XL inst_cellmath__203_0_I3793 (.Y(N11813), .A(N11240), .B(N11681), .S0(N11192));
NOR2BX1 inst_cellmath__203_0_I3794 (.Y(N12847), .AN(N12019), .B(N22540));
MXI2XL inst_cellmath__203_0_I3795 (.Y(N12199), .A(N11240), .B(N11681), .S0(N12847));
XNOR2X1 inst_cellmath__203_0_I3796 (.Y(N11978), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
NAND2XL inst_cellmath__203_0_I3797 (.Y(N12783), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
NOR2XL inst_cellmath__203_0_I3798 (.Y(N11832), .A(inst_cellmath__61[12]), .B(inst_cellmath__61[13]));
AND2XL inst_cellmath__203_0_I3799 (.Y(N12701), .A(N12783), .B(inst_cellmath__61[14]));
OR2XL inst_cellmath__203_0_I3800 (.Y(N11713), .A(N11832), .B(inst_cellmath__61[14]));
INVXL inst_cellmath__203_0_I3801 (.Y(N11270), .A(N12701));
NOR2XL inst_cellmath__203_0_I3802 (.Y(N12524), .A(N12534), .B(N11978));
MXI2XL inst_cellmath__203_0_I3803 (.Y(N12503), .A(N11270), .B(N11713), .S0(N12524));
MXI2XL inst_cellmath__203_0_I3804 (.Y(N12459), .A(N11170), .B(N12534), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3805 (.Y(N12858), .A(N11270), .B(N11713), .S0(N12459));
MXI2XL inst_cellmath__203_0_I3806 (.Y(N12399), .A(N11553), .B(N11170), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3807 (.Y(N11521), .A(N11270), .B(N11713), .S0(N12399));
MXI2XL inst_cellmath__203_0_I3808 (.Y(N12337), .A(N11944), .B(N11553), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3809 (.Y(N11910), .A(N11270), .B(N11713), .S0(N12337));
MXI2XL inst_cellmath__203_0_I3810 (.Y(N12277), .A(N12320), .B(N11944), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3811 (.Y(N12292), .A(N11270), .B(N11713), .S0(N12277));
MXI2XL inst_cellmath__203_0_I3812 (.Y(N12212), .A(N12675), .B(N12320), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3813 (.Y(N12648), .A(N11270), .B(N11713), .S0(N12212));
MXI2XL inst_cellmath__203_0_I3814 (.Y(N12146), .A(N11330), .B(N12675), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3815 (.Y(N11298), .A(N11270), .B(N11713), .S0(N12146));
MXI2XL inst_cellmath__203_0_I3816 (.Y(N12086), .A(N11705), .B(N11330), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3817 (.Y(N11672), .A(N11270), .B(N11713), .S0(N12086));
MXI2XL inst_cellmath__203_0_I3818 (.Y(N12021), .A(N12104), .B(N11705), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3819 (.Y(N12072), .A(N11270), .B(N11713), .S0(N12021));
MXI2XL inst_cellmath__203_0_I3820 (.Y(N11952), .A(N12470), .B(N12104), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3821 (.Y(N12441), .A(N11270), .B(N11713), .S0(N11952));
MXI2XL inst_cellmath__203_0_I3822 (.Y(N11885), .A(N12823), .B(N12470), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3823 (.Y(N12792), .A(N11270), .B(N11713), .S0(N11885));
MXI2XL inst_cellmath__203_0_I3824 (.Y(N11819), .A(N11489), .B(N12823), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3825 (.Y(N11460), .A(N11270), .B(N11713), .S0(N11819));
MXI2XL inst_cellmath__203_0_I3826 (.Y(N11744), .A(N11876), .B(N11489), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3827 (.Y(N11844), .A(N11270), .B(N11713), .S0(N11744));
MXI2XL inst_cellmath__203_0_I3828 (.Y(N11677), .A(N12258), .B(N11876), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3829 (.Y(N12229), .A(N11270), .B(N11713), .S0(N11677));
MXI2XL inst_cellmath__203_0_I3830 (.Y(N11617), .A(N12617), .B(N12258), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3831 (.Y(N12589), .A(N11270), .B(N11713), .S0(N11617));
MXI2XL inst_cellmath__203_0_I3832 (.Y(N11554), .A(N11265), .B(N12617), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3833 (.Y(N11233), .A(N11270), .B(N11713), .S0(N11554));
MXI2XL inst_cellmath__203_0_I3834 (.Y(N11490), .A(N11643), .B(N11265), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3835 (.Y(N11613), .A(N11270), .B(N11713), .S0(N11490));
MXI2XL inst_cellmath__203_0_I3836 (.Y(N11424), .A(N12040), .B(N11643), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3837 (.Y(N12012), .A(N11270), .B(N11713), .S0(N11424));
MXI2XL inst_cellmath__203_0_I3838 (.Y(N11356), .A(N12412), .B(N12040), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3839 (.Y(N12381), .A(N11270), .B(N11713), .S0(N11356));
MXI2XL inst_cellmath__203_0_I3840 (.Y(N11294), .A(N12760), .B(N12412), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3841 (.Y(N12730), .A(N11270), .B(N11713), .S0(N11294));
MXI2XL inst_cellmath__203_0_I3842 (.Y(N11230), .A(N11423), .B(N12760), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3843 (.Y(N11389), .A(N11270), .B(N11713), .S0(N11230));
MXI2XL inst_cellmath__203_0_I3844 (.Y(N11165), .A(N22540), .B(N11423), .S0(N11978));
MXI2XL inst_cellmath__203_0_I3845 (.Y(N11771), .A(N11270), .B(N11713), .S0(N11165));
NOR2BX1 inst_cellmath__203_0_I3846 (.Y(N12817), .AN(N11978), .B(N22540));
MXI2XL inst_cellmath__203_0_I3847 (.Y(N12270), .A(N11270), .B(N11713), .S0(N12817));
XNOR2X1 inst_cellmath__203_0_I3848 (.Y(N11940), .A(inst_cellmath__61[14]), .B(inst_cellmath__61[15]));
NAND2XL inst_cellmath__203_0_I3849 (.Y(N12753), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
NOR2XL inst_cellmath__203_0_I3850 (.Y(N11796), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
AND2XL inst_cellmath__203_0_I3851 (.Y(N12674), .A(N12753), .B(inst_cellmath__115__W1[0]));
OR2XL inst_cellmath__203_0_I3852 (.Y(N11742), .A(N11796), .B(inst_cellmath__115__W1[0]));
INVXL inst_cellmath__203_0_I3853 (.Y(inst_cellmath__203__W0[42]), .A(N12674));
NOR2XL inst_cellmath__203_0_I3854 (.Y(N12494), .A(N12534), .B(N11940));
MXI2XL inst_cellmath__203_0_I3855 (.Y(N12467), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12494));
MXI2XL inst_cellmath__203_0_I3856 (.Y(N12432), .A(N11170), .B(N12534), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3857 (.Y(N12819), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12432));
MXI2XL inst_cellmath__203_0_I3858 (.Y(N12370), .A(N11553), .B(N11170), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3859 (.Y(N11485), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12370));
MXI2XL inst_cellmath__203_0_I3860 (.Y(N12310), .A(N11944), .B(N11553), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3861 (.Y(N11871), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12310));
MXI2XL inst_cellmath__203_0_I3862 (.Y(N12246), .A(N12320), .B(N11944), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3863 (.Y(N12254), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12246));
MXI2XL inst_cellmath__203_0_I3864 (.Y(N12181), .A(N12675), .B(N12320), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3865 (.Y(N12614), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12181));
MXI2XL inst_cellmath__203_0_I3866 (.Y(N12120), .A(N11330), .B(N12675), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3867 (.Y(N11262), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12120));
MXI2XL inst_cellmath__203_0_I3868 (.Y(N12055), .A(N11705), .B(N11330), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3869 (.Y(N11638), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12055));
MXI2XL inst_cellmath__203_0_I3870 (.Y(N11988), .A(N12104), .B(N11705), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3871 (.Y(N12035), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11988));
MXI2XL inst_cellmath__203_0_I3872 (.Y(N11921), .A(N12470), .B(N12104), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3873 (.Y(N12408), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11921));
MXI2XL inst_cellmath__203_0_I3874 (.Y(N11855), .A(N12823), .B(N12470), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3875 (.Y(N12756), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11855));
MXI2XL inst_cellmath__203_0_I3876 (.Y(N11781), .A(N11489), .B(N12823), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3877 (.Y(N11418), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11781));
MXI2XL inst_cellmath__203_0_I3878 (.Y(N11712), .A(N11876), .B(N11489), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3879 (.Y(N11803), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11712));
MXI2XL inst_cellmath__203_0_I3880 (.Y(N11650), .A(N12258), .B(N11876), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3881 (.Y(N12190), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11650));
MXI2XL inst_cellmath__203_0_I3882 (.Y(N11585), .A(N12617), .B(N12258), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3883 (.Y(N12556), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11585));
MXI2XL inst_cellmath__203_0_I3884 (.Y(N11524), .A(N11265), .B(N12617), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3885 (.Y(N11195), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11524));
MXI2XL inst_cellmath__203_0_I3886 (.Y(N11461), .A(N11643), .B(N11265), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3887 (.Y(N11575), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11461));
MXI2XL inst_cellmath__203_0_I3888 (.Y(N11390), .A(N12040), .B(N11643), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3889 (.Y(N11968), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11390));
MXI2XL inst_cellmath__203_0_I3890 (.Y(N11327), .A(N12412), .B(N12040), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3891 (.Y(N12345), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11327));
MXI2XL inst_cellmath__203_0_I3892 (.Y(N11263), .A(N12760), .B(N12412), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3893 (.Y(N12695), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11263));
MXI2XL inst_cellmath__203_0_I3894 (.Y(N11196), .A(N11423), .B(N12760), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3895 (.Y(N11352), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N11196));
MXI2XL inst_cellmath__203_0_I3896 (.Y(N12850), .A(N22540), .B(N11423), .S0(N11940));
MXI2XL inst_cellmath__203_0_I3897 (.Y(N11730), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12850));
NOR2BX1 inst_cellmath__203_0_I3898 (.Y(N12786), .AN(N11940), .B(N22540));
MXI2XL inst_cellmath__203_0_I3899 (.Y(inst_cellmath__203__W1[42]), .A(inst_cellmath__203__W0[42]), .B(N11742), .S0(N12786));
ADDHX1 inst_cellmath__203_0_I3900 (.CO(N11343), .S(inst_cellmath__203__W1[1]), .A(N12835), .B(inst_cellmath__198[19]));
ADDHX1 inst_cellmath__203_0_I3901 (.CO(inst_cellmath__203__W0[3]), .S(inst_cellmath__203__W1[2]), .A(N11889), .B(N11343));
ADDHX1 inst_cellmath__203_0_I3902 (.CO(N12841), .S(N12490), .A(N12628), .B(N12702));
ADDFX1 inst_cellmath__203_0_I3903 (.CO(N11895), .S(inst_cellmath__203__W1[3]), .A(N12490), .B(N12324), .CI(N12504));
ADDFX1 inst_cellmath__203_0_I3904 (.CO(N12632), .S(inst_cellmath__203__W0[4]), .A(N11653), .B(N12137), .CI(N12680));
ADDFX1 inst_cellmath__203_0_I3905 (.CO(inst_cellmath__203__W0[5]), .S(inst_cellmath__203__W1[4]), .A(N12856), .B(N12841), .CI(N11895));
ADDFX1 inst_cellmath__203_0_I3906 (.CO(N12428), .S(N12058), .A(N12860), .B(N3662), .CI(N12696));
ADDFX1 inst_cellmath__203_0_I3907 (.CO(N11438), .S(N12778), .A(N12422), .B(N12058), .CI(N11938));
ADDFX1 inst_cellmath__203_0_I3908 (.CO(N12214), .S(N11824), .A(N11701), .B(N11332), .CI(N11522));
ADDFXL inst_cellmath__203_0_I3909 (.CO(inst_cellmath__203__W0[6]), .S(inst_cellmath__203__W1[5]), .A(N12632), .B(N12778), .CI(N11824));
ADDFX1 inst_cellmath__203_0_I3910 (.CO(N11991), .S(N11593), .A(N11355), .B(N11914), .CI(N12428));
ADDFX1 inst_cellmath__203_0_I3911 (.CO(N12716), .S(N12364), .A(N11435), .B(N11593), .CI(N11711));
ADDFXL inst_cellmath__203_0_I3912 (.CO(N11753), .S(N11367), .A(N11438), .B(N11911), .CI(N12101));
ADDFXL inst_cellmath__203_0_I3913 (.CO(inst_cellmath__203__W0[7]), .S(inst_cellmath__203__W1[6]), .A(N12214), .B(N12364), .CI(N11367));
ADDFX1 inst_cellmath__203_0_I3914 (.CO(N11533), .S(N12867), .A(N12651), .B(N11164), .CI(N11733));
ADDFX1 inst_cellmath__203_0_I3915 (.CO(N12305), .S(N11923), .A(N12867), .B(N12671), .CI(N11991));
ADDFX1 inst_cellmath__203_0_I3916 (.CO(N11309), .S(N12662), .A(N11923), .B(N12208), .CI(N12848));
ADDFX1 inst_cellmath__203_0_I3917 (.CO(N12088), .S(N11684), .A(N12290), .B(N12109), .CI(N12641));
ADDFX1 inst_cellmath__203_0_I3918 (.CO(N12806), .S(N12452), .A(N12662), .B(N12465), .CI(N12716));
ADDFX1 inst_cellmath__203_0_I3919 (.CO(inst_cellmath__203__W0[8]), .S(inst_cellmath__203__W1[7]), .A(N11684), .B(N11753), .CI(N12452));
ADDFX1 inst_cellmath__203_0_I3920 (.CO(N12599), .S(N12242), .A(N12128), .B(N11676), .CI(N11321));
ADDFX1 inst_cellmath__203_0_I3921 (.CO(N11624), .S(N11244), .A(N12242), .B(N11533), .CI(N12305));
ADDFX1 inst_cellmath__203_0_I3922 (.CO(N12391), .S(N12023), .A(N11244), .B(N11209), .CI(N12473));
ADDFX1 inst_cellmath__203_0_I3923 (.CO(N11399), .S(N12743), .A(N11309), .B(N12649), .CI(N11290));
ADDFX1 inst_cellmath__203_0_I3924 (.CO(N12175), .S(N11783), .A(N12023), .B(N12820), .CI(N12088));
ADDFX1 inst_cellmath__203_0_I3925 (.CO(inst_cellmath__203__W0[9]), .S(inst_cellmath__203__W1[8]), .A(N12743), .B(N12806), .CI(N11783));
ADDFX1 inst_cellmath__203_0_I3926 (.CO(N11954), .S(N11560), .A(N12444), .B(N12843), .CI(N11696));
ADDFX1 inst_cellmath__203_0_I3927 (.CO(N12685), .S(N12331), .A(N12636), .B(N12498), .CI(N12599));
ADDFX1 inst_cellmath__203_0_I3928 (.CO(N11719), .S(N11336), .A(N12331), .B(N11560), .CI(N11986));
ADDFX1 inst_cellmath__203_0_I3929 (.CO(N12480), .S(N12114), .A(N11624), .B(N12095), .CI(N11336));
ADDFX1 inst_cellmath__203_0_I3930 (.CO(N11498), .S(N12833), .A(N12826), .B(N11861), .CI(N11299));
ADDFX1 inst_cellmath__203_0_I3931 (.CO(N12271), .S(N11887), .A(N11486), .B(N11663), .CI(N12114));
ADDFX1 inst_cellmath__203_0_I3932 (.CO(N11273), .S(N12625), .A(N11399), .B(N12391), .CI(N12833));
ADDFXL inst_cellmath__203_0_I3933 (.CO(inst_cellmath__203__W0[10]), .S(inst_cellmath__203__W1[9]), .A(N12175), .B(N11887), .CI(N12625));
ADDFX1 inst_cellmath__203_0_I3934 (.CO(N12772), .S(N12420), .A(N12097), .B(N11462), .CI(N11284));
ADDFX1 inst_cellmath__203_0_I3935 (.CO(N11820), .S(N11433), .A(N11954), .B(N12852), .CI(N12420));
ADDFX1 inst_cellmath__203_0_I3936 (.CO(N12565), .S(N12206), .A(N11433), .B(N12685), .CI(N12709));
ADDFX1 inst_cellmath__203_0_I3937 (.CO(N11588), .S(N11205), .A(N12206), .B(N11719), .CI(N11494));
ADDFXL inst_cellmath__203_0_I3938 (.CO(N12355), .S(N11983), .A(N11673), .B(N12250), .CI(N12480));
ADDFX1 inst_cellmath__203_0_I3939 (.CO(N11361), .S(N12708), .A(N11869), .B(N12064), .CI(N11205));
ADDFXL inst_cellmath__203_0_I3940 (.CO(N12140), .S(N11745), .A(N12271), .B(N11498), .CI(N11983));
ADDFXL inst_cellmath__203_0_I3941 (.CO(inst_cellmath__203__W0[11]), .S(inst_cellmath__203__W1[10]), .A(N11273), .B(N12708), .CI(N11745));
ADDFX1 inst_cellmath__203_0_I3942 (.CO(N11917), .S(N11527), .A(N12232), .B(N12808), .CI(N11514));
ADDFX1 inst_cellmath__203_0_I3943 (.CO(N12656), .S(N12296), .A(N12461), .B(N11660), .CI(N12602));
ADDFX1 inst_cellmath__203_0_I3944 (.CO(N11678), .S(N11302), .A(N11527), .B(N12772), .CI(N12296));
ADDFX1 inst_cellmath__203_0_I3945 (.CO(N12445), .S(N12079), .A(N11302), .B(N11820), .CI(N11749));
ADDFX1 inst_cellmath__203_0_I3946 (.CO(N11465), .S(N12796), .A(N12079), .B(N12565), .CI(N11281));
ADDFX1 inst_cellmath__203_0_I3947 (.CO(N12234), .S(N11849), .A(N12073), .B(N11879), .CI(N12608));
ADDFX1 inst_cellmath__203_0_I3948 (.CO(N11238), .S(N12594), .A(N12255), .B(N12436), .CI(N12776));
ADDFX1 inst_cellmath__203_0_I3949 (.CO(N12016), .S(N11618), .A(N11588), .B(N12796), .CI(N12355));
ADDFX1 inst_cellmath__203_0_I3950 (.CO(N12735), .S(N12385), .A(N11361), .B(N11849), .CI(N12594));
ADDFX1 inst_cellmath__203_0_I3951 (.CO(inst_cellmath__203__W0[12]), .S(inst_cellmath__203__W1[11]), .A(N12140), .B(N11618), .CI(N12385));
ADDFX1 inst_cellmath__203_0_I3952 (.CO(N12535), .S(N12167), .A(N11904), .B(N11237), .CI(N12060));
ADDFX1 inst_cellmath__203_0_I3953 (.CO(N11555), .S(N11171), .A(N11247), .B(N12816), .CI(N11917));
ADDFX1 inst_cellmath__203_0_I3954 (.CO(N12321), .S(N11946), .A(N12167), .B(N12656), .CI(N11171));
ADDFX1 inst_cellmath__203_0_I3955 (.CO(N11331), .S(N12676), .A(N12509), .B(N11678), .CI(N11946));
ADDFX1 inst_cellmath__203_0_I3956 (.CO(N12105), .S(N11707), .A(N12263), .B(N12445), .CI(N12676));
ADDFX1 inst_cellmath__203_0_I3957 (.CO(N12824), .S(N12472), .A(N11253), .B(N12442), .CI(N11465));
ADDFX1 inst_cellmath__203_0_I3958 (.CO(N11877), .S(N11491), .A(N12615), .B(N12784), .CI(N11439));
ADDFX1 inst_cellmath__203_0_I3959 (.CO(N12618), .S(N12259), .A(N11707), .B(N12234), .CI(N11238));
ADDFX1 inst_cellmath__203_0_I3960 (.CO(N11645), .S(N11266), .A(N11491), .B(N12472), .CI(N12016));
ADDFX1 inst_cellmath__203_0_I3961 (.CO(inst_cellmath__203__W0[13]), .S(inst_cellmath__203__W1[12]), .A(N12735), .B(N12259), .CI(N11266));
ADDFX1 inst_cellmath__203_0_I3962 (.CO(N11425), .S(N12761), .A(N12013), .B(N12773), .CI(N11479));
ADDFX1 inst_cellmath__203_0_I3963 (.CO(N12196), .S(N11809), .A(N12431), .B(N11627), .CI(N12567));
ADDFX1 inst_cellmath__203_0_I3964 (.CO(N11199), .S(N12559), .A(N12535), .B(N12286), .CI(N12761));
ADDFX1 inst_cellmath__203_0_I3965 (.CO(N11973), .S(N11582), .A(N11555), .B(N11809), .CI(N12559));
ADDFX1 inst_cellmath__203_0_I3966 (.CO(N12700), .S(N12348), .A(N12321), .B(N11528), .CI(N11582));
ADDFX1 inst_cellmath__203_0_I3967 (.CO(N11737), .S(N11357), .A(N12621), .B(N11331), .CI(N12243));
ADDFX1 inst_cellmath__203_0_I3968 (.CO(N12499), .S(N12134), .A(N12348), .B(N12793), .CI(N11632));
ADDFX1 inst_cellmath__203_0_I3969 (.CO(N11519), .S(N12854), .A(N11260), .B(N11448), .CI(N11825));
ADDFX1 inst_cellmath__203_0_I3970 (.CO(N12288), .S(N11906), .A(N12105), .B(N12022), .CI(N11357));
ADDFX1 inst_cellmath__203_0_I3971 (.CO(N11295), .S(N12647), .A(N11877), .B(N12824), .CI(N12134));
ADDFX1 inst_cellmath__203_0_I3972 (.CO(N12071), .S(N11670), .A(N12618), .B(N12854), .CI(N11906));
ADDFXL inst_cellmath__203_0_I3973 (.CO(inst_cellmath__203__W0[14]), .S(inst_cellmath__203__W1[13]), .A(N11645), .B(N12647), .CI(N11670));
ADDFX1 inst_cellmath__203_0_I3974 (.CO(N11840), .S(N11456), .A(N11863), .B(N12733), .CI(N12025));
ADDFX1 inst_cellmath__203_0_I3975 (.CO(N12586), .S(N12226), .A(N11208), .B(N12780), .CI(N12643));
ADDFX1 inst_cellmath__203_0_I3976 (.CO(N11610), .S(N11231), .A(N12196), .B(N11425), .CI(N11456));
ADDFX1 inst_cellmath__203_0_I3977 (.CO(N12379), .S(N12008), .A(N11199), .B(N12226), .CI(N11231));
ADDFX1 inst_cellmath__203_0_I3978 (.CO(N11385), .S(N12728), .A(N11973), .B(N12301), .CI(N12008));
ADDFXL inst_cellmath__203_0_I3979 (.CO(N12161), .S(N11768), .A(N11267), .B(N12700), .CI(N11458));
ADDFX1 inst_cellmath__203_0_I3980 (.CO(N11166), .S(N12529), .A(N12028), .B(N11639), .CI(N11834));
ADDFX1 inst_cellmath__203_0_I3981 (.CO(N11937), .S(N11547), .A(N12213), .B(N12728), .CI(N12392));
ADDFXL inst_cellmath__203_0_I3982 (.CO(N12673), .S(N12316), .A(N12499), .B(N11737), .CI(N11768));
ADDFX1 inst_cellmath__203_0_I3983 (.CO(N11698), .S(N11325), .A(N12529), .B(N11519), .CI(N12288));
ADDFX1 inst_cellmath__203_0_I3984 (.CO(N12464), .S(N12099), .A(N11295), .B(N11547), .CI(N12316));
ADDFXL inst_cellmath__203_0_I3985 (.CO(inst_cellmath__203__W0[15]), .S(inst_cellmath__203__W1[14]), .A(N11325), .B(N12071), .CI(N12099));
ADDHX1 inst_cellmath__203_0_I3986 (.CO(N12253), .S(N11868), .A(N12737), .B(N11775));
ADDFX1 inst_cellmath__203_0_I3987 (.CO(N11258), .S(N12612), .A(N11442), .B(N11868), .CI(N11292));
ADDFX1 inst_cellmath__203_0_I3988 (.CO(N12033), .S(N11636), .A(N12394), .B(N11590), .CI(N12537));
ADDFX1 inst_cellmath__203_0_I3989 (.CO(N12754), .S(N12405), .A(N11840), .B(N12252), .CI(N12586));
ADDFX1 inst_cellmath__203_0_I3990 (.CO(N11800), .S(N11415), .A(N11636), .B(N12612), .CI(N11610));
ADDFX1 inst_cellmath__203_0_I3991 (.CO(N12554), .S(N12188), .A(N11305), .B(N12405), .CI(N12379));
ADDFX1 inst_cellmath__203_0_I3992 (.CO(N11572), .S(N11191), .A(N11648), .B(N11415), .CI(N12706));
ADDFX1 inst_cellmath__203_0_I3993 (.CO(N12343), .S(N11966), .A(N12188), .B(N11385), .CI(N11845));
ADDFX1 inst_cellmath__203_0_I3994 (.CO(N11349), .S(N12693), .A(N12220), .B(N12400), .CI(N12036));
ADDFX1 inst_cellmath__203_0_I3995 (.CO(N12125), .S(N11728), .A(N12744), .B(N12570), .CI(N12161));
ADDFXL inst_cellmath__203_0_I3996 (.CO(N12846), .S(N12496), .A(N11166), .B(N11191), .CI(N11966));
ADDFX1 inst_cellmath__203_0_I3997 (.CO(N11900), .S(N11509), .A(N12693), .B(N11937), .CI(N12673));
ADDFXL inst_cellmath__203_0_I3998 (.CO(N12639), .S(N12283), .A(N12496), .B(N11728), .CI(N11698));
ADDFXL inst_cellmath__203_0_I3999 (.CO(inst_cellmath__203__W0[16]), .S(inst_cellmath__203__W1[15]), .A(N12464), .B(N11509), .CI(N12283));
ADDFX1 inst_cellmath__203_0_I4000 (.CO(N12433), .S(N12062), .A(N12253), .B(N12531), .CI(N11828));
ADDFX1 inst_cellmath__203_0_I4001 (.CO(N11445), .S(N12782), .A(N11985), .B(N11666), .CI(N12611));
ADDFX1 inst_cellmath__203_0_I4002 (.CO(N12218), .S(N11830), .A(N11173), .B(N12746), .CI(N11258));
ADDFXL inst_cellmath__203_0_I4003 (.CO(N11220), .S(N12578), .A(N12062), .B(N12033), .CI(N12782));
ADDFXL inst_cellmath__203_0_I4004 (.CO(N11998), .S(N11599), .A(N11830), .B(N12754), .CI(N12578));
ADDFX1 inst_cellmath__203_0_I4005 (.CO(N12719), .S(N12371), .A(N11800), .B(N12081), .CI(N11599));
ADDFX1 inst_cellmath__203_0_I4006 (.CO(N11758), .S(N11376), .A(N12045), .B(N12554), .CI(N12230));
ADDFXL inst_cellmath__203_0_I4007 (.CO(N12522), .S(N12153), .A(N11746), .B(N12750), .CI(N12580));
ADDFX1 inst_cellmath__203_0_I4008 (.CO(N11538), .S(N12872), .A(N12371), .B(N12406), .CI(N11215));
ADDFX1 inst_cellmath__203_0_I4009 (.CO(N12311), .S(N11929), .A(N11572), .B(N11397), .CI(N12343));
ADDFX1 inst_cellmath__203_0_I4010 (.CO(N11316), .S(N12665), .A(N11349), .B(N11376), .CI(N12153));
ADDFX1 inst_cellmath__203_0_I4011 (.CO(N12091), .S(N11688), .A(N12125), .B(N12872), .CI(N11929));
ADDFX1 inst_cellmath__203_0_I4012 (.CO(N12810), .S(N12458), .A(N12665), .B(N12846), .CI(N11900));
ADDFX1 inst_cellmath__203_0_I4013 (.CO(inst_cellmath__203__W0[17]), .S(inst_cellmath__203__W1[16]), .A(N12639), .B(N11688), .CI(N12458));
ADDFXL inst_cellmath__203_0_I4014 (.CO(N12604), .S(N12247), .A(N11552), .B(N12701), .CI(N12066));
ADDFX1 inst_cellmath__203_0_I4015 (.CO(N11628), .S(N11251), .A(N11557), .B(N11402), .CI(N12358));
ADDFX1 inst_cellmath__203_0_I4016 (.CO(N12398), .S(N12026), .A(N12503), .B(N11256), .CI(N12216));
ADDFX1 inst_cellmath__203_0_I4017 (.CO(N11404), .S(N12748), .A(N11445), .B(N12433), .CI(N12247));
ADDFX1 inst_cellmath__203_0_I4018 (.CO(N12182), .S(N11790), .A(N12026), .B(N11251), .CI(N12218));
ADDFX1 inst_cellmath__203_0_I4019 (.CO(N11182), .S(N12545), .A(N12748), .B(N11220), .CI(N12800));
ADDFX1 inst_cellmath__203_0_I4020 (.CO(N11958), .S(N11564), .A(N11790), .B(N11998), .CI(N12545));
ADDFXL inst_cellmath__203_0_I4021 (.CO(N12688), .S(N12336), .A(N12719), .B(N12414), .CI(N12587));
ADDFXL inst_cellmath__203_0_I4022 (.CO(N11722), .S(N11340), .A(N12507), .B(N11408), .CI(N11225));
ADDFX1 inst_cellmath__203_0_I4023 (.CO(N12486), .S(N12121), .A(N11592), .B(N12757), .CI(N11564));
ADDFX1 inst_cellmath__203_0_I4024 (.CO(N11502), .S(N12838), .A(N11758), .B(N11784), .CI(N12522));
ADDFXL inst_cellmath__203_0_I4025 (.CO(N12276), .S(N11892), .A(N11538), .B(N12336), .CI(N11340));
ADDFXL inst_cellmath__203_0_I4026 (.CO(N11277), .S(N12629), .A(N12121), .B(N12311), .CI(N11316));
ADDFX1 inst_cellmath__203_0_I4027 (.CO(N12056), .S(N11655), .A(N11892), .B(N12838), .CI(N12091));
ADDFX1 inst_cellmath__203_0_I4028 (.CO(inst_cellmath__203__W0[18]), .S(inst_cellmath__203__W1[17]), .A(N12810), .B(N12629), .CI(N11655));
ADDFX1 inst_cellmath__203_0_I4029 (.CO(N11823), .S(N11436), .A(N11786), .B(N12319), .CI(N12711));
ADDFX1 inst_cellmath__203_0_I4030 (.CO(N12568), .S(N12211), .A(N11949), .B(N11634), .CI(N12573));
ADDFXL inst_cellmath__203_0_I4031 (.CO(N11591), .S(N11211), .A(N12858), .B(N12438), .CI(N12604));
ADDFX1 inst_cellmath__203_0_I4032 (.CO(N12360), .S(N11989), .A(N12398), .B(N11628), .CI(N11436));
ADDFX1 inst_cellmath__203_0_I4033 (.CO(N11364), .S(N12712), .A(N12211), .B(N11211), .CI(N11404));
ADDFXL inst_cellmath__203_0_I4034 (.CO(N12145), .S(N11750), .A(N11989), .B(N12182), .CI(N11853));
ADDFXL inst_cellmath__203_0_I4035 (.CO(N12864), .S(N12512), .A(N11182), .B(N12712), .CI(N11750));
ADDFXL inst_cellmath__203_0_I4036 (.CO(N11922), .S(N11530), .A(N12764), .B(N11958), .CI(N11234));
ADDFXL inst_cellmath__203_0_I4037 (.CO(N12659), .S(N12303), .A(N11791), .B(N11526), .CI(N11601));
ADDFX1 inst_cellmath__203_0_I4038 (.CO(N11682), .S(N11307), .A(N11992), .B(N11419), .CI(N12512));
ADDFX1 inst_cellmath__203_0_I4039 (.CO(N12449), .S(N12085), .A(N12688), .B(N12176), .CI(N11722));
ADDFXL inst_cellmath__203_0_I4040 (.CO(N11468), .S(N12802), .A(N11530), .B(N12486), .CI(N12303));
ADDFXL inst_cellmath__203_0_I4041 (.CO(N12239), .S(N11856), .A(N11502), .B(N11307), .CI(N12276));
ADDFXL inst_cellmath__203_0_I4042 (.CO(N11242), .S(N12597), .A(N12802), .B(N12085), .CI(N11277));
ADDFX1 inst_cellmath__203_0_I4043 (.CO(inst_cellmath__203__W0[19]), .S(inst_cellmath__203__W1[18]), .A(N12056), .B(N11856), .CI(N12597));
ADDFX1 inst_cellmath__203_0_I4044 (.CO(N12740), .S(N12389), .A(N11329), .B(N12674), .CI(N12030));
ADDFXL inst_cellmath__203_0_I4045 (.CO(N11782), .S(N11396), .A(N11521), .B(N11362), .CI(N12323));
ADDFX1 inst_cellmath__203_0_I4046 (.CO(N12538), .S(N12172), .A(N11217), .B(N12789), .CI(N12179));
ADDFX1 inst_cellmath__203_0_I4047 (.CO(N11558), .S(N11176), .A(N11823), .B(N12467), .CI(N12568));
ADDFX1 inst_cellmath__203_0_I4048 (.CO(N12327), .S(N11951), .A(N11396), .B(N12389), .CI(N11591));
ADDFX1 inst_cellmath__203_0_I4049 (.CO(N11335), .S(N12682), .A(N12360), .B(N12172), .CI(N11176));
ADDFXL inst_cellmath__203_0_I4050 (.CO(N12111), .S(N11716), .A(N11951), .B(N11364), .CI(N12595));
ADDFXL inst_cellmath__203_0_I4051 (.CO(N12829), .S(N12477), .A(N12145), .B(N12682), .CI(N11716));
ADDFXL inst_cellmath__203_0_I4052 (.CO(N11884), .S(N11495), .A(N11614), .B(N11429), .CI(N12864));
ADDFXL inst_cellmath__203_0_I4053 (.CO(N12623), .S(N12267), .A(N12297), .B(N12183), .CI(N12000));
ADDFX1 inst_cellmath__203_0_I4054 (.CO(N11652), .S(N11272), .A(N12365), .B(N11801), .CI(N12477));
ADDFX1 inst_cellmath__203_0_I4055 (.CO(N12418), .S(N12047), .A(N11922), .B(N12539), .CI(N12659));
ADDFXL inst_cellmath__203_0_I4056 (.CO(N11430), .S(N12768), .A(N11682), .B(N11495), .CI(N12267));
ADDFXL inst_cellmath__203_0_I4057 (.CO(N12204), .S(N11816), .A(N12449), .B(N11272), .CI(N11468));
ADDFHXL inst_cellmath__203_0_I4058 (.CO(N11203), .S(N12563), .A(N12047), .B(N12768), .CI(N12239));
ADDFHXL inst_cellmath__203_0_I4059 (.CO(inst_cellmath__203__W0[20]), .S(inst_cellmath__203__W1[19]), .A(N11816), .B(N11242), .CI(N12563));
INVXL inst_cellmath__203_0_I4060 (.Y(N12723), .A(N11743));
ADDFX1 inst_cellmath__203_0_I4061 (.CO(N12705), .S(N12352), .A(N11595), .B(N11748), .CI(N12723));
ADDFX1 inst_cellmath__203_0_I4062 (.CO(N12506), .S(N12138), .A(N12679), .B(N11910), .CI(N12542));
ADDFX1 inst_cellmath__203_0_I4063 (.CO(N11525), .S(N12859), .A(N11451), .B(N12402), .CI(N12819));
ADDFXL inst_cellmath__203_0_I4064 (.CO(N12293), .S(N11913), .A(N11782), .B(N12740), .CI(N12538));
ADDFX1 inst_cellmath__203_0_I4065 (.CO(N11301), .S(N12653), .A(N12859), .B(N12138), .CI(N12352));
ADDFXL inst_cellmath__203_0_I4066 (.CO(N12076), .S(N11675), .A(N11558), .B(N12327), .CI(N11913));
ADDFX1 inst_cellmath__203_0_I4067 (.CO(N12794), .S(N12443), .A(N12653), .B(N11631), .CI(N11335));
ADDFX1 inst_cellmath__203_0_I4068 (.CO(N11847), .S(N11463), .A(N12111), .B(N11675), .CI(N12443));
ADDFXL inst_cellmath__203_0_I4069 (.CO(N12591), .S(N12231), .A(N11811), .B(N12009), .CI(N12548));
ADDFXL inst_cellmath__203_0_I4070 (.CO(N11616), .S(N11236), .A(N12829), .B(N11303), .CI(N12374));
ADDFX1 inst_cellmath__203_0_I4071 (.CO(N12384), .S(N12014), .A(N12714), .B(N12191), .CI(N11178));
ADDFX1 inst_cellmath__203_0_I4072 (.CO(N11391), .S(N12732), .A(N11884), .B(N11463), .CI(N12623));
ADDFXL inst_cellmath__203_0_I4073 (.CO(N12164), .S(N11774), .A(N11652), .B(N12231), .CI(N11236));
ADDFX1 inst_cellmath__203_0_I4074 (.CO(N11169), .S(N12533), .A(N12418), .B(N12014), .CI(N11430));
ADDFXL cynw_cm_float_sin_I28147 (.CO(N43947), .S(N11551), .A(N11774), .B(N12732), .CI(N12204));
ADDFXL inst_cellmath__203_0_I4076 (.CO(inst_cellmath__203__W0[21]), .S(inst_cellmath__203__W1[20]), .A(N11203), .B(N12533), .CI(N11551));
INVXL inst_cellmath__203_0_I4077 (.Y(N12669), .A(N12469));
ADDFX1 inst_cellmath__203_0_I4078 (.CO(N11704), .S(N11328), .A(N11993), .B(N11743), .CI(N12669));
ADDFX1 inst_cellmath__203_0_I4079 (.CO(N11488), .S(N12822), .A(N11837), .B(N11333), .CI(N12292));
ADDFX1 inst_cellmath__203_0_I4080 (.CO(N12257), .S(N11873), .A(N11180), .B(N11485), .CI(N12752));
ADDFX1 inst_cellmath__203_0_I4081 (.CO(N11264), .S(N12616), .A(N12705), .B(N12143), .CI(N11525));
ADDFX1 inst_cellmath__203_0_I4082 (.CO(N12038), .S(N11642), .A(N12822), .B(N12506), .CI(N11873));
ADDFX1 inst_cellmath__203_0_I4083 (.CO(N12759), .S(N12410), .A(N12293), .B(N11328), .CI(N12616));
ADDFXL inst_cellmath__203_0_I4084 (.CO(N11805), .S(N11421), .A(N11642), .B(N11301), .CI(N12076));
ADDFX1 inst_cellmath__203_0_I4085 (.CO(N12558), .S(N12194), .A(N12794), .B(N12410), .CI(N12200));
ADDFXL inst_cellmath__203_0_I4086 (.CO(N11579), .S(N11197), .A(N12382), .B(N11421), .CI(N11184));
ADDFXL inst_cellmath__203_0_I4087 (.CO(N12346), .S(N11971), .A(N12078), .B(N12721), .CI(N12557));
ADDFX1 inst_cellmath__203_0_I4088 (.CO(N11354), .S(N12697), .A(N11368), .B(N11847), .CI(N11561));
ADDFX1 inst_cellmath__203_0_I4089 (.CO(N12130), .S(N11732), .A(N12591), .B(N12194), .CI(N11616));
ADDFX1 inst_cellmath__203_0_I4090 (.CO(N12851), .S(N12497), .A(N11971), .B(N11197), .CI(N12384));
ADDFXL inst_cellmath__203_0_I4094 (.CO(N12437), .S(N12068), .A(N11874), .B(N12469), .CI(N12224));
ADDFXL inst_cellmath__203_0_I4095 (.CO(N11453), .S(N12788), .A(N11563), .B(N11710), .CI(N12648));
ADDFX1 inst_cellmath__203_0_I4096 (.CO(N12223), .S(N11836), .A(N12368), .B(N11871), .CI(N12508));
ADDFX1 inst_cellmath__203_0_I4097 (.CO(N11227), .S(N12584), .A(N11704), .B(N11411), .CI(N12257));
ADDFX1 inst_cellmath__203_0_I4098 (.CO(N12004), .S(N11605), .A(N11488), .B(N12068), .CI(N12788));
ADDFX1 inst_cellmath__203_0_I4099 (.CO(N12725), .S(N12375), .A(N11264), .B(N11836), .CI(N12584));
ADDFX1 inst_cellmath__203_0_I4100 (.CO(N11765), .S(N11382), .A(N11605), .B(N12038), .CI(N12759));
ADDFXL inst_cellmath__203_0_I4101 (.CO(N12527), .S(N12158), .A(N12488), .B(N12375), .CI(N11805));
ADDFXL inst_cellmath__203_0_I4102 (.CO(N11544), .S(N11163), .A(N12731), .B(N11382), .CI(N11566));
ADDFXL inst_cellmath__203_0_I4103 (.CO(N12315), .S(N11934), .A(N11193), .B(N12797), .CI(N11378));
ADDFX1 inst_cellmath__203_0_I4104 (.CO(N11322), .S(N12670), .A(N12158), .B(N11754), .CI(N12558));
ADDFXL inst_cellmath__203_0_I4105 (.CO(N12096), .S(N11695), .A(N11955), .B(N11579), .CI(N12346));
ADDFX1 inst_cellmath__203_0_I4106 (.CO(N12815), .S(N12462), .A(N11354), .B(N11163), .CI(N11934));
INVXL inst_cellmath__203_0_I4110 (.Y(N12609), .A(N11410));
ADDFX1 inst_cellmath__203_0_I4111 (.CO(N12403), .S(N12029), .A(N12582), .B(N11957), .CI(N12609));
ADDFX1 inst_cellmath__203_0_I4112 (.CO(N12185), .S(N11795), .A(N11793), .B(N11298), .CI(N12254));
ADDFX1 inst_cellmath__203_0_I4113 (.CO(N11187), .S(N12551), .A(N12717), .B(N12862), .CI(N12108));
ADDFXL inst_cellmath__203_0_I4114 (.CO(N11962), .S(N11569), .A(N11453), .B(N12437), .CI(N12223));
ADDFX1 inst_cellmath__203_0_I4115 (.CO(N12692), .S(N12340), .A(N12029), .B(N11795), .CI(N12551));
ADDFXL inst_cellmath__203_0_I4116 (.CO(N11725), .S(N11346), .A(N11227), .B(N12004), .CI(N11569));
ADDFX1 inst_cellmath__203_0_I4117 (.CO(N12493), .S(N12124), .A(N12725), .B(N12340), .CI(N11346));
ADDFXL inst_cellmath__203_0_I4118 (.CO(N11508), .S(N12842), .A(N11387), .B(N11765), .CI(N12527));
ADDFX1 inst_cellmath__203_0_I4119 (.CO(N12281), .S(N11896), .A(N11960), .B(N11850), .CI(N12124));
ADDFX1 inst_cellmath__203_0_I4120 (.CO(N11283), .S(N12637), .A(N11576), .B(N11763), .CI(N12148));
ADDFXL inst_cellmath__203_0_I4121 (.CO(N12061), .S(N11659), .A(N11544), .B(N12329), .CI(N12315));
ADDFXL inst_cellmath__203_0_I4122 (.CO(N12779), .S(N12430), .A(N12842), .B(N11322), .CI(N11896));
INVXL inst_cellmath__203_0_I4126 (.Y(N12549), .A(N11373));
ADDFX1 inst_cellmath__203_0_I4127 (.CO(N12367), .S(N11994), .A(N11228), .B(N11410), .CI(N12549));
ADDFX1 inst_cellmath__203_0_I4128 (.CO(N12150), .S(N11756), .A(N11672), .B(N12186), .CI(N12614));
ADDFX1 inst_cellmath__203_0_I4129 (.CO(N12870), .S(N12519), .A(N12333), .B(N11529), .CI(N11371));
ADDFX1 inst_cellmath__203_0_I4130 (.CO(N11927), .S(N11535), .A(N12403), .B(N12475), .CI(N12185));
ADDFX1 inst_cellmath__203_0_I4131 (.CO(N12663), .S(N12308), .A(N11756), .B(N11187), .CI(N12519));
ADDFX1 inst_cellmath__203_0_I4132 (.CO(N11687), .S(N11314), .A(N11962), .B(N11994), .CI(N11535));
ADDFXL inst_cellmath__203_0_I4133 (.CO(N12455), .S(N12089), .A(N12308), .B(N12692), .CI(N11725));
ADDFXL inst_cellmath__203_0_I4134 (.CO(N11472), .S(N12807), .A(N11990), .B(N11314), .CI(N12089));
ADDFX1 inst_cellmath__203_0_I4135 (.CO(N12245), .S(N11859), .A(N12592), .B(N12493), .CI(N12338));
ADDFX1 inst_cellmath__203_0_I4136 (.CO(N11249), .S(N12601), .A(N12155), .B(N11969), .CI(N12515));
ADDFXL inst_cellmath__203_0_I4137 (.CO(N12024), .S(N11626), .A(N12807), .B(N11508), .CI(N12686));
ADDFX1 inst_cellmath__203_0_I4138 (.CO(N12745), .S(N12395), .A(N11283), .B(N12281), .CI(N11859));
ADDFX1 inst_cellmath__203_0_I4139 (.CO(N11788), .S(N11401), .A(N12061), .B(N12601), .CI(N11626));
ADDFXL cynw_cm_float_sin_I28154 (.CO(N11827), .S(N43935), .A(N12096), .B(N12637), .CI(N11659));
ADDFHXL inst_cellmath__203_0_I4140 (.CO(N12541), .S(N12178), .A(N12779), .B(N12395), .CI(N11827));
ADDFXL cynw_cm_float_sin_I28151 (.CO(N43997), .S(N43982), .A(N12670), .B(N12130), .CI(N11695));
ADDFHXL cynw_cm_float_sin_I28155 (.CO(N12574), .S(N43964), .A(N12815), .B(N12430), .CI(N43997));
ADDFHXL inst_cellmath__203_0_I4141 (.CO(inst_cellmath__203__W0[25]), .S(inst_cellmath__203__W1[24]), .A(N12574), .B(N11401), .CI(N12178));
XNOR2X1 inst_cellmath__203_0_I4142 (.Y(N11956), .A(N12411), .B(N11373));
OR2XL inst_cellmath__203_0_I4143 (.Y(N12334), .A(N12411), .B(N11373));
ADDFX1 inst_cellmath__203_0_I4144 (.CO(N12118), .S(N11721), .A(N11919), .B(N11956), .CI(N11262));
ADDFX1 inst_cellmath__203_0_I4145 (.CO(N12837), .S(N12483), .A(N12552), .B(N11606), .CI(N11757));
ADDFX1 inst_cellmath__203_0_I4146 (.CO(N11890), .S(N11500), .A(N12687), .B(N12825), .CI(N12072));
ADDFX1 inst_cellmath__203_0_I4147 (.CO(N12627), .S(N12274), .A(N12150), .B(N12367), .CI(N12870));
ADDFX1 inst_cellmath__203_0_I4148 (.CO(N11654), .S(N11275), .A(N12483), .B(N11721), .CI(N11500));
ADDFX1 inst_cellmath__203_0_I4149 (.CO(N12423), .S(N12053), .A(N11927), .B(N12663), .CI(N12274));
ADDFXL inst_cellmath__203_0_I4150 (.CO(N11434), .S(N12775), .A(N11687), .B(N11275), .CI(N12053));
ADDFX1 inst_cellmath__203_0_I4151 (.CO(N12209), .S(N11821), .A(N12455), .B(N11619), .CI(N12690));
ADDFX1 inst_cellmath__203_0_I4152 (.CO(N11207), .S(N12566), .A(N12775), .B(N12344), .CI(N12525));
ADDFXL inst_cellmath__203_0_I4153 (.CO(N11987), .S(N11589), .A(N11472), .B(N12868), .CI(N11337));
ADDFXL inst_cellmath__203_0_I4154 (.CO(N12710), .S(N12357), .A(N11249), .B(N12245), .CI(N11821));
ADDFX1 inst_cellmath__203_0_I4155 (.CO(N11747), .S(N11363), .A(N12024), .B(N12566), .CI(N11589));
ADDFXL inst_cellmath__203_0_I4156 (.CO(N12511), .S(N12142), .A(N12357), .B(N12745), .CI(N11788));
ADDFXL inst_cellmath__203_0_I4157 (.CO(inst_cellmath__203__W0[26]), .S(inst_cellmath__203__W1[25]), .A(N12541), .B(N11363), .CI(N12142));
ADDHX1 inst_cellmath__203_0_I4158 (.CO(N12299), .S(N11920), .A(N12334), .B(N12001));
ADDFX1 inst_cellmath__203_0_I4159 (.CO(N11306), .S(N12657), .A(N11188), .B(N12151), .CI(N11920));
ADDFX1 inst_cellmath__203_0_I4160 (.CO(N12082), .S(N11679), .A(N11493), .B(N11638), .CI(N12300));
ADDFX1 inst_cellmath__203_0_I4161 (.CO(N12798), .S(N12448), .A(N12441), .B(N11339), .CI(N12118));
ADDFHXL inst_cellmath__203_0_I4162 (.CO(N11854), .S(N11466), .A(N12837), .B(N11890), .CI(N12657));
ADDFX1 inst_cellmath__203_0_I4163 (.CO(N12596), .S(N12236), .A(N12627), .B(N11679), .CI(N12448));
ADDFX1 inst_cellmath__203_0_I4164 (.CO(N11621), .S(N11239), .A(N11466), .B(N11654), .CI(N12236));
ADDFX1 inst_cellmath__203_0_I4165 (.CO(N12388), .S(N12018), .A(N12451), .B(N12423), .CI(N11434));
ADDFX1 inst_cellmath__203_0_I4166 (.CO(N11395), .S(N12736), .A(N12386), .B(N11239), .CI(N11344));
ADDFXL inst_cellmath__203_0_I4167 (.CO(N12170), .S(N11780), .A(N11161), .B(N11531), .CI(N11718));
ADDFX1 inst_cellmath__203_0_I4168 (.CO(N11174), .S(N12536), .A(N12209), .B(N12018), .CI(N11207));
ADDFX1 inst_cellmath__203_0_I4169 (.CO(N11948), .S(N11556), .A(N11987), .B(N12736), .CI(N11780));
ADDFXL inst_cellmath__203_0_I4170 (.CO(N12678), .S(N12326), .A(N12536), .B(N12710), .CI(N11747));
ADDFXL inst_cellmath__203_0_I4171 (.CO(inst_cellmath__203__W0[27]), .S(inst_cellmath__203__W1[26]), .A(N12511), .B(N11556), .CI(N12326));
XNOR2X1 inst_cellmath__203_0_I4172 (.Y(N12107), .A(N12376), .B(N11881));
OR2XL inst_cellmath__203_0_I4173 (.Y(N12474), .A(N12376), .B(N11881));
ADDFX1 inst_cellmath__203_0_I4174 (.CO(N12265), .S(N11880), .A(N12518), .B(N11570), .CI(N11720));
ADDFX1 inst_cellmath__203_0_I4175 (.CO(N11268), .S(N12619), .A(N12792), .B(N12299), .CI(N12658));
ADDFX1 inst_cellmath__203_0_I4176 (.CO(N12043), .S(N11649), .A(N12035), .B(N12107), .CI(N11306));
ADDFX1 inst_cellmath__203_0_I4177 (.CO(N12765), .S(N12415), .A(N11880), .B(N12082), .CI(N12619));
ADDFXL inst_cellmath__203_0_I4178 (.CO(N11812), .S(N11427), .A(N11854), .B(N12798), .CI(N11649));
ADDFXL inst_cellmath__203_0_I4179 (.CO(N12561), .S(N12202), .A(N12415), .B(N12596), .CI(N11427));
ADDFX1 inst_cellmath__203_0_I4180 (.CO(N11584), .S(N11201), .A(N11393), .B(N11621), .CI(N11723));
ADDFXL inst_cellmath__203_0_I4181 (.CO(N12351), .S(N11977), .A(N11541), .B(N12202), .CI(N11924));
ADDFX1 inst_cellmath__203_0_I4182 (.CO(N11360), .S(N12703), .A(N12115), .B(N12388), .CI(N11395));
ADDFX1 inst_cellmath__203_0_I4183 (.CO(N12136), .S(N11740), .A(N12170), .B(N11201), .CI(N11977));
ADDFXL inst_cellmath__203_0_I4184 (.CO(N12857), .S(N12502), .A(N12703), .B(N11174), .CI(N11948));
ADDFXL inst_cellmath__203_0_I4185 (.CO(inst_cellmath__203__W0[28]), .S(inst_cellmath__203__W1[27]), .A(N12678), .B(N11740), .CI(N12502));
INVXL inst_cellmath__203_0_I4186 (.Y(N11826), .A(N11668));
ADDFX1 inst_cellmath__203_0_I4187 (.CO(N12650), .S(N12291), .A(N12871), .B(N11963), .CI(N11826));
ADDFX1 inst_cellmath__203_0_I4188 (.CO(N12440), .S(N12075), .A(N11460), .B(N12119), .CI(N12262));
ADDFX1 inst_cellmath__203_0_I4189 (.CO(N11459), .S(N12791), .A(N12408), .B(N11304), .CI(N12474));
ADDFX1 inst_cellmath__203_0_I4190 (.CO(N12228), .S(N11843), .A(N11268), .B(N12265), .CI(N12075));
ADDFXL inst_cellmath__203_0_I4191 (.CO(N11235), .S(N12588), .A(N12791), .B(N12291), .CI(N12043));
ADDFXL inst_cellmath__203_0_I4192 (.CO(N12011), .S(N11612), .A(N11843), .B(N12765), .CI(N12588));
ADDFX1 inst_cellmath__203_0_I4193 (.CO(N12729), .S(N12383), .A(N11177), .B(N11812), .CI(N11612));
ADDFX1 inst_cellmath__203_0_I4194 (.CO(N11772), .S(N11388), .A(N12168), .B(N12561), .CI(N12122));
ADDFXL inst_cellmath__203_0_I4195 (.CO(N12530), .S(N12162), .A(N12481), .B(N12306), .CI(N12383));
ADDFX1 inst_cellmath__203_0_I4196 (.CO(N11549), .S(N11168), .A(N12351), .B(N11584), .CI(N11388));
ADDFXL inst_cellmath__203_0_I4197 (.CO(N12318), .S(N11939), .A(N12162), .B(N11360), .CI(N12136));
ADDFXL inst_cellmath__203_0_I4198 (.CO(inst_cellmath__203__W0[29]), .S(inst_cellmath__203__W1[28]), .A(N12857), .B(N11168), .CI(N11939));
ADDFX1 inst_cellmath__203_0_I4199 (.CO(N12100), .S(N11702), .A(N12341), .B(N11668), .CI(N11844));
ADDFX1 inst_cellmath__203_0_I4200 (.CO(N12821), .S(N12466), .A(N12484), .B(N11536), .CI(N11680));
ADDFX1 inst_cellmath__203_0_I4201 (.CO(N11870), .S(N11484), .A(N12620), .B(N12756), .CI(N12650));
ADDFX1 inst_cellmath__203_0_I4202 (.CO(N12613), .S(N12256), .A(N11702), .B(N12440), .CI(N11459));
ADDFX1 inst_cellmath__203_0_I4203 (.CO(N11640), .S(N11261), .A(N11484), .B(N12466), .CI(N12228));
ADDFX1 inst_cellmath__203_0_I4204 (.CO(N12407), .S(N12034), .A(N11235), .B(N12256), .CI(N11261));
ADDFXL inst_cellmath__203_0_I4205 (.CO(N11417), .S(N12758), .A(N11172), .B(N12011), .CI(N12491));
ADDFX1 inst_cellmath__203_0_I4206 (.CO(N12192), .S(N11802), .A(N12729), .B(N12034), .CI(N12660));
ADDFX1 inst_cellmath__203_0_I4207 (.CO(N11194), .S(N12555), .A(N11772), .B(N12831), .CI(N12758));
ADDFX1 inst_cellmath__203_0_I4208 (.CO(N11967), .S(N11577), .A(N12530), .B(N11802), .CI(N11549));
ADDFX1 inst_cellmath__203_0_I4209 (.CO(inst_cellmath__203__W0[30]), .S(inst_cellmath__203__W1[29]), .A(N12318), .B(N12555), .CI(N11577));
INVXL inst_cellmath__203_0_I4210 (.Y(N11755), .A(N11413));
ADDFX1 inst_cellmath__203_0_I4211 (.CO(N11729), .S(N11351), .A(N12834), .B(N11926), .CI(N11755));
ADDFX1 inst_cellmath__203_0_I4212 (.CO(N11512), .S(N12849), .A(N11418), .B(N12083), .CI(N12229));
ADDFX1 inst_cellmath__203_0_I4213 (.CO(N12284), .S(N11901), .A(N12100), .B(N11269), .CI(N12821));
ADDFX1 inst_cellmath__203_0_I4214 (.CO(N11289), .S(N12642), .A(N11351), .B(N12849), .CI(N11870));
ADDFX1 inst_cellmath__203_0_I4215 (.CO(N12065), .S(N11664), .A(N11901), .B(N12613), .CI(N12642));
ADDFX1 inst_cellmath__203_0_I4216 (.CO(N12785), .S(N12435), .A(N11664), .B(N11640), .CI(N12769));
ADDFX1 inst_cellmath__203_0_I4217 (.CO(N11833), .S(N11449), .A(N11945), .B(N12407), .CI(N11310));
ADDFX1 inst_cellmath__203_0_I4218 (.CO(N12581), .S(N12221), .A(N11499), .B(N12435), .CI(N11417));
ADDFX1 inst_cellmath__203_0_I4219 (.CO(N11602), .S(N11224), .A(N11449), .B(N12192), .CI(N11194));
ADDFX1 inst_cellmath__203_0_I4220 (.CO(inst_cellmath__203__W0[31]), .S(inst_cellmath__203__W1[30]), .A(N11967), .B(N12221), .CI(N11224));
ADDFX1 inst_cellmath__203_0_I4221 (.CO(N11379), .S(N12722), .A(N12309), .B(N11413), .CI(N11803));
ADDFX1 inst_cellmath__203_0_I4222 (.CO(N12156), .S(N11762), .A(N12446), .B(N11501), .CI(N11647));
ADDFX1 inst_cellmath__203_0_I4223 (.CO(N11160), .S(N12526), .A(N11729), .B(N12589), .CI(N11512));
ADDFX1 inst_cellmath__203_0_I4224 (.CO(N11932), .S(N11542), .A(N11762), .B(N12722), .CI(N12284));
ADDFX1 inst_cellmath__203_0_I4225 (.CO(N12668), .S(N12314), .A(N11289), .B(N12526), .CI(N11542));
ADDFX1 inst_cellmath__203_0_I4226 (.CO(N11692), .S(N11319), .A(N12314), .B(N12065), .CI(N12677));
ADDFX1 inst_cellmath__203_0_I4227 (.CO(N12460), .S(N12094), .A(N11685), .B(N12785), .CI(N11888));
ADDFX1 inst_cellmath__203_0_I4228 (.CO(N11476), .S(N12813), .A(N11319), .B(N11833), .CI(N12581));
ADDFX1 inst_cellmath__203_0_I4229 (.CO(inst_cellmath__203__W0[32]), .S(inst_cellmath__203__W1[31]), .A(N11602), .B(N12094), .CI(N12813));
INVXL inst_cellmath__203_0_I4230 (.Y(N11686), .A(N12576));
ADDFX1 inst_cellmath__203_0_I4231 (.CO(N11254), .S(N12607), .A(N12799), .B(N11891), .CI(N11686));
ADDFX1 inst_cellmath__203_0_I4232 (.CO(N12751), .S(N12401), .A(N12190), .B(N12044), .CI(N11233));
ADDFX1 inst_cellmath__203_0_I4233 (.CO(N11792), .S(N11407), .A(N12156), .B(N11379), .CI(N12607));
ADDFX1 inst_cellmath__203_0_I4234 (.CO(N12547), .S(N12184), .A(N11160), .B(N12401), .CI(N11932));
ADDFX1 inst_cellmath__203_0_I4235 (.CO(N11568), .S(N11185), .A(N12668), .B(N11407), .CI(N12184));
ADDFXL inst_cellmath__203_0_I4236 (.CO(N12339), .S(N11959), .A(N11708), .B(N11915), .CI(N11185));
ADDFXL inst_cellmath__203_0_I4237 (.CO(N11342), .S(N12691), .A(N11692), .B(N12269), .CI(N11959));
ADDFX1 inst_cellmath__203_0_I4238 (.CO(inst_cellmath__203__W1[33]), .S(inst_cellmath__203__W1[32]), .A(N12691), .B(N12460), .CI(N11476));
ADDFX1 inst_cellmath__203_0_I4239 (.CO(N12840), .S(N12489), .A(N12273), .B(N12576), .CI(N11467));
ADDFX1 inst_cellmath__203_0_I4240 (.CO(N11894), .S(N11506), .A(N11613), .B(N12416), .CI(N12556));
ADDFX1 inst_cellmath__203_0_I4241 (.CO(N12634), .S(N12280), .A(N12751), .B(N11254), .CI(N12489));
ADDFX1 inst_cellmath__203_0_I4242 (.CO(N11657), .S(N11280), .A(N11792), .B(N11506), .CI(N12280));
ADDFX1 inst_cellmath__203_0_I4243 (.CO(N12427), .S(N12059), .A(N11280), .B(N12547), .CI(N11568));
ADDFX1 inst_cellmath__203_0_I4244 (.CO(N11441), .S(N12777), .A(N12626), .B(N12471), .CI(N12059));
ADDFX1 inst_cellmath__203_0_I4245 (.CO(inst_cellmath__203__W1[34]), .S(inst_cellmath__203__W0[33]), .A(N12777), .B(N12339), .CI(N11342));
INVXL inst_cellmath__203_0_I4246 (.Y(N11625), .A(N12747));
ADDFX1 inst_cellmath__203_0_I4247 (.CO(N11214), .S(N12571), .A(N12763), .B(N11852), .CI(N11625));
ADDFX1 inst_cellmath__203_0_I4248 (.CO(N12715), .S(N12363), .A(N11195), .B(N12012), .CI(N12840));
ADDFX1 inst_cellmath__203_0_I4249 (.CO(N11752), .S(N11370), .A(N12571), .B(N11894), .CI(N12634));
ADDFX1 inst_cellmath__203_0_I4250 (.CO(N12516), .S(N12149), .A(N11657), .B(N12363), .CI(N11370));
ADDFX1 inst_cellmath__203_0_I4251 (.CO(N11532), .S(N12866), .A(N11492), .B(N12149), .CI(N12734));
ADDFX1 inst_cellmath__203_0_I4252 (.CO(inst_cellmath__203__W1[35]), .S(inst_cellmath__203__W0[34]), .A(N12866), .B(N12427), .CI(N11441));
ADDFX1 inst_cellmath__203_0_I4253 (.CO(N11312), .S(N12661), .A(N12237), .B(N12747), .CI(N11428));
ADDFX1 inst_cellmath__203_0_I4254 (.CO(N12087), .S(N11683), .A(N11575), .B(N12381), .CI(N11214));
ADDFX1 inst_cellmath__203_0_I4255 (.CO(N12805), .S(N12453), .A(N12715), .B(N12661), .CI(N11683));
ADDFX1 inst_cellmath__203_0_I4256 (.CO(N11858), .S(N11470), .A(N12453), .B(N11752), .CI(N12516));
ADDFX1 inst_cellmath__203_0_I4257 (.CO(inst_cellmath__203__W1[36]), .S(inst_cellmath__203__W0[35]), .A(N11470), .B(N12260), .CI(N11532));
INVXL inst_cellmath__203_0_I4258 (.Y(N11562), .A(N11210));
ADDFX1 inst_cellmath__203_0_I4259 (.CO(N11623), .S(N11246), .A(N12730), .B(N11813), .CI(N11562));
ADDFX1 inst_cellmath__203_0_I4260 (.CO(N11398), .S(N12742), .A(N11312), .B(N11968), .CI(N11246));
ADDFX1 inst_cellmath__203_0_I4261 (.CO(N12174), .S(N11785), .A(N12742), .B(N12087), .CI(N12805));
ADDFX1 inst_cellmath__203_0_I4262 (.CO(inst_cellmath__203__W1[37]), .S(inst_cellmath__203__W0[36]), .A(N12749), .B(N11785), .CI(N11858));
ADDFX1 inst_cellmath__203_0_I4263 (.CO(N11953), .S(N11559), .A(N12199), .B(N11210), .CI(N11389));
ADDFX1 inst_cellmath__203_0_I4264 (.CO(N12684), .S(N12330), .A(N11623), .B(N12345), .CI(N11559));
ADDFX1 inst_cellmath__203_0_I4265 (.CO(inst_cellmath__203__W1[38]), .S(inst_cellmath__203__W0[37]), .A(N12330), .B(N11398), .CI(N12174));
ADDFX1 inst_cellmath__203_0_I4266 (.CO(N12479), .S(N12116), .A(N11771), .B(N11240), .CI(N12695));
ADDFX1 inst_cellmath__203_0_I4267 (.CO(inst_cellmath__203__W1[39]), .S(inst_cellmath__203__W0[38]), .A(N12116), .B(N11953), .CI(N12684));
INVXL inst_cellmath__203_0_I4268 (.Y(N11886), .A(N12270));
ADDFX1 inst_cellmath__203_0_I4269 (.CO(inst_cellmath__203__W1[40]), .S(inst_cellmath__203__W0[39]), .A(N11352), .B(N11886), .CI(N12479));
ADDFX1 inst_cellmath__203_0_I4270 (.CO(inst_cellmath__203__W1[41]), .S(inst_cellmath__203__W0[40]), .A(N12270), .B(N11270), .CI(N11730));
INVXL inst_cellmath__203_0_I4271 (.Y(inst_cellmath__203__W0[41]), .A(inst_cellmath__203__W1[42]));
ADDHX1 cynw_cm_float_sin_I4274 (.CO(N14718), .S(N14599), .A(inst_cellmath__203__W0[18]), .B(inst_cellmath__195[0]));
ADDFHXL cynw_cm_float_sin_I4275 (.CO(N14970), .S(N14845), .A(inst_cellmath__203__W0[19]), .B(inst_cellmath__195[1]), .CI(inst_cellmath__203__W1[19]));
ADDFXL cynw_cm_float_sin_I4276 (.CO(N14650), .S(N14520), .A(inst_cellmath__195[2]), .B(inst_cellmath__203__W0[20]), .CI(inst_cellmath__203__W1[20]));
ADDFXL cynw_cm_float_sin_I28148 (.CO(N43976), .S(N43960), .A(N12697), .B(N11391), .CI(N12164));
ADDFHXL cynw_cm_float_sin_I28149 (.CO(N43938), .S(N43990), .A(N11732), .B(N12497), .CI(N11169));
ADDFHXL cynw_cm_float_sin_I28150 (.CO(N43967), .S(inst_cellmath__203__W1[21]), .A(N43947), .B(N43960), .CI(N43990));
ADDFHXL cynw_cm_float_sin_I4277 (.CO(N14895), .S(N14772), .A(inst_cellmath__195[3]), .B(inst_cellmath__203__W0[21]), .CI(inst_cellmath__203__W1[21]));
ADDFXL cynw_cm_float_sin_I28152 (.CO(N43957), .S(N43944), .A(N12462), .B(N12851), .CI(N43976));
ADDFHXL cynw_cm_float_sin_I28156 (.CO(inst_cellmath__203__W0[24]), .S(N43994), .A(N43935), .B(N43957), .CI(N43964));
ADDFHXL cynw_cm_float_sin_I4280 (.CO(N15074), .S(N14948), .A(inst_cellmath__195[6]), .B(inst_cellmath__203__W0[24]), .CI(inst_cellmath__203__W1[24]));
ADDFHX1 cynw_cm_float_sin_I4281 (.CO(N14749), .S(N14628), .A(inst_cellmath__195[7]), .B(inst_cellmath__203__W0[25]), .CI(inst_cellmath__203__W1[25]));
ADDFXL cynw_cm_float_sin_I4282 (.CO(N14998), .S(N14874), .A(inst_cellmath__203__W0[26]), .B(inst_cellmath__195[8]), .CI(inst_cellmath__203__W1[26]));
ADDFHX1 cynw_cm_float_sin_I4283 (.CO(N14682), .S(N14554), .A(inst_cellmath__203__W0[27]), .B(inst_cellmath__195[9]), .CI(inst_cellmath__203__W1[27]));
ADDFXL cynw_cm_float_sin_I4284 (.CO(N14927), .S(N14801), .A(inst_cellmath__203__W0[28]), .B(inst_cellmath__195[10]), .CI(inst_cellmath__203__W1[28]));
ADDFHXL cynw_cm_float_sin_I4285 (.CO(N14607), .S(N15058), .A(inst_cellmath__203__W0[29]), .B(inst_cellmath__195[11]), .CI(inst_cellmath__203__W1[29]));
ADDFX1 cynw_cm_float_sin_I4286 (.CO(N14855), .S(N14728), .A(inst_cellmath__203__W0[30]), .B(inst_cellmath__195[12]), .CI(inst_cellmath__203__W1[30]));
ADDFX1 cynw_cm_float_sin_I4287 (.CO(N14535), .S(N14978), .A(inst_cellmath__203__W0[31]), .B(inst_cellmath__195[13]), .CI(inst_cellmath__203__W1[31]));
ADDFX1 cynw_cm_float_sin_I4288 (.CO(N14779), .S(N14661), .A(inst_cellmath__195[14]), .B(inst_cellmath__203__W0[32]), .CI(inst_cellmath__203__W1[32]));
ADDFX1 cynw_cm_float_sin_I4289 (.CO(N15034), .S(N14909), .A(inst_cellmath__203__W1[33]), .B(inst_cellmath__195[15]), .CI(inst_cellmath__203__W0[33]));
ADDFX1 cynw_cm_float_sin_I4290 (.CO(N14710), .S(N14586), .A(inst_cellmath__203__W0[34]), .B(inst_cellmath__195[16]), .CI(inst_cellmath__203__W1[34]));
ADDFX1 cynw_cm_float_sin_I4291 (.CO(N14956), .S(N14836), .A(inst_cellmath__203__W1[35]), .B(inst_cellmath__195[17]), .CI(inst_cellmath__203__W0[35]));
ADDFX1 cynw_cm_float_sin_I4292 (.CO(N14640), .S(N15087), .A(inst_cellmath__203__W0[36]), .B(inst_cellmath__195[18]), .CI(inst_cellmath__203__W1[36]));
ADDFX1 cynw_cm_float_sin_I4293 (.CO(N14885), .S(N14758), .A(inst_cellmath__203__W0[37]), .B(inst_cellmath__195[19]), .CI(inst_cellmath__203__W1[37]));
ADDFX1 cynw_cm_float_sin_I4294 (.CO(N14562), .S(N15011), .A(inst_cellmath__203__W0[38]), .B(inst_cellmath__195[20]), .CI(inst_cellmath__203__W1[38]));
ADDFX1 cynw_cm_float_sin_I4295 (.CO(N14813), .S(N14692), .A(inst_cellmath__203__W0[39]), .B(inst_cellmath__195[21]), .CI(inst_cellmath__203__W1[39]));
ADDFX1 cynw_cm_float_sin_I4296 (.CO(N15066), .S(N14934), .A(inst_cellmath__203__W0[40]), .B(inst_cellmath__195[22]), .CI(inst_cellmath__203__W1[40]));
ADDFX1 cynw_cm_float_sin_I4297 (.CO(N14736), .S(N14616), .A(inst_cellmath__203__W0[41]), .B(inst_cellmath__195[23]), .CI(inst_cellmath__203__W1[41]));
ADDFX1 cynw_cm_float_sin_I4298 (.CO(N14987), .S(N14865), .A(inst_cellmath__203__W1[42]), .B(inst_cellmath__203__W0[42]), .CI(inst_cellmath__195[24]));
ADDHX1 cynw_cm_float_sin_I4299 (.CO(N14671), .S(N14541), .A(1'B1), .B(inst_cellmath__195[25]));
ADDHX1 cynw_cm_float_sin_I4300 (.CO(N14914), .S(N14788), .A(1'B1), .B(inst_cellmath__195[26]));
ADDHX1 cynw_cm_float_sin_I4301 (.CO(N14596), .S(N15043), .A(1'B1), .B(inst_cellmath__195[27]));
INVXL hap1_A_I28351 (.Y(N14716), .A(inst_cellmath__195[28]));
OR2XL hap1_A_I10792 (.Y(N14843), .A(1'B0), .B(inst_cellmath__195[28]));
INVXL cynw_cm_float_sin_I4303 (.Y(N14966), .A(inst_cellmath__195[29]));
NOR2XL cynw_cm_float_sin_I4307 (.Y(N14697), .A(N11504), .B(inst_cellmath__203__W1[2]));
NOR2XL cynw_cm_float_sin_I4309 (.Y(N14944), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
NAND2XL cynw_cm_float_sin_I4310 (.Y(N15072), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
NOR2XL cynw_cm_float_sin_I4311 (.Y(N14625), .A(inst_cellmath__203__W0[4]), .B(inst_cellmath__203__W1[4]));
NAND2XL cynw_cm_float_sin_I4312 (.Y(N14745), .A(inst_cellmath__203__W0[4]), .B(inst_cellmath__203__W1[4]));
NOR2XL cynw_cm_float_sin_I4313 (.Y(N14871), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
NOR2XL cynw_cm_float_sin_I4315 (.Y(N14551), .A(inst_cellmath__203__W0[6]), .B(inst_cellmath__203__W1[6]));
NAND2X1 cynw_cm_float_sin_I4316 (.Y(N14679), .A(inst_cellmath__203__W0[6]), .B(inst_cellmath__203__W1[6]));
NOR2XL cynw_cm_float_sin_I4317 (.Y(N14797), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
NAND2XL cynw_cm_float_sin_I4318 (.Y(N14924), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
OR2XL cynw_cm_float_sin_I4319 (.Y(N15055), .A(inst_cellmath__203__W0[8]), .B(inst_cellmath__203__W1[8]));
AND2XL cynw_cm_float_sin_I4320 (.Y(N14604), .A(inst_cellmath__203__W0[8]), .B(inst_cellmath__203__W1[8]));
NOR2XL cynw_cm_float_sin_I4321 (.Y(N14724), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
NAND2XL cynw_cm_float_sin_I4322 (.Y(N14853), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
NOR2XL cynw_cm_float_sin_I4323 (.Y(N14974), .A(inst_cellmath__203__W0[10]), .B(inst_cellmath__203__W1[10]));
NAND2X1 cynw_cm_float_sin_I4324 (.Y(N14530), .A(inst_cellmath__203__W0[10]), .B(inst_cellmath__203__W1[10]));
OR2XL cynw_cm_float_sin_I4325 (.Y(N14658), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
AND2XL cynw_cm_float_sin_I4326 (.Y(N14777), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
NOR2XL cynw_cm_float_sin_I4327 (.Y(N14904), .A(inst_cellmath__203__W0[12]), .B(inst_cellmath__203__W1[12]));
NAND2XL cynw_cm_float_sin_I4328 (.Y(N15031), .A(inst_cellmath__203__W0[12]), .B(inst_cellmath__203__W1[12]));
NOR2XL cynw_cm_float_sin_I4329 (.Y(N14582), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NAND2X1 cynw_cm_float_sin_I4330 (.Y(N14707), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NOR2XL cynw_cm_float_sin_I4331 (.Y(N14834), .A(inst_cellmath__203__W0[14]), .B(inst_cellmath__203__W1[14]));
NOR2XL cynw_cm_float_sin_I4333 (.Y(N15083), .A(inst_cellmath__203__W0[15]), .B(inst_cellmath__203__W1[15]));
NAND2X1 cynw_cm_float_sin_I4334 (.Y(N14638), .A(inst_cellmath__203__W0[15]), .B(inst_cellmath__203__W1[15]));
NOR2XL cynw_cm_float_sin_I4335 (.Y(N14756), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
NAND2XL cynw_cm_float_sin_I4336 (.Y(N14882), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
AND2XL cynw_cm_float_sin_I28352 (.Y(N14690), .A(inst_cellmath__203__W0[1]), .B(inst_cellmath__203__W1[1]));
AOI21XL cynw_cm_float_sin_I4338 (.Y(N14615), .A0(N15072), .A1(N14697), .B0(N14944));
OAI2BB1X1 cynw_cm_float_sin_I10151 (.Y(N14733), .A0N(N11504), .A1N(inst_cellmath__203__W1[2]), .B0(N15072));
OAI21XL cynw_cm_float_sin_I4340 (.Y(N15041), .A0(N14733), .A1(N14690), .B0(N14615));
AOI21XL cynw_cm_float_sin_I4341 (.Y(N14572), .A0(N14745), .A1(N15041), .B0(N14625));
AOI21XL cynw_cm_float_sin_I4342 (.Y(N15069), .A0(N14679), .A1(N14871), .B0(N14551));
OAI2BB1X1 cynw_cm_float_sin_I10569 (.Y(N14623), .A0N(inst_cellmath__203__W0[5]), .A1N(inst_cellmath__203__W1[5]), .B0(N14679));
OAI21XL cynw_cm_float_sin_I4344 (.Y(N14529), .A0(N14623), .A1(N14572), .B0(N15069));
AOI21X1 cynw_cm_float_sin_I4345 (.Y(N14807), .A0(N14924), .A1(N14529), .B0(N14797));
OAI21X1 cynw_cm_float_sin_I4348 (.Y(N15016), .A0(N14604), .A1(N14807), .B0(N15055));
AOI21XL cynw_cm_float_sin_I4349 (.Y(N14940), .A0(N14530), .A1(N14724), .B0(N14974));
INVXL cynw_cm_float_sin_I4350 (.Y(N14763), .A(N14940));
AND2XL cynw_cm_float_sin_I4351 (.Y(N14887), .A(N14530), .B(N14853));
AOI21X1 cynw_cm_float_sin_I4353 (.Y(N14751), .A0(N14887), .A1(N15016), .B0(N14763));
OAI21X2 cynw_cm_float_sin_I4356 (.Y(N14565), .A0(N14777), .A1(N14751), .B0(N14658));
AO21XL cynw_cm_float_sin_I4357 (.Y(N15075), .A0(N14707), .A1(N14904), .B0(N14582));
AND2XL cynw_cm_float_sin_I4358 (.Y(N14627), .A(N15031), .B(N14707));
AOI21X2 cynw_cm_float_sin_I4360 (.Y(N15057), .A0(N14627), .A1(N14565), .B0(N15075));
AOI21X1 cynw_cm_float_sin_I4362 (.Y(N14977), .A0(N14638), .A1(N14834), .B0(N15083));
OAI2BB1X1 cynw_cm_float_sin_I10157 (.Y(N14534), .A0N(inst_cellmath__203__W0[14]), .A1N(inst_cellmath__203__W1[14]), .B0(N14638));
OAI21X2 cynw_cm_float_sin_I4364 (.Y(N14965), .A0(N14534), .A1(N15057), .B0(N14977));
AOI21X2 cynw_cm_float_sin_I4371 (.Y(N14635), .A0(N14882), .A1(N14965), .B0(N14756));
INVX1 cynw_cm_float_sin_I4405 (.Y(N14621), .A(N14635));
NOR2XL cynw_cm_float_sin_I4406 (.Y(N14867), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
NAND2XL cynw_cm_float_sin_I4407 (.Y(N14992), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
NOR2XL cynw_cm_float_sin_I4408 (.Y(N14545), .A(N14599), .B(inst_cellmath__203__W1[18]));
NAND2XL cynw_cm_float_sin_I4409 (.Y(N14673), .A(N14599), .B(inst_cellmath__203__W1[18]));
NOR2XL cynw_cm_float_sin_I4410 (.Y(N14792), .A(N14718), .B(N14845));
NAND2X2 cynw_cm_float_sin_I4411 (.Y(N14918), .A(N14718), .B(N14845));
NOR2X2 cynw_cm_float_sin_I4412 (.Y(N15048), .A(N14970), .B(N14520));
NAND2X1 cynw_cm_float_sin_I4413 (.Y(N14601), .A(N14970), .B(N14520));
NOR2X1 cynw_cm_float_sin_I4414 (.Y(N14719), .A(N14650), .B(N14772));
NAND2X4 cynw_cm_float_sin_I4415 (.Y(N14847), .A(N14650), .B(N14772));
NOR4X1 cynw_cm_float_sin_I28363 (.Y(N43963), .A(N7697), .B(N7931), .C(N8393), .D(N8230));
NOR4BBX1 cynw_cm_float_sin_I28139 (.Y(N43949), .AN(N8037), .BN(N8307), .C(N7934), .D(N8734));
NAND4XL cynw_cm_float_sin_I28364 (.Y(N43993), .A(N8727), .B(N8531), .C(N43963), .D(N43949));
ADDFXL cynw_cm_float_sin_I28153 (.CO(N43987), .S(N43973), .A(N43938), .B(N43982), .CI(N43944));
ADDFHXL cynw_cm_float_sin_I28157 (.CO(N14577), .S(N15022), .A(N43967), .B(N43993), .CI(N43973));
NOR2X2 cynw_cm_float_sin_I4416 (.Y(N14971), .A(N14895), .B(N15022));
NAND2X1 cynw_cm_float_sin_I4417 (.Y(N14522), .A(N14895), .B(N15022));
OR2XL cynw_cm_float_sin_I28365 (.Y(N43970), .A(N8397), .B(N8145));
NAND3XL hyperpropagate_4_1_A_I28634 (.Y(N44116), .A(N8638), .B(N8360), .C(N8554));
NOR2XL hyperpropagate_4_1_A_I28635 (.Y(N43954), .A(N7760), .B(N44116));
NOR2XL cynw_cm_float_sin_I28143 (.Y(N43941), .A(N8301), .B(N7882));
NAND4BXL cynw_cm_float_sin_I28146 (.Y(N43985), .AN(N43970), .B(N43954), .C(N8215), .D(N43941));
ADDFHXL cynw_cm_float_sin_I28158 (.CO(N14823), .S(N14699), .A(N43987), .B(N43985), .CI(N43994));
NOR2X1 cynw_cm_float_sin_I4418 (.Y(N14651), .A(N14577), .B(N14699));
NAND2X4 cynw_cm_float_sin_I28159 (.Y(N14773), .A(N14577), .B(N14699));
NOR2X2 cynw_cm_float_sin_I4420 (.Y(N14897), .A(N14823), .B(N14948));
NAND2X1 cynw_cm_float_sin_I4421 (.Y(N15023), .A(N14823), .B(N14948));
NOR2X1 cynw_cm_float_sin_I4422 (.Y(N14578), .A(N15074), .B(N14628));
NAND2X4 cynw_cm_float_sin_I4423 (.Y(N14701), .A(N15074), .B(N14628));
NOR2X1 cynw_cm_float_sin_I4424 (.Y(N14824), .A(N14749), .B(N14874));
NAND2X1 cynw_cm_float_sin_I4425 (.Y(N14949), .A(N14749), .B(N14874));
NOR2X1 cynw_cm_float_sin_I4426 (.Y(N15076), .A(N14998), .B(N14554));
NAND2X4 cynw_cm_float_sin_I4427 (.Y(N14629), .A(N14998), .B(N14554));
NOR2X1 cynw_cm_float_sin_I4428 (.Y(N14750), .A(N14682), .B(N14801));
NAND2X1 cynw_cm_float_sin_I4429 (.Y(N14875), .A(N14682), .B(N14801));
NOR2XL cynw_cm_float_sin_I4430 (.Y(N14999), .A(N14927), .B(N15058));
NAND2X2 cynw_cm_float_sin_I4431 (.Y(N14556), .A(N14927), .B(N15058));
NOR2XL cynw_cm_float_sin_I4432 (.Y(N14683), .A(N14607), .B(N14728));
NAND2XL cynw_cm_float_sin_I4433 (.Y(N14802), .A(N14607), .B(N14728));
NOR2XL cynw_cm_float_sin_I4434 (.Y(N14928), .A(N14855), .B(N14978));
NAND2X1 cynw_cm_float_sin_I4435 (.Y(N15059), .A(N14855), .B(N14978));
NOR2XL cynw_cm_float_sin_I4436 (.Y(N14608), .A(N14535), .B(N14661));
NAND2XL cynw_cm_float_sin_I4437 (.Y(N14729), .A(N14535), .B(N14661));
NOR2XL cynw_cm_float_sin_I4438 (.Y(N14856), .A(N14909), .B(N14779));
NAND2XL cynw_cm_float_sin_I4439 (.Y(N14979), .A(N14909), .B(N14779));
NOR2XL cynw_cm_float_sin_I4440 (.Y(N14536), .A(N14586), .B(N15034));
NAND2XL cynw_cm_float_sin_I4441 (.Y(N14663), .A(N14586), .B(N15034));
NOR2XL cynw_cm_float_sin_I4442 (.Y(N14780), .A(N14710), .B(N14836));
NAND2XL cynw_cm_float_sin_I4443 (.Y(N14910), .A(N14710), .B(N14836));
NOR2XL cynw_cm_float_sin_I4444 (.Y(N15036), .A(N15087), .B(N14956));
NAND2XL cynw_cm_float_sin_I4445 (.Y(N14587), .A(N15087), .B(N14956));
NOR2XL cynw_cm_float_sin_I4446 (.Y(N14711), .A(N14758), .B(N14640));
NAND2XL cynw_cm_float_sin_I4447 (.Y(N14838), .A(N14758), .B(N14640));
NOR2XL cynw_cm_float_sin_I4448 (.Y(N14957), .A(N15011), .B(N14885));
NAND2XL cynw_cm_float_sin_I4449 (.Y(N15088), .A(N15011), .B(N14885));
NOR2XL cynw_cm_float_sin_I4450 (.Y(N14641), .A(N14692), .B(N14562));
NAND2XL cynw_cm_float_sin_I4451 (.Y(N14759), .A(N14692), .B(N14562));
NOR2XL cynw_cm_float_sin_I4452 (.Y(N14886), .A(N14934), .B(N14813));
NAND2XL cynw_cm_float_sin_I4453 (.Y(N15012), .A(N14934), .B(N14813));
NOR2XL cynw_cm_float_sin_I4454 (.Y(N14563), .A(N14616), .B(N15066));
NAND2XL cynw_cm_float_sin_I4455 (.Y(N14693), .A(N14616), .B(N15066));
NOR2XL cynw_cm_float_sin_I4456 (.Y(N14814), .A(N14865), .B(N14736));
NAND2XL cynw_cm_float_sin_I4457 (.Y(N14935), .A(N14865), .B(N14736));
NOR2XL cynw_cm_float_sin_I4458 (.Y(N15067), .A(N14987), .B(N14541));
NAND2XL cynw_cm_float_sin_I4459 (.Y(N14617), .A(N14987), .B(N14541));
NOR2XL cynw_cm_float_sin_I4460 (.Y(N14737), .A(N14671), .B(N14788));
NAND2XL cynw_cm_float_sin_I4461 (.Y(N14866), .A(N14671), .B(N14788));
NOR2XL cynw_cm_float_sin_I4462 (.Y(N14988), .A(N14914), .B(N15043));
NAND2XL cynw_cm_float_sin_I4463 (.Y(N14542), .A(N14914), .B(N15043));
NOR2XL cynw_cm_float_sin_I4464 (.Y(N14672), .A(N14596), .B(N14716));
NAND2XL cynw_cm_float_sin_I4465 (.Y(N14789), .A(N14596), .B(N14716));
NOR2XL cynw_cm_float_sin_I4466 (.Y(N14915), .A(N14966), .B(N14843));
NAND2XL cynw_cm_float_sin_I4467 (.Y(N15045), .A(N14966), .B(N14843));
AOI21X2 cynw_cm_float_sin_I4468 (.Y(N14967), .A0(N14992), .A1(N14621), .B0(N14867));
AOI21X2 cynw_cm_float_sin_I4469 (.Y(N14893), .A0(N14918), .A1(N14545), .B0(N14792));
NAND2X1 cynw_cm_float_sin_I4470 (.Y(N15020), .A(N14673), .B(N14918));
AOI21X4 cynw_cm_float_sin_I4471 (.Y(N14821), .A0(N15048), .A1(N14847), .B0(N14719));
NAND2X2 cynw_cm_float_sin_I4472 (.Y(N14945), .A(N14601), .B(N14847));
AOI21X4 cynw_cm_float_sin_I4473 (.Y(N14746), .A0(N14971), .A1(N14773), .B0(N14651));
NAND2X4 cynw_cm_float_sin_I4474 (.Y(N14872), .A(N14522), .B(N14773));
AOI21X4 cynw_cm_float_sin_I4475 (.Y(N14680), .A0(N14701), .A1(N14897), .B0(N14578));
NAND2X2 cynw_cm_float_sin_I4476 (.Y(N14799), .A(N14701), .B(N15023));
AOI21X2 cynw_cm_float_sin_I4477 (.Y(N14605), .A0(N14629), .A1(N14824), .B0(N15076));
NAND2X4 cynw_cm_float_sin_I4478 (.Y(N14725), .A(N14629), .B(N14949));
AOI21X1 cynw_cm_float_sin_I4479 (.Y(N14531), .A0(N14556), .A1(N14750), .B0(N14999));
NAND2X2 cynw_cm_float_sin_I4480 (.Y(N14660), .A(N14556), .B(N14875));
AOI21XL cynw_cm_float_sin_I4481 (.Y(N15033), .A0(N15059), .A1(N14683), .B0(N14928));
NAND2X1 cynw_cm_float_sin_I4482 (.Y(N14583), .A(N15059), .B(N14802));
AOI21XL cynw_cm_float_sin_I4483 (.Y(N14954), .A0(N14979), .A1(N14608), .B0(N14856));
NAND2X1 cynw_cm_float_sin_I4484 (.Y(N15084), .A(N14979), .B(N14729));
AOI21XL cynw_cm_float_sin_I4485 (.Y(N14883), .A0(N14910), .A1(N14536), .B0(N14780));
NAND2XL cynw_cm_float_sin_I4486 (.Y(N15010), .A(N14910), .B(N14663));
INVXL cynw_cm_float_sin_I4487 (.Y(N14975), .A(N14587));
AOI21XL cynw_cm_float_sin_I4488 (.Y(N14812), .A0(N14838), .A1(N15036), .B0(N14711));
NAND2XL cynw_cm_float_sin_I4489 (.Y(N14931), .A(N14838), .B(N14587));
AOI21XL cynw_cm_float_sin_I4490 (.Y(N14595), .A0(N14759), .A1(N14957), .B0(N14641));
NAND2XL cynw_cm_float_sin_I4491 (.Y(N14714), .A(N14759), .B(N15088));
INVXL cynw_cm_float_sin_I4492 (.Y(N14832), .A(N15012));
AOI21XL cynw_cm_float_sin_I4493 (.Y(N14515), .A0(N14693), .A1(N14886), .B0(N14563));
NAND2XL cynw_cm_float_sin_I4494 (.Y(N14646), .A(N14693), .B(N15012));
AOI21XL cynw_cm_float_sin_I4495 (.Y(N14869), .A0(N14617), .A1(N14814), .B0(N15067));
NAND2XL cynw_cm_float_sin_I4496 (.Y(N14994), .A(N14617), .B(N14935));
INVXL cynw_cm_float_sin_I4497 (.Y(N14689), .A(N14866));
AOI21XL cynw_cm_float_sin_I4498 (.Y(N14795), .A0(N14542), .A1(N14737), .B0(N14988));
NAND2XL cynw_cm_float_sin_I4499 (.Y(N14923), .A(N14542), .B(N14866));
AOI21XL cynw_cm_float_sin_I4500 (.Y(N14580), .A0(N15045), .A1(N14672), .B0(N14915));
NAND2XL cynw_cm_float_sin_I4501 (.Y(N14706), .A(N15045), .B(N14789));
INVXL cynw_cm_float_sin_I4502 (.Y(N14985), .A(N14966));
NOR2X1 cynw_cm_float_sin_I4503 (.Y(N15006), .A(N14580), .B(N14985));
NOR2XL cynw_cm_float_sin_I4504 (.Y(N14557), .A(N14975), .B(N14883));
NOR2XL cynw_cm_float_sin_I4505 (.Y(N14963), .A(N14557), .B(N15036));
OA21X1 cynw_cm_float_sin_I4506 (.Y(N14645), .A0(N14931), .A1(N14883), .B0(N14812));
OR2XL cynw_cm_float_sin_I4507 (.Y(N14767), .A(N14931), .B(N15010));
NOR2XL cynw_cm_float_sin_I4508 (.Y(N14858), .A(N14832), .B(N14595));
NOR2XL cynw_cm_float_sin_I4509 (.Y(N14817), .A(N14858), .B(N14886));
OA21X1 cynw_cm_float_sin_I4510 (.Y(N15070), .A0(N14646), .A1(N14595), .B0(N14515));
OR2XL cynw_cm_float_sin_I4511 (.Y(N14622), .A(N14646), .B(N14714));
NOR2XL cynw_cm_float_sin_I4512 (.Y(N14588), .A(N14689), .B(N14869));
OA21X1 cynw_cm_float_sin_I4514 (.Y(N14922), .A0(N14923), .A1(N14869), .B0(N14795));
OR2XL cynw_cm_float_sin_I4515 (.Y(N15052), .A(N14923), .B(N14994));
OR2XL cynw_cm_float_sin_I4516 (.Y(N14655), .A(N14985), .B(N14706));
INVXL cynw_cm_float_sin_I4517 (.Y(N14775), .A(N14967));
OAI21X2 cynw_cm_float_sin_I4518 (.Y(N14794), .A0(N15020), .A1(N14967), .B0(N14893));
OAI21X1 cynw_cm_float_sin_I4519 (.Y(N15050), .A0(N14945), .A1(N14893), .B0(N14821));
NOR2XL cynw_cm_float_sin_I4520 (.Y(N14602), .A(N15020), .B(N14945));
OAI21X4 cynw_cm_float_sin_I4521 (.Y(N14722), .A0(N14872), .A1(N14821), .B0(N14746));
NOR2X2 cynw_cm_float_sin_I4522 (.Y(N14849), .A(N14945), .B(N14872));
OAI21X2 cynw_cm_float_sin_I4523 (.Y(N14972), .A0(N14799), .A1(N14746), .B0(N14680));
NOR2X2 cynw_cm_float_sin_I4524 (.Y(N14526), .A(N14799), .B(N14872));
OAI21X4 cynw_cm_float_sin_I4525 (.Y(N14653), .A0(N14725), .A1(N14680), .B0(N14605));
NOR2X2 cynw_cm_float_sin_I4526 (.Y(N14774), .A(N14725), .B(N14799));
OAI21X1 cynw_cm_float_sin_I4527 (.Y(N14900), .A0(N14660), .A1(N14605), .B0(N14531));
NOR2XL cynw_cm_float_sin_I4528 (.Y(N15025), .A(N14660), .B(N14725));
OAI21X1 cynw_cm_float_sin_I4529 (.Y(N14579), .A0(N14583), .A1(N14531), .B0(N15033));
NOR2X1 cynw_cm_float_sin_I4530 (.Y(N14704), .A(N14583), .B(N14660));
OAI21XL cynw_cm_float_sin_I4531 (.Y(N14827), .A0(N15084), .A1(N15033), .B0(N14954));
NOR2XL cynw_cm_float_sin_I4532 (.Y(N14950), .A(N15084), .B(N14583));
OAI21XL cynw_cm_float_sin_I4533 (.Y(N15080), .A0(N14767), .A1(N14954), .B0(N14645));
NOR2XL cynw_cm_float_sin_I4534 (.Y(N14631), .A(N14767), .B(N15084));
OAI21XL cynw_cm_float_sin_I4535 (.Y(N14752), .A0(N14622), .A1(N14645), .B0(N15070));
NOR2XL cynw_cm_float_sin_I4536 (.Y(N14878), .A(N14622), .B(N14767));
OAI21XL cynw_cm_float_sin_I4537 (.Y(N15001), .A0(N15052), .A1(N15070), .B0(N14922));
NOR2XL cynw_cm_float_sin_I4538 (.Y(N14558), .A(N15052), .B(N14622));
INVXL cynw_cm_float_sin_I4539 (.Y(N14902), .A(N14775));
INVXL cynw_cm_float_sin_I4540 (.Y(N15028), .A(N14794));
AOI21XL cynw_cm_float_sin_I4541 (.Y(N14610), .A0(N14602), .A1(N14775), .B0(N15050));
AOI21X2 cynw_cm_float_sin_I4542 (.Y(N14861), .A0(N14849), .A1(N14794), .B0(N14722));
AOI21X2 cynw_cm_float_sin_I4543 (.Y(N14537), .A0(N14526), .A1(N15050), .B0(N14972));
NAND2X1 cynw_cm_float_sin_I4544 (.Y(N14666), .A(N14526), .B(N14602));
AOI21X2 cynw_cm_float_sin_I4545 (.Y(N14783), .A0(N14774), .A1(N14722), .B0(N14653));
NAND2XL cynw_cm_float_sin_I4546 (.Y(N14911), .A(N14774), .B(N14849));
AOI21XL cynw_cm_float_sin_I4547 (.Y(N15039), .A0(N15025), .A1(N14972), .B0(N14900));
NAND2XL cynw_cm_float_sin_I4548 (.Y(N14590), .A(N15025), .B(N14526));
AOI21X2 cynw_cm_float_sin_I4549 (.Y(N14712), .A0(N14704), .A1(N14653), .B0(N14579));
NAND2X2 cynw_cm_float_sin_I4550 (.Y(N14841), .A(N14704), .B(N14774));
AOI21X1 cynw_cm_float_sin_I4551 (.Y(N14959), .A0(N14950), .A1(N14900), .B0(N14827));
NAND2X1 cynw_cm_float_sin_I4552 (.Y(N15089), .A(N15025), .B(N14950));
AOI21X1 cynw_cm_float_sin_I4553 (.Y(N14644), .A0(N14631), .A1(N14579), .B0(N15080));
NAND2XL cynw_cm_float_sin_I4554 (.Y(N14761), .A(N14631), .B(N14704));
AOI21X1 cynw_cm_float_sin_I4555 (.Y(N14888), .A0(N14878), .A1(N14827), .B0(N14752));
NAND2XL cynw_cm_float_sin_I4556 (.Y(N15015), .A(N14878), .B(N14950));
AOI21X1 cynw_cm_float_sin_I4557 (.Y(N14566), .A0(N14558), .A1(N15080), .B0(N15001));
NAND2X1 cynw_cm_float_sin_I4558 (.Y(N14694), .A(N14631), .B(N14558));
INVXL cynw_cm_float_sin_I4559 (.Y(N14830), .A(N14902));
INVXL cynw_cm_float_sin_I4560 (.Y(N14951), .A(N15028));
INVX2 cynw_cm_float_sin_I4562 (.Y(N14634), .A(N14861));
OAI21X2 cynw_cm_float_sin_I4563 (.Y(N14521), .A0(N15089), .A1(N14537), .B0(N14959));
NOR2X1 cynw_cm_float_sin_I4564 (.Y(N14649), .A(N14666), .B(N15089));
OAI21X1 cynw_cm_float_sin_I4565 (.Y(N14771), .A0(N14761), .A1(N14783), .B0(N14644));
NOR2X1 cynw_cm_float_sin_I4566 (.Y(N14896), .A(N14761), .B(N14911));
OAI21X2 cynw_cm_float_sin_I4569 (.Y(N14700), .A0(N14694), .A1(N14712), .B0(N14566));
NOR2X2 cynw_cm_float_sin_I4570 (.Y(N14822), .A(N14694), .B(N14841));
INVXL cynw_cm_float_sin_I10793 (.Y(N22732), .A(N14634));
OA21X1 cynw_cm_float_sin_I4575 (.Y(N14687), .A0(N14902), .A1(N14666), .B0(N14537));
OA21X1 cynw_cm_float_sin_I4576 (.Y(N14808), .A0(N14911), .A1(N15028), .B0(N14783));
OA21X1 cynw_cm_float_sin_I4577 (.Y(N14929), .A0(N14590), .A1(N14610), .B0(N15039));
OA21X1 cynw_cm_float_sin_I4578 (.Y(N15063), .A0(N14841), .A1(N14861), .B0(N14712));
AOI21X2 cynw_cm_float_sin_I4580 (.Y(N14908), .A0(N14896), .A1(N14951), .B0(N14771));
AOI21X2 cynw_cm_float_sin_I4582 (.Y(N14837), .A0(N14822), .A1(N14634), .B0(N14700));
NAND2BXL cynw_cm_float_sin_I4593 (.Y(N14810), .AN(N14578), .B(N14701));
NAND2BXL cynw_cm_float_sin_I4594 (.Y(N14614), .AN(N14824), .B(N14949));
NAND2BXL cynw_cm_float_sin_I4595 (.Y(N14986), .AN(N15076), .B(N14629));
NAND2BXL cynw_cm_float_sin_I4596 (.Y(N14787), .AN(N14750), .B(N14875));
NAND2BXL cynw_cm_float_sin_I4597 (.Y(N14594), .AN(N14999), .B(N14556));
NAND2BXL cynw_cm_float_sin_I4598 (.Y(N14964), .AN(N14683), .B(N14802));
NAND2BXL cynw_cm_float_sin_I4599 (.Y(N14768), .AN(N14928), .B(N15059));
NAND2BXL cynw_cm_float_sin_I4600 (.Y(N14571), .AN(N14608), .B(N14729));
NAND2BXL cynw_cm_float_sin_I4601 (.Y(N14943), .AN(N14856), .B(N14979));
NAND2BXL cynw_cm_float_sin_I4603 (.Y(N14550), .AN(N14780), .B(N14910));
NAND2BXL cynw_cm_float_sin_I4604 (.Y(N15003), .AN(N15036), .B(N14587));
NAND2BXL cynw_cm_float_sin_I4605 (.Y(N14667), .AN(N14711), .B(N14838));
NAND2BXL cynw_cm_float_sin_I4606 (.Y(N14528), .AN(N14957), .B(N15088));
NAND2BXL cynw_cm_float_sin_I4607 (.Y(N14903), .AN(N14641), .B(N14759));
NAND2BXL cynw_cm_float_sin_I4608 (.Y(N14620), .AN(N14886), .B(N15012));
NAND2BXL cynw_cm_float_sin_I4609 (.Y(N14846), .AN(N14563), .B(N14693));
NAND2BXL cynw_cm_float_sin_I4610 (.Y(N14881), .AN(N14814), .B(N14935));
NAND2BXL cynw_cm_float_sin_I4611 (.Y(N14688), .AN(N15067), .B(N14617));
NAND2BXL cynw_cm_float_sin_I4612 (.Y(N14803), .AN(N14737), .B(N14866));
NAND2BXL cynw_cm_float_sin_I4614 (.Y(N14669), .AN(N14672), .B(N14789));
NAND2BXL cynw_cm_float_sin_I4615 (.Y(N15040), .AN(N14915), .B(N15045));
XNOR2XL cynw_cm_float_sin_I4621 (.Y(inst_cellmath__201[26]), .A(N14614), .B(N14687));
XOR2XL cynw_cm_float_sin_I4622 (.Y(inst_cellmath__201[28]), .A(N14787), .B(N14808));
XOR2XL cynw_cm_float_sin_I4623 (.Y(inst_cellmath__201[30]), .A(N14964), .B(N14929));
XOR2XL cynw_cm_float_sin_I4624 (.Y(inst_cellmath__201[32]), .A(N14571), .B(N15063));
XOR2XL cynw_cm_float_sin_I4626 (.Y(inst_cellmath__201[38]), .A(N14528), .B(N14908));
NOR2X1 inst_cellmath__200_0_I27962 (.Y(N43441), .A(N15015), .B(N14590));
INVXL inst_cellmath__200_0_I27960 (.Y(N43426), .A(N14610));
OAI21X1 inst_cellmath__200_0_I27961 (.Y(N43433), .A0(N15015), .A1(N15039), .B0(N14888));
AOI21X2 inst_cellmath__200_0_I27963 (.Y(N14585), .A0(N43441), .A1(N43426), .B0(N43433));
XOR2XL cynw_cm_float_sin_I4627 (.Y(inst_cellmath__201[42]), .A(N14585), .B(N14881));
XOR2XL cynw_cm_float_sin_I4628 (.Y(inst_cellmath__201[46]), .A(N14837), .B(N14669));
XNOR2X1 cynw_cm_float_sin_I4638 (.Y(N14652), .A(N15023), .B(N14810));
XNOR2X1 cynw_cm_float_sin_I4639 (.Y(N14525), .A(N14897), .B(N14810));
MXI2XL cynw_cm_float_sin_I28375 (.Y(inst_cellmath__201[25]), .A(N14652), .B(N14525), .S0(N22732));
XNOR2X1 cynw_cm_float_sin_I4641 (.Y(N15024), .A(N14949), .B(N14986));
XNOR2X1 cynw_cm_float_sin_I4642 (.Y(N14899), .A(N14824), .B(N14986));
MXI2XL cynw_cm_float_sin_I4643 (.Y(inst_cellmath__201[27]), .A(N15024), .B(N14899), .S0(N14687));
XNOR2X1 cynw_cm_float_sin_I4644 (.Y(N14826), .A(N14594), .B(N14875));
XNOR2X1 cynw_cm_float_sin_I4645 (.Y(N14703), .A(N14594), .B(N14750));
MX2XL cynw_cm_float_sin_I4646 (.Y(inst_cellmath__201[29]), .A(N14826), .B(N14703), .S0(N14808));
XNOR2X1 cynw_cm_float_sin_I4647 (.Y(N14630), .A(N14768), .B(N14802));
XNOR2X1 cynw_cm_float_sin_I4648 (.Y(N15079), .A(N14768), .B(N14683));
MX2XL cynw_cm_float_sin_I4649 (.Y(inst_cellmath__201[31]), .A(N14630), .B(N15079), .S0(N14929));
XNOR2X1 cynw_cm_float_sin_I4650 (.Y(N15000), .A(N14943), .B(N14729));
XNOR2X1 cynw_cm_float_sin_I4651 (.Y(N14877), .A(N14943), .B(N14608));
MX2XL cynw_cm_float_sin_I4652 (.Y(inst_cellmath__201[33]), .A(N15000), .B(N14877), .S0(N15063));
XOR2XL cynw_cm_float_sin_I4656 (.Y(N15061), .A(N15003), .B(N14883));
NAND2XL cynw_cm_float_sin_I4657 (.Y(N14753), .A(N15010), .B(N14883));
XNOR2X1 cynw_cm_float_sin_I4658 (.Y(N14609), .A(N15003), .B(N14753));
AOI21X2 inst_cellmath__200_0_I28105 (.Y(N14662), .A0(N14649), .A1(N14830), .B0(N14521));
MX2XL cynw_cm_float_sin_I4659 (.Y(inst_cellmath__201[36]), .A(N14609), .B(N15061), .S0(N14662));
XOR2XL cynw_cm_float_sin_I4660 (.Y(N14859), .A(N14667), .B(N14963));
OAI21XL cynw_cm_float_sin_I4661 (.Y(N14982), .A0(N14975), .A1(N15010), .B0(N14963));
XNOR2X1 cynw_cm_float_sin_I4662 (.Y(N14980), .A(N14667), .B(N14982));
MXI2XL mx2a_A_I28636 (.Y(N44122), .A(N14980), .B(N14859), .S0(N14662));
INVXL mx2a_A_I28637 (.Y(inst_cellmath__201[37]), .A(N44122));
XNOR2X1 cynw_cm_float_sin_I4664 (.Y(N14782), .A(N14903), .B(N15088));
XNOR2X1 cynw_cm_float_sin_I4665 (.Y(N14665), .A(N14903), .B(N14957));
MXI2XL cynw_cm_float_sin_I4666 (.Y(inst_cellmath__201[39]), .A(N14782), .B(N14665), .S0(N14908));
XOR2XL cynw_cm_float_sin_I4667 (.Y(N15038), .A(N14620), .B(N14595));
NAND2XL cynw_cm_float_sin_I4668 (.Y(N14938), .A(N14714), .B(N14595));
XNOR2X1 cynw_cm_float_sin_I4669 (.Y(N14589), .A(N14620), .B(N14938));
MXI2XL cynw_cm_float_sin_I4670 (.Y(inst_cellmath__201[40]), .A(N14589), .B(N15038), .S0(N14908));
XOR2XL cynw_cm_float_sin_I4671 (.Y(N14840), .A(N14846), .B(N14817));
OAI21XL cynw_cm_float_sin_I4672 (.Y(N14600), .A0(N14832), .A1(N14714), .B0(N14817));
XNOR2X1 cynw_cm_float_sin_I4673 (.Y(N14958), .A(N14846), .B(N14600));
MXI2XL cynw_cm_float_sin_I4674 (.Y(inst_cellmath__201[41]), .A(N14958), .B(N14840), .S0(N14908));
XNOR2X1 cynw_cm_float_sin_I4675 (.Y(N14760), .A(N14688), .B(N14935));
XNOR2X1 cynw_cm_float_sin_I4676 (.Y(N14643), .A(N14688), .B(N14814));
MXI2XL cynw_cm_float_sin_I4677 (.Y(inst_cellmath__201[43]), .A(N14760), .B(N14643), .S0(N14585));
XOR2XL cynw_cm_float_sin_I4678 (.Y(N15014), .A(N14803), .B(N14869));
NAND2XL cynw_cm_float_sin_I4679 (.Y(N14555), .A(N14994), .B(N14869));
XNOR2X1 cynw_cm_float_sin_I4680 (.Y(N14564), .A(N14803), .B(N14555));
MX2XL cynw_cm_float_sin_I4681 (.Y(inst_cellmath__201[44]), .A(N14564), .B(N15014), .S0(N14585));
XNOR2X1 cynw_cm_float_sin_I4686 (.Y(N14739), .A(N15040), .B(N14789));
XNOR2X1 cynw_cm_float_sin_I4687 (.Y(N14619), .A(N15040), .B(N14672));
MX2XL cynw_cm_float_sin_I4688 (.Y(inst_cellmath__201[47]), .A(N14739), .B(N14619), .S0(N14837));
XOR2XL cynw_cm_float_sin_I4689 (.Y(N14990), .A(N14985), .B(N14580));
NAND2XL cynw_cm_float_sin_I4690 (.Y(N14738), .A(N14706), .B(N14580));
XNOR2X1 cynw_cm_float_sin_I4691 (.Y(N14543), .A(N14985), .B(N14738));
MXI2XL cynw_cm_float_sin_I4692 (.Y(inst_cellmath__201[48]), .A(N14543), .B(N14990), .S0(N14837));
NOR2XL inst_cellmath__200_0_I27959 (.Y(N43449), .A(N14737), .B(N14588));
NAND2BXL inst_cellmath__200_0_I27964 (.Y(N43424), .AN(N14988), .B(N14542));
XNOR2X1 inst_cellmath__200_0_I28376 (.Y(N43432), .A(N43449), .B(N43424));
OAI21XL inst_cellmath__200_0_I27967 (.Y(N43438), .A0(N14689), .A1(N14994), .B0(N43449));
XOR2XL inst_cellmath__200_0_I28377 (.Y(N43446), .A(N43424), .B(N43438));
INVX1 inst_cellmath__200_0_I27970 (.Y(N43434), .A(N14585));
NAND2BXL inst_cellmath__200_0_I28106 (.Y(N43811), .AN(N14536), .B(N14663));
XOR2XL inst_cellmath__200_0_I28107 (.Y(N43817), .A(N43811), .B(N14662));
XNOR2X1 inst_cellmath__200_0_I28108 (.Y(N43800), .A(N14550), .B(N14663));
XNOR2X1 inst_cellmath__200_0_I28109 (.Y(N43804), .A(N14536), .B(N14550));
MX2XL inst_cellmath__200_0_I28110 (.Y(N43808), .A(N43800), .B(N43804), .S0(N14662));
AOI2BB1X4 inst_cellmath__200_0_I28111 (.Y(N43813), .A0N(N14655), .A1N(N14837), .B0(N15006));
INVX12 inst_cellmath__200_0_I28112 (.Y(N22595), .A(N43813));
NOR2X1 inst_cellmath__200_0_I28113 (.Y(inst_cellmath__210[9]), .A(N22595), .B(N43817));
NOR2X1 inst_cellmath__200_0_I28114 (.Y(inst_cellmath__210[10]), .A(N22595), .B(N43808));
NOR2X2 inst_cellmath__200_0_I28115 (.Y(N15984), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[9]));
MXI2X1 inst_cellmath__200_0_I27972 (.Y(N43448), .A(N43432), .B(N43446), .S0(N43434));
NOR2X2 inst_cellmath__200_0_I27973 (.Y(inst_cellmath__210[20]), .A(N22595), .B(N43448));
NOR2BX1 inst_cellmath__200_0_I4743 (.Y(inst_cellmath__210[0]), .AN(inst_cellmath__201[25]), .B(N22595));
NOR2BX1 inst_cellmath__200_0_I4744 (.Y(inst_cellmath__210[1]), .AN(inst_cellmath__201[26]), .B(N22595));
NOR2BX1 inst_cellmath__200_0_I4745 (.Y(inst_cellmath__210[2]), .AN(inst_cellmath__201[27]), .B(N22595));
NOR2X2 inst_cellmath__200_0_I4746 (.Y(inst_cellmath__210[3]), .A(inst_cellmath__201[28]), .B(N22595));
NOR2X2 inst_cellmath__200_0_I4747 (.Y(inst_cellmath__210[4]), .A(inst_cellmath__201[29]), .B(N22595));
NOR2X1 inst_cellmath__200_0_I4748 (.Y(inst_cellmath__210[5]), .A(inst_cellmath__201[30]), .B(N22595));
NOR2X2 inst_cellmath__200_0_I4749 (.Y(inst_cellmath__210[6]), .A(N22595), .B(inst_cellmath__201[31]));
NOR2X2 inst_cellmath__200_0_I4750 (.Y(inst_cellmath__210[7]), .A(inst_cellmath__201[32]), .B(N22595));
NOR2X1 inst_cellmath__200_0_I4751 (.Y(inst_cellmath__210[8]), .A(inst_cellmath__201[33]), .B(N22595));
NOR2X2 inst_cellmath__200_0_I4754 (.Y(inst_cellmath__210[11]), .A(N22595), .B(inst_cellmath__201[36]));
NOR2X2 inst_cellmath__200_0_I4755 (.Y(inst_cellmath__210[12]), .A(N22595), .B(inst_cellmath__201[37]));
NOR2X2 inst_cellmath__200_0_I4756 (.Y(inst_cellmath__210[13]), .A(N22595), .B(inst_cellmath__201[38]));
NOR2BX2 inst_cellmath__200_0_I4757 (.Y(inst_cellmath__210[14]), .AN(inst_cellmath__201[39]), .B(N22595));
NOR2BX1 inst_cellmath__200_0_I4758 (.Y(inst_cellmath__210[15]), .AN(inst_cellmath__201[40]), .B(N22595));
NOR2BXL inst_cellmath__200_0_I4759 (.Y(inst_cellmath__210[16]), .AN(inst_cellmath__201[41]), .B(N22595));
NOR2X1 inst_cellmath__200_0_I4760 (.Y(inst_cellmath__210[17]), .A(N22595), .B(inst_cellmath__201[42]));
NOR2BX1 inst_cellmath__200_0_I4761 (.Y(inst_cellmath__210[18]), .AN(inst_cellmath__201[43]), .B(N22595));
NOR2X1 inst_cellmath__200_0_I4762 (.Y(inst_cellmath__210[19]), .A(N22595), .B(inst_cellmath__201[44]));
NOR2X1 inst_cellmath__200_0_I4764 (.Y(inst_cellmath__210[21]), .A(inst_cellmath__201[46]), .B(N22595));
NOR2XL inst_cellmath__200_0_I4765 (.Y(inst_cellmath__210[22]), .A(inst_cellmath__201[47]), .B(N22595));
NAND2XL inst_cellmath__19_0_I4768 (.Y(N15746), .A(a_exp[6]), .B(a_exp[5]));
NAND2XL inst_cellmath__19_0_I4769 (.Y(N15749), .A(a_exp[4]), .B(a_exp[3]));
NAND2XL inst_cellmath__19_0_I4770 (.Y(N15737), .A(a_exp[2]), .B(a_exp[1]));
NOR2XL inst_cellmath__19_0_I4772 (.Y(N15744), .A(N15749), .B(N15737));
NAND3XL hyperpropagate_4_1_A_I10795 (.Y(N22738), .A(a_exp[7]), .B(a_exp[0]), .C(N15744));
NOR2XL hyperpropagate_4_1_A_I10796 (.Y(inst_cellmath__19), .A(N15746), .B(N22738));
NOR2XL inst_cellmath__24_0_I4774 (.Y(N15790), .A(a_man[0]), .B(a_man[1]));
NOR2XL inst_cellmath__24_0_I4776 (.Y(N15763), .A(a_man[20]), .B(a_man[19]));
NOR2XL inst_cellmath__24_0_I4777 (.Y(N15773), .A(a_man[18]), .B(a_man[17]));
NOR2XL inst_cellmath__24_0_I4778 (.Y(N15784), .A(a_man[16]), .B(a_man[15]));
NOR2XL inst_cellmath__24_0_I4779 (.Y(N15794), .A(a_man[14]), .B(a_man[13]));
NOR2XL inst_cellmath__24_0_I4780 (.Y(N15804), .A(a_man[12]), .B(a_man[11]));
NOR2XL inst_cellmath__24_0_I4781 (.Y(N15767), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__24_0_I4782 (.Y(N15777), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__24_0_I4783 (.Y(N15788), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__24_0_I4784 (.Y(N15798), .A(a_man[4]), .B(a_man[3]));
NAND2XL inst_cellmath__24_0_I4786 (.Y(N15771), .A(N5956), .B(N15790));
AND4XL inst_cellmath__24_0_I28385 (.Y(N15796), .A(N15804), .B(N15773), .C(N15784), .D(N15794));
NAND3XL hyperpropagate_4_1_A_I10797 (.Y(N22746), .A(N6053), .B(N15763), .C(N15796));
NOR2XL hyperpropagate_4_1_A_I10798 (.Y(N15769), .A(N15771), .B(N22746));
AND4XL inst_cellmath__24_0_I28387 (.Y(N15780), .A(N15798), .B(N15767), .C(N15777), .D(N15788));
NAND2XL inst_cellmath__24_0_I4796 (.Y(inst_cellmath__24), .A(N15780), .B(N15769));
INVXL inst_cellmath__66_0_I4797 (.Y(N15829), .A(a_sign));
NAND2XL inst_cellmath__66_0_I4798 (.Y(N15832), .A(N15829), .B(inst_cellmath__19));
NAND2XL cynw_cm_float_sin_I4800 (.Y(N15839), .A(a_sign), .B(inst_cellmath__19));
AOI21XL cynw_cm_float_sin_I28389 (.Y(inst_cellmath__68), .A0(N15839), .A1(N15832), .B0(inst_cellmath__24));
INVXL inst_cellmath__82_0_I10172 (.Y(N15854), .A(inst_cellmath__19));
INVXL inst_cellmath__82_0_I4806 (.Y(inst_cellmath__82), .A(N15854));
OR4X1 inst_cellmath__17_0_I28390 (.Y(N15863), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 inst_cellmath__17_0_I28391 (.Y(N15867), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NOR2XL inst_cellmath__17_0_I4813 (.Y(inst_cellmath__17), .A(N15863), .B(N15867));
OR2XL cynw_cm_float_sin_I4814 (.Y(N487), .A(inst_cellmath__17), .B(inst_cellmath__68));
OR3XL cynw_cm_float_sin_I4815 (.Y(N759), .A(inst_cellmath__82), .B(inst_cellmath__68), .C(N487));
NAND2XL inst_cellmath__216__184__I4817 (.Y(N15898), .A(a_exp[5]), .B(a_exp[6]));
NOR2XL inst_cellmath__216__184__I4818 (.Y(N15891), .A(N15749), .B(N15898));
NOR2X1 inst_cellmath__216__184__I4819 (.Y(N639), .A(a_exp[7]), .B(N15891));
NAND2XL hyperpropagate_3_1_A_I10799 (.Y(N22752), .A(inst_cellmath__201[48]), .B(inst_cellmath__61[22]));
NOR2XL hyperpropagate_3_1_A_I10800 (.Y(inst_cellmath__219), .A(N22595), .B(N22752));
INVX1 inst_cellmath__211__182__I4821 (.Y(N15983), .A(inst_cellmath__210[22]));
INVX1 inst_cellmath__211__182__I4822 (.Y(N15920), .A(inst_cellmath__210[0]));
INVX1 inst_cellmath__211__182__I4823 (.Y(N15959), .A(inst_cellmath__210[2]));
OAI21X1 inst_cellmath__211__182__I4824 (.Y(N15978), .A0(N15920), .A1(inst_cellmath__210[1]), .B0(N15959));
OR2XL inst_cellmath__211__182__I4825 (.Y(N15982), .A(inst_cellmath__210[1]), .B(inst_cellmath__210[2]));
INVX1 inst_cellmath__211__182__I4826 (.Y(N15945), .A(inst_cellmath__210[3]));
NOR2X1 inst_cellmath__211__182__I4827 (.Y(N15967), .A(inst_cellmath__210[4]), .B(N15945));
INVX1 inst_cellmath__211__182__I4828 (.Y(N15987), .A(inst_cellmath__210[6]));
OAI21X1 inst_cellmath__211__182__I4829 (.Y(N15917), .A0(inst_cellmath__210[5]), .A1(N15967), .B0(N15987));
NOR2X1 inst_cellmath__211__182__I4830 (.Y(N15934), .A(inst_cellmath__210[3]), .B(inst_cellmath__210[4]));
NOR2X2 inst_cellmath__211__182__I4831 (.Y(N15954), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[5]));
NOR2BX1 inst_cellmath__211__182__I10588 (.Y(N15994), .AN(inst_cellmath__210[7]), .B(inst_cellmath__210[8]));
INVXL inst_cellmath__211__182__I4834 (.Y(N15923), .A(inst_cellmath__210[10]));
OAI21X1 inst_cellmath__211__182__I4835 (.Y(N15941), .A0(inst_cellmath__210[9]), .A1(N15994), .B0(N15923));
NOR2X2 inst_cellmath__211__182__I4836 (.Y(N15963), .A(inst_cellmath__210[7]), .B(inst_cellmath__210[8]));
NOR2BX1 inst_cellmath__211__182__I10589 (.Y(N15931), .AN(inst_cellmath__210[11]), .B(inst_cellmath__210[12]));
INVXL inst_cellmath__211__182__I4840 (.Y(N15950), .A(inst_cellmath__210[14]));
OAI21X2 inst_cellmath__211__182__I4841 (.Y(N15972), .A0(inst_cellmath__210[13]), .A1(N15931), .B0(N15950));
NOR2X2 inst_cellmath__211__182__I4842 (.Y(N15992), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[11]));
NOR2X2 inst_cellmath__211__182__I4843 (.Y(N15921), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[13]));
NOR2BX1 inst_cellmath__211__182__I4844 (.Y(N15960), .AN(inst_cellmath__210[15]), .B(inst_cellmath__210[16]));
INVXL inst_cellmath__211__182__I4845 (.Y(N15980), .A(inst_cellmath__210[18]));
OAI21X1 inst_cellmath__211__182__I4846 (.Y(N15911), .A0(inst_cellmath__210[17]), .A1(N15960), .B0(N15980));
NOR2X1 inst_cellmath__211__182__I4847 (.Y(N15944), .A(inst_cellmath__210[15]), .B(inst_cellmath__210[16]));
NOR2X2 inst_cellmath__211__182__I4848 (.Y(N15946), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[17]));
INVX1 inst_cellmath__211__182__I4849 (.Y(N15970), .A(inst_cellmath__210[19]));
NOR2X1 inst_cellmath__211__182__I4850 (.Y(N15989), .A(N15970), .B(inst_cellmath__210[20]));
OAI21X2 inst_cellmath__211__182__I4851 (.Y(N15937), .A0(inst_cellmath__210[21]), .A1(N15989), .B0(N15983));
INVXL inst_cellmath__211__182__I4854 (.Y(N15928), .A(N15954));
NAND2X2 inst_cellmath__211__182__I4856 (.Y(N15990), .A(N15954), .B(N15934));
NAND2BXL inst_cellmath__211__182__I4857 (.Y(N15938), .AN(N15963), .B(N15984));
INVXL inst_cellmath__211__182__I4858 (.Y(N15958), .A(N15921));
NAND2X4 inst_cellmath__211__182__I4861 (.Y(N15926), .A(N15921), .B(N15992));
NOR2X1 cynw_cm_float_sin_I27925 (.Y(N15976), .A(inst_cellmath__210[21]), .B(inst_cellmath__210[22]));
NOR2X1 cynw_cm_float_sin_I27924 (.Y(N15956), .A(inst_cellmath__210[19]), .B(inst_cellmath__210[20]));
NAND2X2 cynw_cm_float_sin_I28062 (.Y(N15996), .A(N15984), .B(N15963));
NOR2X4 cynw_cm_float_sin_I27929 (.Y(N15935), .A(N15926), .B(N15996));
NAND2X2 cynw_cm_float_sin_I28064 (.Y(N15953), .A(N15976), .B(N15956));
NAND2X2 cynw_cm_float_sin_I28063 (.Y(N43693), .A(N15944), .B(N15946));
NOR2X2 cynw_cm_float_sin_I28069 (.Y(N15969), .A(N43693), .B(N15953));
NAND2BXL inst_cellmath__211__182__I4871 (.Y(N544), .AN(N15935), .B(N15969));
OAI21X2 inst_cellmath__211__182__I4878 (.Y(N15962), .A0(N15990), .A1(N15978), .B0(N15917));
OAI21X1 inst_cellmath__211__182__I4879 (.Y(N15913), .A0(N15926), .A1(N15941), .B0(N15972));
OAI21X2 inst_cellmath__211__182__I4880 (.Y(N15949), .A0(N15953), .A1(N15911), .B0(N15937));
AOI21XL cynw_cm_float_sin_I27926 (.Y(N43367), .A0(N15934), .A1(N15982), .B0(N15928));
AOI21X1 cynw_cm_float_sin_I27927 (.Y(N43337), .A0(N15992), .A1(N15938), .B0(N15958));
NAND2BXL cynw_cm_float_sin_I27928 (.Y(N43345), .AN(N15944), .B(N15946));
INVXL cynw_cm_float_sin_I28065 (.Y(N43708), .A(N15990));
INVXL cynw_cm_float_sin_I28066 (.Y(N43717), .A(N15926));
OAI21XL cynw_cm_float_sin_I28067 (.Y(N43689), .A0(N43708), .A1(N15996), .B0(N43717));
NAND2BXL cynw_cm_float_sin_I28068 (.Y(N43696), .AN(N15953), .B(N43693));
CLKINVX4 cynw_cm_float_sin_I28070 (.Y(N15952), .A(N15969));
OAI21X1 cynw_cm_float_sin_I28071 (.Y(N543), .A0(N43689), .A1(N15952), .B0(N43696));
AOI21X1 cynw_cm_float_sin_I28072 (.Y(N43706), .A0(N43367), .A1(N15935), .B0(N43337));
OAI2BB1X1 cynw_cm_float_sin_I28073 (.Y(N43715), .A0N(N15956), .A1N(N43345), .B0(N15976));
OAI21X2 cynw_cm_float_sin_I28074 (.Y(N542), .A0(N15952), .A1(N43706), .B0(N43715));
AOI21X2 cynw_cm_float_sin_I28075 (.Y(N43365), .A0(N15935), .A1(N15962), .B0(N15913));
INVX2 cynw_cm_float_sin_I28076 (.Y(N43335), .A(N15949));
OAI21X4 cynw_cm_float_sin_I28077 (.Y(N541), .A0(N15952), .A1(N43365), .B0(N43335));
AND2XL cynw_cm_float_sin_I28078 (.Y(N16062), .A(N542), .B(N541));
NAND2XL cynw_cm_float_sin_I28079 (.Y(N43713), .A(N541), .B(N542));
CLKXOR2X1 cynw_cm_float_sin_I28080 (.Y(inst_cellmath__215[2]), .A(N543), .B(N43713));
NAND2XL cynw_cm_float_sin_I4886 (.Y(N16065), .A(N542), .B(N543));
INVX2 cynw_cm_float_sin_I27941 (.Y(inst_cellmath__215[0]), .A(N541));
NOR2XL cynw_cm_float_sin_I4887 (.Y(N16069), .A(inst_cellmath__215[0]), .B(N16065));
INVXL gen2_alt_A_I28638 (.Y(N44129), .A(N544));
OAI2BB1X1 gen2_alt_A_I28639 (.Y(N16072), .A0N(N543), .A1N(N16062), .B0(N44129));
NOR2X1 cynw_cm_float_sin_I27937 (.Y(N43361), .A(N15952), .B(N43365));
INVXL cynw_cm_float_sin_I27938 (.Y(N43353), .A(N43335));
NOR2X1 cynw_cm_float_sin_I27939 (.Y(N43346), .A(N43353), .B(N43361));
MXI2X2 cynw_cm_float_sin_I27942 (.Y(inst_cellmath__215[1]), .A(N43346), .B(N541), .S0(N542));
XOR2XL cynw_cm_float_sin_I4892 (.Y(inst_cellmath__215[3]), .A(N16069), .B(N544));
INVX1 cynw_cm_float_sin_I4893 (.Y(N16063), .A(N16072));
MXI2X1 cynw_cm_float_sin_I4894 (.Y(inst_cellmath__215[4]), .A(N16063), .B(N16072), .S0(N15952));
CLKINVX4 inst_cellmath__220__188__I4895 (.Y(N16142), .A(inst_cellmath__215[0]));
AND2XL inst_cellmath__220__188__I4896 (.Y(N16241), .A(N16142), .B(inst_cellmath__210[0]));
MX2XL inst_cellmath__220__188__I4897 (.Y(N16154), .A(inst_cellmath__210[0]), .B(inst_cellmath__210[1]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4898 (.Y(N16188), .A(inst_cellmath__210[1]), .B(inst_cellmath__210[2]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4899 (.Y(N16222), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[3]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4900 (.Y(N16100), .A(inst_cellmath__210[3]), .B(inst_cellmath__210[4]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4901 (.Y(N16132), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[5]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4902 (.Y(N16169), .A(inst_cellmath__210[5]), .B(inst_cellmath__210[6]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4903 (.Y(N16203), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[7]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4904 (.Y(N16236), .A(inst_cellmath__210[7]), .B(inst_cellmath__210[8]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4905 (.Y(N16115), .A(inst_cellmath__210[8]), .B(inst_cellmath__210[9]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4906 (.Y(N16147), .A(inst_cellmath__210[9]), .B(inst_cellmath__210[10]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4907 (.Y(N16183), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[11]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4908 (.Y(N16214), .A(inst_cellmath__210[11]), .B(inst_cellmath__210[12]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4909 (.Y(N16093), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[13]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4910 (.Y(N16126), .A(inst_cellmath__210[13]), .B(inst_cellmath__210[14]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4911 (.Y(N16163), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[15]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4912 (.Y(N16197), .A(inst_cellmath__210[15]), .B(inst_cellmath__210[16]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4913 (.Y(N16231), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[17]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4914 (.Y(N16109), .A(inst_cellmath__210[17]), .B(inst_cellmath__210[18]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4915 (.Y(N16140), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[19]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4916 (.Y(N16176), .A(inst_cellmath__210[19]), .B(inst_cellmath__210[20]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4917 (.Y(N16208), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[21]), .S0(N16142));
MX2XL inst_cellmath__220__188__I4918 (.Y(N16087), .A(inst_cellmath__210[21]), .B(inst_cellmath__210[22]), .S0(N16142));
CLKINVX8 inst_cellmath__220__188__I4919 (.Y(N16178), .A(inst_cellmath__215[1]));
NAND2XL inst_cellmath__220__188__I4920 (.Y(N16105), .A(N16241), .B(N16178));
NAND2XL inst_cellmath__220__188__I4921 (.Y(N16175), .A(N16154), .B(N16178));
MXI2XL inst_cellmath__220__188__I4922 (.Y(N16240), .A(N16241), .B(N16188), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4923 (.Y(N16119), .A(N16154), .B(N16222), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4924 (.Y(N16153), .A(N16188), .B(N16100), .S0(N16178));
MXI2X1 inst_cellmath__220__188__I4925 (.Y(N16187), .A(N16222), .B(N16132), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4926 (.Y(N16220), .A(N16100), .B(N16169), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4927 (.Y(N16098), .A(N16132), .B(N16203), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4928 (.Y(N16131), .A(N16169), .B(N16236), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4929 (.Y(N16168), .A(N16203), .B(N16115), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4930 (.Y(N16202), .A(N16236), .B(N16147), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4931 (.Y(N16235), .A(N16115), .B(N16183), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4932 (.Y(N16114), .A(N16147), .B(N16214), .S0(N16178));
MXI2X1 inst_cellmath__220__188__I4933 (.Y(N16146), .A(N16183), .B(N16093), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4934 (.Y(N16182), .A(N16214), .B(N16126), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4935 (.Y(N16213), .A(N16093), .B(N16163), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4936 (.Y(N16092), .A(N16126), .B(N16197), .S0(N16178));
MXI2X1 inst_cellmath__220__188__I4937 (.Y(N16125), .A(N16163), .B(N16231), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4938 (.Y(N16162), .A(N16197), .B(N16109), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4939 (.Y(N16196), .A(N16231), .B(N16140), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4940 (.Y(N16230), .A(N16109), .B(N16176), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4941 (.Y(N16108), .A(N16140), .B(N16208), .S0(N16178));
MXI2XL inst_cellmath__220__188__I4942 (.Y(N16139), .A(N16176), .B(N16087), .S0(N16178));
INVX2 inst_cellmath__220__188__I4944 (.Y(N16104), .A(inst_cellmath__215[2]));
INVX2 inst_cellmath__220__188__I9974 (.Y(N22596), .A(N16104));
INVX1 inst_cellmath__220__188__I9978 (.Y(N22600), .A(N22596));
INVX1 inst_cellmath__220__188__I9977 (.Y(N22599), .A(N22596));
INVX1 inst_cellmath__220__188__I9976 (.Y(N22598), .A(N22596));
INVX2 inst_cellmath__220__188__I9975 (.Y(N22597), .A(N22596));
NOR2BX1 inst_cellmath__220__188__I10594 (.Y(N16158), .AN(N22596), .B(N16105));
NOR2XL inst_cellmath__220__188__I4948 (.Y(N16225), .A(N16175), .B(N22600));
NOR2XL inst_cellmath__220__188__I4949 (.Y(N16136), .A(N16240), .B(N22600));
NOR2XL inst_cellmath__220__188__I4950 (.Y(N16206), .A(N16119), .B(N22597));
MXI2XL inst_cellmath__220__188__I4951 (.Y(N16118), .A(N16153), .B(N16105), .S0(N22597));
MXI2X1 inst_cellmath__220__188__I4952 (.Y(N16151), .A(N16187), .B(N16175), .S0(N22597));
MXI2XL inst_cellmath__220__188__I4953 (.Y(N16186), .A(N16220), .B(N16240), .S0(N22597));
MXI2XL inst_cellmath__220__188__I4954 (.Y(N16218), .A(N16098), .B(N16119), .S0(N22598));
MXI2XL inst_cellmath__220__188__I4955 (.Y(N16096), .A(N16131), .B(N16153), .S0(N22598));
MXI2XL inst_cellmath__220__188__I4956 (.Y(N16130), .A(N16168), .B(N16187), .S0(N22598));
MXI2XL inst_cellmath__220__188__I4957 (.Y(N16166), .A(N16202), .B(N16220), .S0(N22599));
MXI2XL inst_cellmath__220__188__I4958 (.Y(N16201), .A(N16235), .B(N16098), .S0(N22599));
MXI2XL inst_cellmath__220__188__I4959 (.Y(N16234), .A(N16114), .B(N16131), .S0(N22599));
MXI2XL inst_cellmath__220__188__I4960 (.Y(N16113), .A(N16146), .B(N16168), .S0(N22599));
MXI2XL inst_cellmath__220__188__I4961 (.Y(N16144), .A(N16182), .B(N16202), .S0(N22599));
MXI2XL inst_cellmath__220__188__I4962 (.Y(N16181), .A(N16213), .B(N16235), .S0(N22597));
MXI2XL inst_cellmath__220__188__I4963 (.Y(N16212), .A(N16092), .B(N16114), .S0(N22598));
MXI2X1 inst_cellmath__220__188__I4964 (.Y(N16091), .A(N16125), .B(N16146), .S0(N16104));
MXI2XL inst_cellmath__220__188__I4965 (.Y(N16124), .A(N16162), .B(N16182), .S0(N22598));
MXI2XL inst_cellmath__220__188__I4966 (.Y(N16161), .A(N16196), .B(N16213), .S0(N22600));
MXI2XL inst_cellmath__220__188__I4967 (.Y(N16195), .A(N16230), .B(N16092), .S0(N22600));
MXI2XL inst_cellmath__220__188__I4968 (.Y(N16229), .A(N16108), .B(N16125), .S0(N16104));
MXI2XL inst_cellmath__220__188__I4969 (.Y(N16107), .A(N16139), .B(N16162), .S0(N22600));
INVX3 inst_cellmath__220__188__I4971 (.Y(N16219), .A(inst_cellmath__215[4]));
NAND2XL inst_cellmath__220__188__I4973 (.Y(N16121), .A(N16158), .B(N16219));
NAND2X1 inst_cellmath__220__188__I4974 (.Y(N16192), .A(N16225), .B(N16219));
NAND2XL inst_cellmath__220__188__I4975 (.Y(N16103), .A(N16136), .B(N16219));
NAND2XL inst_cellmath__220__188__I4976 (.Y(N16172), .A(N16206), .B(N16219));
NAND2XL inst_cellmath__220__188__I4977 (.Y(N16239), .A(N16118), .B(N16219));
NAND2XL inst_cellmath__220__188__I4978 (.Y(N16150), .A(N16151), .B(N16219));
NAND2XL inst_cellmath__220__188__I4979 (.Y(N16216), .A(N16186), .B(N16219));
NAND2XL inst_cellmath__220__188__I4980 (.Y(N16129), .A(N16218), .B(N16219));
NAND2XL inst_cellmath__220__188__I4981 (.Y(N16200), .A(N16096), .B(N16219));
NAND2XL inst_cellmath__220__188__I4982 (.Y(N16111), .A(N16130), .B(N16219));
NAND2XL inst_cellmath__220__188__I4983 (.Y(N16180), .A(N16166), .B(N16219));
NAND2XL inst_cellmath__220__188__I4984 (.Y(N16090), .A(N16201), .B(N16219));
NAND2XL inst_cellmath__220__188__I4985 (.Y(N16159), .A(N16234), .B(N16219));
NAND2XL inst_cellmath__220__188__I4986 (.Y(N16228), .A(N16113), .B(N16219));
NAND2XL inst_cellmath__220__188__I4987 (.Y(N16138), .A(N16144), .B(N16219));
NAND2XL inst_cellmath__220__188__I4988 (.Y(N16207), .A(N16181), .B(N16219));
MXI2XL inst_cellmath__220__188__I4989 (.Y(N16120), .A(N16158), .B(N16212), .S0(N16219));
MXI2X1 inst_cellmath__220__188__I4990 (.Y(N16155), .A(N16225), .B(N16091), .S0(N16219));
MXI2XL inst_cellmath__220__188__I4991 (.Y(N16189), .A(N16136), .B(N16124), .S0(N16219));
MXI2XL inst_cellmath__220__188__I4992 (.Y(N16221), .A(N16206), .B(N16161), .S0(N16219));
MXI2XL inst_cellmath__220__188__I4993 (.Y(N16099), .A(N16118), .B(N16195), .S0(N16219));
MXI2XL inst_cellmath__220__188__I4994 (.Y(N16133), .A(N16151), .B(N16229), .S0(N16219));
MXI2XL inst_cellmath__220__188__I4995 (.Y(N16170), .A(N16186), .B(N16107), .S0(N16219));
CLKINVX4 inst_cellmath__220__188__I4997 (.Y(N16145), .A(inst_cellmath__215[3]));
NOR2XL inst_cellmath__220__188__I4999 (.Y(N679), .A(N16121), .B(N16145));
NOR2X1 inst_cellmath__220__188__I5000 (.Y(N680), .A(N16145), .B(N16192));
NOR2X1 inst_cellmath__220__188__I5001 (.Y(N681), .A(N16145), .B(N16103));
NOR2XL inst_cellmath__220__188__I5002 (.Y(N682), .A(N16172), .B(N16145));
NOR2XL inst_cellmath__220__188__I5003 (.Y(N683), .A(N16145), .B(N16239));
NOR2XL inst_cellmath__220__188__I5004 (.Y(N684), .A(N16150), .B(N16145));
NOR2XL inst_cellmath__220__188__I5005 (.Y(N685), .A(N16216), .B(N16145));
NOR2XL inst_cellmath__220__188__I5006 (.Y(N686), .A(N16129), .B(N16145));
MXI2XL inst_cellmath__220__188__I5007 (.Y(N687), .A(N16200), .B(N16121), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5008 (.Y(N688), .A(N16111), .B(N16192), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5009 (.Y(N689), .A(N16180), .B(N16103), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5010 (.Y(N690), .A(N16090), .B(N16172), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5011 (.Y(N691), .A(N16159), .B(N16239), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5012 (.Y(N692), .A(N16228), .B(N16150), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5013 (.Y(N693), .A(N16138), .B(N16216), .S0(N16145));
MXI2X1 inst_cellmath__220__188__I5014 (.Y(N694), .A(N16207), .B(N16129), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5015 (.Y(N695), .A(N16120), .B(N16200), .S0(N16145));
MXI2X1 inst_cellmath__220__188__I5016 (.Y(N696), .A(N16155), .B(N16111), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5017 (.Y(N697), .A(N16189), .B(N16180), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5018 (.Y(N698), .A(N16221), .B(N16090), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5019 (.Y(N699), .A(N16099), .B(N16159), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5020 (.Y(N700), .A(N16133), .B(N16228), .S0(N16145));
MXI2XL inst_cellmath__220__188__I5021 (.Y(N701), .A(N16170), .B(N16138), .S0(N16145));
INVX1 cynw_cm_float_sin_I5026 (.Y(N675), .A(inst_cellmath__215[4]));
NOR2X1 inst_cellmath__220_2WWMM_I5027 (.Y(N16452), .A(inst_cellmath__219), .B(N639));
AOI22XL inst_cellmath__220_2WWMM_I5028 (.Y(N16405), .A0(a_exp[0]), .A1(N639), .B0(N16452), .B1(N16142));
AOI22XL inst_cellmath__220_2WWMM_I5029 (.Y(N16449), .A0(a_exp[1]), .A1(N639), .B0(N16452), .B1(N16178));
AOI22XL inst_cellmath__220_2WWMM_I5030 (.Y(N16391), .A0(a_exp[2]), .A1(N639), .B0(N16452), .B1(inst_cellmath__215[2]));
AOI22XL inst_cellmath__220_2WWMM_I5031 (.Y(N16436), .A0(a_exp[3]), .A1(N639), .B0(N16452), .B1(inst_cellmath__215[3]));
AOI22X2 inst_cellmath__220_2WWMM_I5032 (.Y(N16482), .A0(a_exp[4]), .A1(N639), .B0(N16452), .B1(N675));
AOI21XL inst_cellmath__220_2WWMM_I5033 (.Y(N16422), .A0(a_exp[5]), .A1(N639), .B0(N16452));
AOI21XL inst_cellmath__220_2WWMM_I5034 (.Y(N16468), .A0(a_exp[6]), .A1(N639), .B0(N16452));
AND2XL inst_cellmath__220_2WWMM_I5035 (.Y(N647), .A(a_exp[7]), .B(N639));
AO22XL inst_cellmath__220_2WWMM_I5036 (.Y(N648), .A0(N639), .A1(a_man[0]), .B0(N16452), .B1(N679));
AO22XL inst_cellmath__220_2WWMM_I5037 (.Y(N649), .A0(N639), .A1(a_man[1]), .B0(N16452), .B1(N680));
AO22XL inst_cellmath__220_2WWMM_I5038 (.Y(N650), .A0(N639), .A1(a_man[2]), .B0(N16452), .B1(N681));
AO22XL inst_cellmath__220_2WWMM_I5039 (.Y(N651), .A0(N639), .A1(a_man[3]), .B0(N16452), .B1(N682));
AO22XL inst_cellmath__220_2WWMM_I5040 (.Y(N652), .A0(N639), .A1(a_man[4]), .B0(N16452), .B1(N683));
AO22XL inst_cellmath__220_2WWMM_I5041 (.Y(N653), .A0(N639), .A1(a_man[5]), .B0(N16452), .B1(N684));
AO22XL inst_cellmath__220_2WWMM_I5042 (.Y(N654), .A0(N639), .A1(a_man[6]), .B0(N16452), .B1(N685));
AO22XL inst_cellmath__220_2WWMM_I5043 (.Y(N655), .A0(N639), .A1(a_man[7]), .B0(N16452), .B1(N686));
AO22XL inst_cellmath__220_2WWMM_I5044 (.Y(N656), .A0(N639), .A1(a_man[8]), .B0(N16452), .B1(N687));
AO22XL inst_cellmath__220_2WWMM_I5045 (.Y(N657), .A0(N639), .A1(a_man[9]), .B0(N16452), .B1(N688));
AO22XL inst_cellmath__220_2WWMM_I5046 (.Y(N658), .A0(N639), .A1(a_man[10]), .B0(N16452), .B1(N689));
AO22XL inst_cellmath__220_2WWMM_I5047 (.Y(N659), .A0(N639), .A1(a_man[11]), .B0(N16452), .B1(N690));
AO22XL inst_cellmath__220_2WWMM_I5048 (.Y(N660), .A0(N639), .A1(a_man[12]), .B0(N16452), .B1(N691));
AO22XL inst_cellmath__220_2WWMM_I5049 (.Y(N661), .A0(N639), .A1(a_man[13]), .B0(N16452), .B1(N692));
AO22XL inst_cellmath__220_2WWMM_I5050 (.Y(N662), .A0(N639), .A1(a_man[14]), .B0(N16452), .B1(N693));
AO22XL inst_cellmath__220_2WWMM_I5051 (.Y(N663), .A0(N639), .A1(a_man[15]), .B0(N16452), .B1(N694));
AO22XL inst_cellmath__220_2WWMM_I5052 (.Y(N664), .A0(N639), .A1(a_man[16]), .B0(N16452), .B1(N695));
AO22XL inst_cellmath__220_2WWMM_I5053 (.Y(N665), .A0(N639), .A1(a_man[17]), .B0(N16452), .B1(N696));
AO22XL inst_cellmath__220_2WWMM_I5054 (.Y(N666), .A0(N639), .A1(a_man[18]), .B0(N16452), .B1(N697));
AO22XL inst_cellmath__220_2WWMM_I5055 (.Y(N667), .A0(N639), .A1(a_man[19]), .B0(N16452), .B1(N698));
AO22XL inst_cellmath__220_2WWMM_I5056 (.Y(N668), .A0(N639), .A1(a_man[20]), .B0(N16452), .B1(N699));
AO22XL inst_cellmath__220_2WWMM_I5057 (.Y(N3584), .A0(N639), .A1(a_man[21]), .B0(N16452), .B1(N700));
AO22XL inst_cellmath__220_2WWMM_I5058 (.Y(N670), .A0(N639), .A1(a_man[22]), .B0(N16452), .B1(N701));
NAND2BXL inst_cellmath__220_2WWMM_I5059 (.Y(N16426), .AN(N639), .B(inst_cellmath__219));
NAND2XL inst_cellmath__220_2WWMM_I5060 (.Y(N640), .A(N16405), .B(N16426));
NAND2XL inst_cellmath__220_2WWMM_I5061 (.Y(N641), .A(N16426), .B(N16449));
NAND2XL inst_cellmath__220_2WWMM_I5062 (.Y(N642), .A(N16426), .B(N16391));
NAND2X1 inst_cellmath__220_2WWMM_I5063 (.Y(N643), .A(N16426), .B(N16436));
NAND2X2 inst_cellmath__220_2WWMM_I5064 (.Y(N644), .A(N16426), .B(N16482));
NAND2XL inst_cellmath__220_2WWMM_I5065 (.Y(N645), .A(N16422), .B(N16426));
NAND2XL inst_cellmath__220_2WWMM_I5066 (.Y(N646), .A(N16468), .B(N16426));
OR4X1 inst_cellmath__223__208__I5067 (.Y(N16530), .A(N647), .B(N645), .C(N646), .D(N640));
NOR3X1 inst_cellmath__223__208__I5068 (.Y(N16565), .A(N641), .B(N642), .C(N16530));
NOR2X1 inst_cellmath__223__208__I5069 (.Y(N16534), .A(N643), .B(N644));
NAND2X1 inst_cellmath__223__208__I5070 (.Y(N16557), .A(N16565), .B(N16534));
NOR3X1 inst_cellmath__223__208__I5071 (.Y(N16576), .A(N16557), .B(N648), .C(N655));
NOR3X2 inst_cellmath__223__208__I5072 (.Y(N16556), .A(N649), .B(N650), .C(N652));
NOR2XL inst_cellmath__223__208__I5073 (.Y(N16568), .A(N663), .B(N656));
NOR2XL inst_cellmath__223__208__I5074 (.Y(N16578), .A(N657), .B(N662));
NOR3XL inst_cellmath__223__208__I5075 (.Y(N16570), .A(N653), .B(N651), .C(N658));
NOR2XL inst_cellmath__223__208__I5076 (.Y(N16560), .A(N664), .B(N668));
NOR2X1 inst_cellmath__223__208__I5077 (.Y(N16572), .A(N665), .B(N3584));
NOR3XL inst_cellmath__223__208__I5078 (.Y(N16542), .A(N660), .B(N659), .C(N667));
OR3XL inst_cellmath__223__208__I5079 (.Y(N16540), .A(N661), .B(N654), .C(N666));
NAND2XL inst_cellmath__223__208__I5080 (.Y(N16535), .A(N16576), .B(N16568));
NAND2XL inst_cellmath__223__208__I5081 (.Y(N16547), .A(N16578), .B(N16560));
NAND2X1 inst_cellmath__223__208__I5082 (.Y(N16558), .A(N16556), .B(N16572));
NAND2XL inst_cellmath__223__208__I5083 (.Y(N16575), .A(N16570), .B(N16542));
NOR2XL inst_cellmath__223__208__I5084 (.Y(N16545), .A(N16540), .B(N16547));
OR2XL inst_cellmath__223__208__I5085 (.Y(N16563), .A(N16535), .B(N16558));
NOR2XL inst_cellmath__223__208__I5086 (.Y(N16532), .A(N16575), .B(N16563));
MXI2XL cynw_cm_float_sin_I5089 (.Y(N577), .A(N15829), .B(a_sign), .S0(N757));
NOR3BX1 inst_cellmath__223__199__I10186 (.Y(N16612), .AN(N577), .B(N487), .C(inst_cellmath__82));
OAI2BB1XL inst_cellmath__223__199__I9909 (.Y(N16607), .A0N(N16545), .A1N(N16532), .B0(N16612));
MXI2XL cynw_cm_float_sin_I5097 (.Y(x[31]), .A(N16607), .B(N15829), .S0(N639));
NAND2BXL cynw_cm_float_sin_I10187 (.Y(N580), .AN(inst_cellmath__82), .B(N487));
INVXL inst_cellmath__228_0_I5100 (.Y(N16646), .A(N759));
AO22XL inst_cellmath__228_0_I5101 (.Y(x[23]), .A0(N759), .A1(N580), .B0(N16646), .B1(N640));
AO22XL inst_cellmath__228_0_I5102 (.Y(x[24]), .A0(N759), .A1(N580), .B0(N16646), .B1(N641));
AO22XL inst_cellmath__228_0_I5103 (.Y(x[25]), .A0(N759), .A1(N580), .B0(N16646), .B1(N642));
AO22XL inst_cellmath__228_0_I5104 (.Y(x[26]), .A0(N759), .A1(N580), .B0(N16646), .B1(N643));
AO22XL inst_cellmath__228_0_I5105 (.Y(x[27]), .A0(N759), .A1(N580), .B0(N16646), .B1(N644));
AO22XL inst_cellmath__228_0_I5106 (.Y(x[28]), .A0(N759), .A1(N580), .B0(N16646), .B1(N645));
AO22XL inst_cellmath__228_0_I5107 (.Y(x[29]), .A0(N759), .A1(N580), .B0(N16646), .B1(N646));
AO22XL inst_cellmath__228_0_I5108 (.Y(x[30]), .A0(N759), .A1(N580), .B0(N16646), .B1(N647));
AO22XL inst_cellmath__231_0_I5110 (.Y(x[0]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N648));
AO22XL inst_cellmath__231_0_I5111 (.Y(x[1]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N649));
AO22XL inst_cellmath__231_0_I5112 (.Y(x[2]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N650));
AO22XL inst_cellmath__231_0_I5113 (.Y(x[3]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N651));
AO22XL inst_cellmath__231_0_I5114 (.Y(x[4]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N652));
AO22XL inst_cellmath__231_0_I5115 (.Y(x[5]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N653));
AO22XL inst_cellmath__231_0_I5116 (.Y(x[6]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N654));
AO22XL inst_cellmath__231_0_I5117 (.Y(x[7]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N655));
AO22XL inst_cellmath__231_0_I5118 (.Y(x[8]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N656));
AO22XL inst_cellmath__231_0_I5119 (.Y(x[9]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N657));
AO22XL inst_cellmath__231_0_I5120 (.Y(x[10]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N658));
AO22XL inst_cellmath__231_0_I5121 (.Y(x[11]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N659));
AO22XL inst_cellmath__231_0_I5122 (.Y(x[12]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N660));
AO22XL inst_cellmath__231_0_I5123 (.Y(x[13]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N661));
AO22XL inst_cellmath__231_0_I5124 (.Y(x[14]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N662));
AO22XL inst_cellmath__231_0_I5125 (.Y(x[15]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N663));
AO22XL inst_cellmath__231_0_I5126 (.Y(x[16]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N664));
AO22XL inst_cellmath__231_0_I5127 (.Y(x[17]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N665));
AO22XL inst_cellmath__231_0_I5128 (.Y(x[18]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N666));
AO22XL inst_cellmath__231_0_I5129 (.Y(x[19]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N667));
AO22XL inst_cellmath__231_0_I5130 (.Y(x[20]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N668));
AO22XL inst_cellmath__231_0_I5131 (.Y(x[21]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N3584));
AO22XL inst_cellmath__231_0_I5132 (.Y(x[22]), .A0(N759), .A1(inst_cellmath__82), .B0(N16646), .B1(N670));
assign inst_cellmath__42[0] = 1'B0;
assign inst_cellmath__42[2] = 1'B0;
assign inst_cellmath__42[3] = 1'B0;
assign inst_cellmath__42[5] = 1'B0;
assign inst_cellmath__42[6] = 1'B0;
assign inst_cellmath__42[7] = 1'B0;
assign inst_cellmath__42[8] = 1'B0;
assign inst_cellmath__61[0] = 1'B0;
assign inst_cellmath__61[3] = 1'B0;
assign inst_cellmath__61[4] = 1'B0;
assign inst_cellmath__61[7] = 1'B0;
assign inst_cellmath__61[8] = 1'B0;
assign inst_cellmath__61[9] = 1'B0;
assign inst_cellmath__61[16] = 1'B0;
assign inst_cellmath__195[4] = 1'B0;
assign inst_cellmath__195[5] = 1'B0;
assign inst_cellmath__197[0] = 1'B0;
assign inst_cellmath__197[1] = 1'B0;
assign inst_cellmath__197[2] = 1'B0;
assign inst_cellmath__197[3] = 1'B0;
assign inst_cellmath__197[4] = 1'B0;
assign inst_cellmath__197[7] = 1'B0;
assign inst_cellmath__197[9] = 1'B0;
assign inst_cellmath__197[10] = 1'B0;
assign inst_cellmath__197[11] = 1'B0;
assign inst_cellmath__197[12] = 1'B0;
assign inst_cellmath__197[13] = 1'B0;
assign inst_cellmath__197[14] = 1'B0;
assign inst_cellmath__197[15] = 1'B0;
assign inst_cellmath__197[17] = 1'B0;
assign inst_cellmath__197[18] = 1'B0;
assign inst_cellmath__197[19] = 1'B0;
assign inst_cellmath__197[20] = 1'B1;
assign inst_cellmath__198[0] = 1'B0;
assign inst_cellmath__198[1] = 1'B0;
assign inst_cellmath__198[2] = 1'B0;
assign inst_cellmath__198[3] = 1'B0;
assign inst_cellmath__198[4] = 1'B0;
assign inst_cellmath__198[5] = 1'B0;
assign inst_cellmath__198[6] = 1'B0;
assign inst_cellmath__198[7] = 1'B0;
assign inst_cellmath__198[8] = 1'B0;
assign inst_cellmath__198[9] = 1'B0;
assign inst_cellmath__198[10] = 1'B0;
assign inst_cellmath__198[11] = 1'B0;
assign inst_cellmath__198[12] = 1'B0;
assign inst_cellmath__198[13] = 1'B0;
assign inst_cellmath__198[14] = 1'B0;
assign inst_cellmath__198[15] = 1'B0;
assign inst_cellmath__198[16] = 1'B0;
assign inst_cellmath__198[17] = 1'B0;
assign inst_cellmath__201[0] = 1'B0;
assign inst_cellmath__201[1] = 1'B0;
assign inst_cellmath__201[2] = 1'B0;
assign inst_cellmath__201[3] = 1'B0;
assign inst_cellmath__201[4] = 1'B0;
assign inst_cellmath__201[5] = 1'B0;
assign inst_cellmath__201[6] = 1'B0;
assign inst_cellmath__201[7] = 1'B0;
assign inst_cellmath__201[8] = 1'B0;
assign inst_cellmath__201[9] = 1'B0;
assign inst_cellmath__201[10] = 1'B0;
assign inst_cellmath__201[11] = 1'B0;
assign inst_cellmath__201[12] = 1'B0;
assign inst_cellmath__201[13] = 1'B0;
assign inst_cellmath__201[14] = 1'B0;
assign inst_cellmath__201[15] = 1'B0;
assign inst_cellmath__201[16] = 1'B0;
assign inst_cellmath__201[17] = 1'B0;
assign inst_cellmath__201[18] = 1'B0;
assign inst_cellmath__201[19] = 1'B0;
assign inst_cellmath__201[20] = 1'B0;
assign inst_cellmath__201[21] = 1'B0;
assign inst_cellmath__201[22] = 1'B0;
assign inst_cellmath__201[23] = 1'B0;
assign inst_cellmath__201[24] = 1'B0;
assign inst_cellmath__201[34] = 1'B0;
assign inst_cellmath__201[35] = 1'B0;
assign inst_cellmath__201[45] = 1'B0;
assign inst_cellmath__201[49] = 1'B0;
assign inst_cellmath__203__W0[0] = 1'B0;
assign inst_cellmath__203__W0[2] = 1'B0;
assign inst_cellmath__203__W0[22] = 1'B0;
assign inst_cellmath__203__W0[23] = 1'B0;
assign inst_cellmath__203__W0[43] = 1'B1;
assign inst_cellmath__203__W0[44] = 1'B1;
assign inst_cellmath__203__W0[45] = 1'B1;
assign inst_cellmath__203__W0[46] = 1'B1;
assign inst_cellmath__203__W1[0] = 1'B0;
assign inst_cellmath__203__W1[22] = 1'B0;
assign inst_cellmath__203__W1[23] = 1'B0;
assign inst_cellmath__203__W1[43] = 1'B0;
assign inst_cellmath__203__W1[44] = 1'B0;
assign inst_cellmath__203__W1[45] = 1'B0;
assign inst_cellmath__203__W1[46] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  v7b4TwHbrBE= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




