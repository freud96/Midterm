/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:12 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_div_ieee_E8_M23_0 (
	clk,
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	accept,
	x
	); /* architecture "gate_level" */ 
input  clk;
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input  accept;
output [31:0] x;
wire [31:0] inst_cellmath__8,
	inst_cellmath__9;
wire  inst_cellmath__11;
wire [3:0] inst_cellmath__12,
	inst_cellmath__13;
wire [25:0] inst_cellmath__14,
	inst_cellmath__16,
	inst_cellmath__17;
wire [4:0] inst_cellmath__22,
	inst_cellmath__23;
wire [6:0] inst_lookup0_cellmath__27;
wire [2:0] inst_lookup0_cellmath__29;
wire [25:0] inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__34,
	inst_cellmath__35,
	inst_cellmath__38__W0,
	inst_cellmath__38__W1,
	inst_cellmath__39__W0,
	inst_cellmath__39__W1;
wire [28:0] inst_cellmath__40,
	inst_cellmath__41,
	inst_cellmath__42,
	inst_cellmath__43,
	inst_cellmath__44,
	inst_cellmath__45,
	inst_cellmath__46,
	inst_cellmath__47;
wire [1:0] inst_cellmath__50;
wire [6:0] inst_it2_lookup1_cellmath__53;
wire [2:0] inst_it2_lookup1_cellmath__55;
wire [25:0] inst_it2_cellmath__56,
	inst_it2_cellmath__57,
	inst_it2_cellmath__60,
	inst_it2_cellmath__61,
	inst_it2_cellmath__62__W0,
	inst_it2_cellmath__62__W1,
	inst_it2_cellmath__63__W1;
wire [1:0] inst_it2_cellmath__66;
wire [9:0] inst_cellmath__67,
	inst_cellmath__68;
wire  inst_cellmath__69,
	inst_cellmath__70,
	inst_cellmath__71,
	inst_cellmath__72,
	inst_cellmath__73,
	inst_cellmath__74,
	inst_cellmath__75,
	inst_cellmath__76,
	inst_cellmath__77,
	inst_cellmath__78,
	inst_cellmath__79,
	inst_cellmath__80,
	inst_cellmath__83,
	inst_cellmath__84,
	inst_cellmath__85,
	inst_cellmath__86,
	inst_cellmath__87,
	inst_cellmath__88,
	inst_cellmath__89,
	inst_cellmath__91,
	inst_cellmath__96,
	inst_cellmath__100,
	inst_cellmath__101,
	inst_cellmath__102,
	inst_cellmath__103,
	inst_cellmath__104,
	inst_cellmath__105,
	inst_cellmath__106,
	inst_cellmath__109;
wire [7:0] inst_cellmath__110,
	inst_cellmath__111;
wire [21:0] inst_cellmath__112;
wire [31:0] inst_cellmath__113;
wire [25:0] inst_cellmath__120;
wire  inst_cellmath__122;
wire [28:0] inst_cellmath__124;
wire [22:0] inst_cellmath__125;
wire  inst_cellmath__126,
	inst_cellmath__127;
wire [22:0] inst_cellmath__129;
wire  inst_cellmath__135,
	inst_cellmath__136,
	inst_cellmath__137;
wire N1322,N1323,N1324,N1325,N1326,N1327,N1386 
	,N1387,N1388,N1417,N1447,N1527,N1528,N1555,N1587 
	,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680 
	,N1681,N1682,N1683,N1685,N1694,N1719,N1750,N1751 
	,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759 
	,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767 
	,N1768,N1769,N1770,N1771,N1772,N1847,N1848,N1873 
	,N1874,N1922,N2045,N2046,N2047,N2048,N2049,N2050 
	,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058 
	,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066 
	,N2067,N2068,N2150,N2151,N2152,N2153,N2154,N2155 
	,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163 
	,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171 
	,N2172,N2173,N2201,N2202,N2203,N2204,N2205,N2206 
	,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214 
	,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222 
	,N2223,N2224,N2254,N2255,N2256,N2257,N2258,N2259 
	,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267 
	,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275 
	,N2276,N2277,N4587,N4594;
EDFFHQX1 inst_cellmath__0_0_0__I0 (.Q(x[0]), .D(inst_cellmath__113[0]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_1__I1 (.Q(x[1]), .D(inst_cellmath__113[1]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_2__I2 (.Q(x[2]), .D(inst_cellmath__113[2]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_3__I3 (.Q(x[3]), .D(inst_cellmath__113[3]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_4__I4 (.Q(x[4]), .D(inst_cellmath__113[4]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_5__I5 (.Q(x[5]), .D(inst_cellmath__113[5]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_6__I6 (.Q(x[6]), .D(inst_cellmath__113[6]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_7__I7 (.Q(x[7]), .D(inst_cellmath__113[7]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_8__I8 (.Q(x[8]), .D(inst_cellmath__113[8]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_9__I9 (.Q(x[9]), .D(inst_cellmath__113[9]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_10__I10 (.Q(x[10]), .D(inst_cellmath__113[10]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_11__I11 (.Q(x[11]), .D(inst_cellmath__113[11]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_12__I12 (.Q(x[12]), .D(inst_cellmath__113[12]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_13__I13 (.Q(x[13]), .D(inst_cellmath__113[13]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_14__I14 (.Q(x[14]), .D(inst_cellmath__113[14]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_15__I15 (.Q(x[15]), .D(inst_cellmath__113[15]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_16__I16 (.Q(x[16]), .D(inst_cellmath__113[16]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_17__I17 (.Q(x[17]), .D(inst_cellmath__113[17]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_18__I18 (.Q(x[18]), .D(inst_cellmath__113[18]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_19__I19 (.Q(x[19]), .D(inst_cellmath__113[19]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_20__I20 (.Q(x[20]), .D(inst_cellmath__113[20]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_21__I21 (.Q(x[21]), .D(inst_cellmath__113[21]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_22__I22 (.Q(x[22]), .D(inst_cellmath__113[22]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_23__I23 (.Q(x[23]), .D(inst_cellmath__113[23]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_24__I24 (.Q(x[24]), .D(inst_cellmath__113[24]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_25__I25 (.Q(x[25]), .D(inst_cellmath__113[25]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_26__I26 (.Q(x[26]), .D(inst_cellmath__113[26]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_27__I27 (.Q(x[27]), .D(inst_cellmath__113[27]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_28__I28 (.Q(x[28]), .D(inst_cellmath__113[28]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_29__I29 (.Q(x[29]), .D(inst_cellmath__113[29]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_30__I30 (.Q(x[30]), .D(inst_cellmath__113[30]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__0_0_31__I31 (.Q(x[31]), .D(inst_cellmath__113[31]), .E(N4594), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_0__I32 (.Q(inst_cellmath__9[0]), .D(b_man[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_1__I33 (.Q(inst_cellmath__9[1]), .D(b_man[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_2__I34 (.Q(inst_cellmath__9[2]), .D(b_man[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_3__I35 (.Q(inst_cellmath__9[3]), .D(b_man[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_4__I36 (.Q(inst_cellmath__9[4]), .D(b_man[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_5__I37 (.Q(inst_cellmath__9[5]), .D(b_man[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_6__I38 (.Q(inst_cellmath__9[6]), .D(b_man[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_7__I39 (.Q(inst_cellmath__9[7]), .D(b_man[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_8__I40 (.Q(inst_cellmath__9[8]), .D(b_man[8]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_9__I41 (.Q(inst_cellmath__9[9]), .D(b_man[9]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_10__I42 (.Q(inst_cellmath__9[10]), .D(b_man[10]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_11__I43 (.Q(inst_cellmath__9[11]), .D(b_man[11]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_12__I44 (.Q(inst_cellmath__9[12]), .D(b_man[12]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_13__I45 (.Q(inst_cellmath__9[13]), .D(b_man[13]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_14__I46 (.Q(inst_cellmath__9[14]), .D(b_man[14]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_15__I47 (.Q(inst_cellmath__9[15]), .D(b_man[15]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_16__I48 (.Q(inst_cellmath__9[16]), .D(b_man[16]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_17__I49 (.Q(inst_cellmath__9[17]), .D(b_man[17]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_18__I50 (.Q(inst_cellmath__9[18]), .D(b_man[18]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_19__I51 (.Q(inst_cellmath__9[19]), .D(b_man[19]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_20__I52 (.Q(inst_cellmath__9[20]), .D(b_man[20]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_21__I53 (.Q(inst_it2_lookup1_cellmath__53[0]), .D(b_man[21]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_22__I54 (.Q(inst_it2_lookup1_cellmath__53[1]), .D(b_man[22]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_23__I55 (.Q(inst_cellmath__9[23]), .D(b_exp[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_24__I56 (.Q(inst_cellmath__9[24]), .D(b_exp[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_25__I57 (.Q(inst_cellmath__9[25]), .D(b_exp[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_26__I58 (.Q(inst_cellmath__9[26]), .D(b_exp[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_27__I59 (.Q(inst_cellmath__9[27]), .D(b_exp[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_28__I60 (.Q(inst_cellmath__9[28]), .D(b_exp[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_29__I61 (.Q(inst_cellmath__9[29]), .D(b_exp[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_30__I62 (.Q(inst_cellmath__9[30]), .D(b_exp[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__9_0_31__I63 (.Q(inst_cellmath__9[31]), .D(b_sign), .E(accept), .CK(clk));
DFFQXL inst_cellmath__11_0_I64 (.Q(inst_cellmath__11), .D(accept), .CK(clk));
DFFQXL inst_cellmath__16_0_1__I65 (.Q(inst_cellmath__16[1]), .D(inst_cellmath__14[1]), .CK(clk));
DFFQXL inst_cellmath__16_0_2__I66 (.Q(inst_cellmath__16[2]), .D(inst_cellmath__14[2]), .CK(clk));
DFFQXL inst_cellmath__16_0_3__I67 (.Q(inst_cellmath__16[3]), .D(inst_cellmath__14[3]), .CK(clk));
DFFQXL inst_cellmath__16_0_4__I68 (.Q(inst_cellmath__16[4]), .D(inst_cellmath__14[4]), .CK(clk));
DFFQXL inst_cellmath__16_0_5__I69 (.Q(inst_cellmath__16[5]), .D(inst_cellmath__14[5]), .CK(clk));
DFFQXL inst_cellmath__16_0_6__I70 (.Q(inst_cellmath__16[6]), .D(inst_cellmath__14[6]), .CK(clk));
DFFQXL inst_cellmath__16_0_7__I71 (.Q(inst_cellmath__16[7]), .D(inst_cellmath__14[7]), .CK(clk));
DFFQXL inst_cellmath__16_0_8__I72 (.Q(inst_cellmath__16[8]), .D(inst_cellmath__14[8]), .CK(clk));
DFFQXL inst_cellmath__16_0_9__I73 (.Q(inst_cellmath__16[9]), .D(inst_cellmath__14[9]), .CK(clk));
DFFQXL inst_cellmath__16_0_10__I74 (.Q(inst_cellmath__16[10]), .D(inst_cellmath__14[10]), .CK(clk));
DFFQXL inst_cellmath__16_0_11__I75 (.Q(inst_cellmath__16[11]), .D(inst_cellmath__14[11]), .CK(clk));
DFFQXL inst_cellmath__16_0_12__I76 (.Q(inst_cellmath__16[12]), .D(inst_cellmath__14[12]), .CK(clk));
DFFQXL inst_cellmath__16_0_13__I77 (.Q(inst_cellmath__16[13]), .D(inst_cellmath__14[13]), .CK(clk));
DFFQXL inst_cellmath__16_0_14__I78 (.Q(inst_cellmath__16[14]), .D(inst_cellmath__14[14]), .CK(clk));
DFFQXL inst_cellmath__16_0_15__I79 (.Q(inst_cellmath__16[15]), .D(inst_cellmath__14[15]), .CK(clk));
DFFQXL inst_cellmath__16_0_16__I80 (.Q(inst_cellmath__16[16]), .D(inst_cellmath__14[16]), .CK(clk));
DFFQXL inst_cellmath__16_0_17__I81 (.Q(inst_cellmath__16[17]), .D(inst_cellmath__14[17]), .CK(clk));
DFFQXL inst_cellmath__16_0_18__I82 (.Q(inst_cellmath__16[18]), .D(inst_cellmath__14[18]), .CK(clk));
DFFQXL inst_cellmath__16_0_19__I83 (.Q(inst_cellmath__16[19]), .D(inst_cellmath__14[19]), .CK(clk));
DFFQXL inst_cellmath__16_0_20__I84 (.Q(inst_cellmath__16[20]), .D(inst_cellmath__14[20]), .CK(clk));
DFFQXL inst_cellmath__16_0_21__I85 (.Q(inst_cellmath__16[21]), .D(inst_cellmath__14[21]), .CK(clk));
DFFQXL inst_cellmath__16_0_22__I86 (.Q(inst_cellmath__16[22]), .D(inst_cellmath__14[22]), .CK(clk));
DFFQXL inst_cellmath__16_0_23__I87 (.Q(inst_cellmath__16[23]), .D(inst_cellmath__14[23]), .CK(clk));
DFFQXL inst_cellmath__16_0_24__I88 (.Q(inst_cellmath__16[24]), .D(inst_cellmath__14[24]), .CK(clk));
DFFQXL inst_cellmath__16_0_25__I89 (.Q(inst_cellmath__16[25]), .D(inst_cellmath__14[25]), .CK(clk));
DFFQXL inst_cellmath__17_0_0__I90 (.Q(inst_cellmath__17[0]), .D(inst_it2_cellmath__63__W1[0]), .CK(clk));
DFFQXL inst_cellmath__17_0_1__I91 (.Q(inst_cellmath__17[1]), .D(inst_it2_cellmath__63__W1[1]), .CK(clk));
DFFQXL inst_cellmath__17_0_2__I92 (.Q(inst_cellmath__17[2]), .D(inst_it2_cellmath__63__W1[2]), .CK(clk));
DFFQXL inst_cellmath__17_0_3__I93 (.Q(inst_cellmath__17[3]), .D(inst_it2_cellmath__63__W1[3]), .CK(clk));
DFFQXL inst_cellmath__17_0_4__I94 (.Q(inst_cellmath__17[4]), .D(inst_it2_cellmath__63__W1[4]), .CK(clk));
DFFQXL inst_cellmath__17_0_5__I95 (.Q(inst_cellmath__17[5]), .D(inst_it2_cellmath__63__W1[5]), .CK(clk));
DFFQXL inst_cellmath__17_0_6__I96 (.Q(inst_cellmath__17[6]), .D(inst_it2_cellmath__63__W1[6]), .CK(clk));
DFFQXL inst_cellmath__17_0_7__I97 (.Q(inst_cellmath__17[7]), .D(inst_it2_cellmath__63__W1[7]), .CK(clk));
DFFQXL inst_cellmath__17_0_8__I98 (.Q(inst_cellmath__17[8]), .D(inst_it2_cellmath__63__W1[8]), .CK(clk));
DFFQXL inst_cellmath__17_0_9__I99 (.Q(inst_cellmath__17[9]), .D(inst_it2_cellmath__63__W1[9]), .CK(clk));
DFFQXL inst_cellmath__17_0_10__I100 (.Q(inst_cellmath__17[10]), .D(inst_it2_cellmath__63__W1[10]), .CK(clk));
DFFQXL inst_cellmath__17_0_11__I101 (.Q(inst_cellmath__17[11]), .D(inst_it2_cellmath__63__W1[11]), .CK(clk));
DFFQXL inst_cellmath__17_0_12__I102 (.Q(inst_cellmath__17[12]), .D(inst_it2_cellmath__63__W1[12]), .CK(clk));
DFFQXL inst_cellmath__17_0_13__I103 (.Q(inst_cellmath__17[13]), .D(inst_it2_cellmath__63__W1[13]), .CK(clk));
DFFQXL inst_cellmath__17_0_14__I104 (.Q(inst_cellmath__17[14]), .D(inst_it2_cellmath__63__W1[14]), .CK(clk));
DFFQXL inst_cellmath__17_0_15__I105 (.Q(inst_cellmath__17[15]), .D(inst_it2_cellmath__63__W1[15]), .CK(clk));
DFFQXL inst_cellmath__17_0_16__I106 (.Q(inst_cellmath__17[16]), .D(inst_it2_cellmath__63__W1[16]), .CK(clk));
DFFQXL inst_cellmath__17_0_17__I107 (.Q(inst_cellmath__17[17]), .D(inst_it2_cellmath__63__W1[17]), .CK(clk));
DFFQXL inst_cellmath__17_0_18__I108 (.Q(inst_cellmath__17[18]), .D(inst_it2_cellmath__63__W1[18]), .CK(clk));
DFFQXL inst_cellmath__17_0_19__I109 (.Q(inst_cellmath__17[19]), .D(inst_it2_cellmath__63__W1[19]), .CK(clk));
DFFQXL inst_cellmath__17_0_20__I110 (.Q(inst_cellmath__17[20]), .D(inst_it2_cellmath__63__W1[20]), .CK(clk));
DFFQXL inst_cellmath__17_0_21__I111 (.Q(inst_cellmath__17[21]), .D(inst_it2_cellmath__63__W1[21]), .CK(clk));
DFFQXL inst_cellmath__17_0_22__I112 (.Q(inst_cellmath__17[22]), .D(inst_it2_cellmath__63__W1[22]), .CK(clk));
DFFQXL inst_cellmath__17_0_23__I113 (.Q(inst_cellmath__17[23]), .D(inst_it2_cellmath__63__W1[23]), .CK(clk));
DFFQXL inst_cellmath__17_0_24__I114 (.Q(inst_cellmath__17[24]), .D(inst_it2_cellmath__63__W1[24]), .CK(clk));
DFFQXL inst_cellmath__17_0_25__I115 (.Q(inst_cellmath__17[25]), .D(inst_it2_cellmath__63__W1[25]), .CK(clk));
cynw_cm_float_div_ieee_inst_cellmath__23_0_bdw410776230_bdw cynw_cm_float_div_ieee_I116 (.inst_cellmath__23_0_out0({inst_cellmath__23[4], inst_cellmath__23[3], inst_cellmath__23[2], inst_cellmath__23[1], inst_cellmath__23[0]}), .inst_cellmath__23_0_in0({inst_cellmath__17[25], inst_cellmath__17[24], inst_cellmath__17[23], inst_cellmath__17[22], inst_cellmath__17[21]}), .inst_cellmath__23_0_in1({inst_cellmath__16[25], inst_cellmath__16[24], inst_cellmath__16[23], inst_cellmath__16[22], inst_cellmath__16[21]}));
EDFFHQX1 inst_cellmath__8_0_0__I117 (.Q(inst_cellmath__8[0]), .D(a_man[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_1__I118 (.Q(inst_cellmath__8[1]), .D(a_man[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_2__I119 (.Q(inst_cellmath__8[2]), .D(a_man[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_3__I120 (.Q(inst_cellmath__8[3]), .D(a_man[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_4__I121 (.Q(inst_cellmath__8[4]), .D(a_man[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_5__I122 (.Q(inst_cellmath__8[5]), .D(a_man[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_6__I123 (.Q(inst_cellmath__8[6]), .D(a_man[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_7__I124 (.Q(inst_cellmath__8[7]), .D(a_man[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_8__I125 (.Q(inst_cellmath__8[8]), .D(a_man[8]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_9__I126 (.Q(inst_cellmath__8[9]), .D(a_man[9]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_10__I127 (.Q(inst_cellmath__8[10]), .D(a_man[10]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_11__I128 (.Q(inst_cellmath__8[11]), .D(a_man[11]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_12__I129 (.Q(inst_cellmath__8[12]), .D(a_man[12]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_13__I130 (.Q(inst_cellmath__8[13]), .D(a_man[13]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_14__I131 (.Q(inst_cellmath__8[14]), .D(a_man[14]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_15__I132 (.Q(inst_cellmath__8[15]), .D(a_man[15]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_16__I133 (.Q(inst_cellmath__8[16]), .D(a_man[16]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_17__I134 (.Q(inst_cellmath__8[17]), .D(a_man[17]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_18__I135 (.Q(inst_cellmath__8[18]), .D(a_man[18]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_19__I136 (.Q(inst_cellmath__8[19]), .D(a_man[19]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_20__I137 (.Q(inst_cellmath__8[20]), .D(a_man[20]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_21__I138 (.Q(inst_cellmath__8[21]), .D(a_man[21]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_22__I139 (.Q(inst_cellmath__8[22]), .D(a_man[22]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_23__I140 (.Q(inst_cellmath__8[23]), .D(a_exp[0]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_24__I141 (.Q(inst_cellmath__8[24]), .D(a_exp[1]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_25__I142 (.Q(inst_cellmath__8[25]), .D(a_exp[2]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_26__I143 (.Q(inst_cellmath__8[26]), .D(a_exp[3]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_27__I144 (.Q(inst_cellmath__8[27]), .D(a_exp[4]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_28__I145 (.Q(inst_cellmath__8[28]), .D(a_exp[5]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_29__I146 (.Q(inst_cellmath__8[29]), .D(a_exp[6]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_30__I147 (.Q(inst_cellmath__8[30]), .D(a_exp[7]), .E(accept), .CK(clk));
EDFFHQX1 inst_cellmath__8_0_31__I148 (.Q(inst_cellmath__8[31]), .D(a_sign), .E(accept), .CK(clk));
INVXL cynw_cm_float_div_ieee_I149 (.Y(N1386), .A(inst_cellmath__9[20]));
INVXL cynw_cm_float_div_ieee_I150 (.Y(N1387), .A(inst_it2_lookup1_cellmath__53[0]));
INVXL cynw_cm_float_div_ieee_I151 (.Y(N1388), .A(inst_it2_lookup1_cellmath__53[1]));
cynw_cm_float_div_ieee_inst_cellmath__22_0_bdw410776230_bdw cynw_cm_float_div_ieee_I152 (.inst_cellmath__22_0_out0({inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}), .inst_cellmath__22_0_in0({inst_cellmath__8[22], inst_cellmath__8[21], inst_cellmath__8[20]}), .inst_cellmath__22_0_in1({N1388, N1387, N1386}));
cynw_cm_float_div_ieee_inst_cellmath__24_0_bdw410776230_bdw cynw_cm_float_div_ieee_I153 (.inst_cellmath__24_0_out0({inst_lookup0_cellmath__27[6], inst_lookup0_cellmath__27[5], inst_lookup0_cellmath__27[4], inst_lookup0_cellmath__27[3], inst_lookup0_cellmath__27[2]}), .inst_cellmath__24_0_in0({inst_cellmath__23[4], inst_cellmath__23[3], inst_cellmath__23[2], inst_cellmath__23[1], inst_cellmath__23[0]}), .inst_cellmath__24_0_in1({inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}), .inst_cellmath__24_0_in2(inst_cellmath__11));
cynw_cm_float_div_ieee_inst_lookup0_cellmath__29_0_bdw410776230_bdw cynw_cm_float_div_ieee_I154 (.inst_lookup0_cellmath__29_0_out0({inst_lookup0_cellmath__29[2], inst_lookup0_cellmath__29[1], inst_lookup0_cellmath__29[0]}), .inst_lookup0_cellmath__29_0_in0({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0]}), .inst_lookup0_cellmath__29_0_in1({inst_lookup0_cellmath__27[6], inst_lookup0_cellmath__27[5], inst_lookup0_cellmath__27[4], inst_lookup0_cellmath__27[3], inst_lookup0_cellmath__27[2]}));
cynw_cm_float_div_ieee_inst_cellmath__30__31__bdw410776230_bdw cynw_cm_float_div_ieee_I155 (.inst_cellmath__30__31__out0({N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N1694}), .inst_cellmath__30__31__in0({inst_lookup0_cellmath__29[0]}), .inst_cellmath__30__31__in1({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}));
cynw_cm_float_div_ieee_inst_cellmath__31__35__bdw410776230_bdw cynw_cm_float_div_ieee_I156 (.inst_cellmath__31__35__out0({N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N1848, N1847}), .inst_cellmath__31__35__in0({inst_lookup0_cellmath__29[1]}), .inst_cellmath__31__35__in1({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}));
cynw_cm_float_div_ieee_inst_cellmath__20_0_bdw410776230_bdw cynw_cm_float_div_ieee_I157 (.inst_cellmath__20_0_out0({inst_cellmath__34[25], inst_cellmath__34[24], inst_cellmath__34[23], inst_cellmath__34[22], inst_cellmath__34[21], inst_cellmath__34[20], inst_cellmath__34[19], inst_cellmath__34[18], inst_cellmath__34[17], inst_cellmath__34[16], inst_cellmath__34[15], inst_cellmath__34[14], inst_cellmath__34[13], inst_cellmath__34[12], inst_cellmath__34[11], inst_cellmath__34[10], inst_cellmath__34[9], inst_cellmath__34[8], inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2]}), .inst_cellmath__20_0_in0({inst_cellmath__8[22], inst_cellmath__8[21], inst_cellmath__8[20], inst_cellmath__8[19], inst_cellmath__8[18], inst_cellmath__8[17], inst_cellmath__8[16], inst_cellmath__8[15], inst_cellmath__8[14], inst_cellmath__8[13], inst_cellmath__8[12], inst_cellmath__8[11], inst_cellmath__8[10], inst_cellmath__8[9], inst_cellmath__8[8], inst_cellmath__8[7], inst_cellmath__8[6], inst_cellmath__8[5], inst_cellmath__8[4], inst_cellmath__8[3], inst_cellmath__8[2], inst_cellmath__8[1], inst_cellmath__8[0]}), .inst_cellmath__20_0_in1({inst_cellmath__16[23], inst_cellmath__16[22], inst_cellmath__16[21], inst_cellmath__16[20], inst_cellmath__16[19], inst_cellmath__16[18], inst_cellmath__16[17], inst_cellmath__16[16], inst_cellmath__16[15], inst_cellmath__16[14], inst_cellmath__16[13], inst_cellmath__16[12], inst_cellmath__16[11], inst_cellmath__16[10], inst_cellmath__16[9], inst_cellmath__16[8], inst_cellmath__16[7], inst_cellmath__16[6], inst_cellmath__16[5], inst_cellmath__16[4], inst_cellmath__16[3], inst_cellmath__16[2], inst_cellmath__16[1], 1'B0}), .inst_cellmath__20_0_in2(inst_cellmath__11));
INVXL cynw_cm_float_div_ieee_I158 (.Y(inst_cellmath__35[0]), .A(inst_lookup0_cellmath__29[2]));
cynw_cm_float_div_ieee_inst_cellmath__21_0_bdw410776230_bdw cynw_cm_float_div_ieee_I159 (.inst_cellmath__21_0_out0({inst_cellmath__35[25], inst_cellmath__35[24], inst_cellmath__35[23], inst_cellmath__35[22], inst_cellmath__35[21], inst_cellmath__35[20], inst_cellmath__35[19], inst_cellmath__35[18], inst_cellmath__35[17], inst_cellmath__35[16], inst_cellmath__35[15], inst_cellmath__35[14], inst_cellmath__35[13], inst_cellmath__35[12], inst_cellmath__35[11], inst_cellmath__35[10], inst_cellmath__35[9], inst_cellmath__35[8], inst_cellmath__35[7], inst_cellmath__35[6], inst_cellmath__35[5], inst_cellmath__35[4], inst_cellmath__35[3], inst_cellmath__35[2]}), .inst_cellmath__21_0_in0({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}), .inst_cellmath__21_0_in1({inst_cellmath__17[23], inst_cellmath__17[22], inst_cellmath__17[21], inst_cellmath__17[20], inst_cellmath__17[19], inst_cellmath__17[18], inst_cellmath__17[17], inst_cellmath__17[16], inst_cellmath__17[15], inst_cellmath__17[14], inst_cellmath__17[13], inst_cellmath__17[12], inst_cellmath__17[11], inst_cellmath__17[10], inst_cellmath__17[9], inst_cellmath__17[8], inst_cellmath__17[7], inst_cellmath__17[6], inst_cellmath__17[5], inst_cellmath__17[4], inst_cellmath__17[3], inst_cellmath__17[2], inst_cellmath__17[1], inst_cellmath__17[0]}), .inst_cellmath__21_0_in2(inst_cellmath__11));
cynw_cm_float_div_ieee_inst_cellmath__30_2mx_bdw410776230_bdw cynw_cm_float_div_ieee_I160 (.inst_cellmath__30_2mx_out0({inst_cellmath__30[25], inst_cellmath__30[24], inst_cellmath__30[23], inst_cellmath__30[22], inst_cellmath__30[21], inst_cellmath__30[20], inst_cellmath__30[19], inst_cellmath__30[18], inst_cellmath__30[17], inst_cellmath__30[16], inst_cellmath__30[15], inst_cellmath__30[14], inst_cellmath__30[13], inst_cellmath__30[12], inst_cellmath__30[11], inst_cellmath__30[10], inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}), .inst_cellmath__30_2mx_in0({inst_lookup0_cellmath__29[2]}), .inst_cellmath__30_2mx_in1({N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045}));
cynw_cm_float_div_ieee_inst_fa_1033_10_bdw410776230_bdw cynw_cm_float_div_ieee_I161 (.inst_fa_1033_10_out0({inst_cellmath__38__W1[25], inst_cellmath__38__W1[24], inst_cellmath__38__W1[23], inst_cellmath__38__W1[22], inst_cellmath__38__W1[21], inst_cellmath__38__W1[20], inst_cellmath__38__W1[19], inst_cellmath__38__W1[18], inst_cellmath__38__W1[17], inst_cellmath__38__W1[16], inst_cellmath__38__W1[15], inst_cellmath__38__W1[14], inst_cellmath__38__W1[13], inst_cellmath__38__W1[12], inst_cellmath__38__W1[11], inst_cellmath__38__W1[10], inst_cellmath__38__W1[9], inst_cellmath__38__W1[8], inst_cellmath__38__W1[7], inst_cellmath__38__W1[6], inst_cellmath__38__W1[5], inst_cellmath__38__W1[4], inst_cellmath__38__W1[3], inst_cellmath__38__W1[2], inst_cellmath__38__W1[1], inst_cellmath__38__W1[0]}), .inst_fa_1033_10_out1({inst_cellmath__38__W0[24], inst_cellmath__38__W0[23], inst_cellmath__38__W0[22], inst_cellmath__38__W0[21], inst_cellmath__38__W0[20], inst_cellmath__38__W0[19], inst_cellmath__38__W0[18], inst_cellmath__38__W0[17], inst_cellmath__38__W0[16], inst_cellmath__38__W0[15], inst_cellmath__38__W0[14], inst_cellmath__38__W0[13], inst_cellmath__38__W0[12], inst_cellmath__38__W0[11], inst_cellmath__38__W0[10], inst_cellmath__38__W0[9], inst_cellmath__38__W0[8], inst_cellmath__38__W0[7], inst_cellmath__38__W0[6], inst_cellmath__38__W0[5], inst_cellmath__38__W0[4], inst_cellmath__38__W0[3], inst_cellmath__38__W0[2], inst_cellmath__38__W0[1], inst_cellmath__38__W0[0]}), .inst_fa_1033_10_in0(inst_cellmath__35[0]), .inst_fa_1033_10_in1({inst_cellmath__30[25], inst_cellmath__30[24], inst_cellmath__30[23], inst_cellmath__30[22], inst_cellmath__30[21], inst_cellmath__30[20], inst_cellmath__30[19], inst_cellmath__30[18], inst_cellmath__30[17], inst_cellmath__30[16], inst_cellmath__30[15], inst_cellmath__30[14], inst_cellmath__30[13], inst_cellmath__30[12], inst_cellmath__30[11], inst_cellmath__30[10], inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}), .inst_fa_1033_10_in2({inst_cellmath__35[25], inst_cellmath__35[24], inst_cellmath__35[23], inst_cellmath__35[22], inst_cellmath__35[21], inst_cellmath__35[20], inst_cellmath__35[19], inst_cellmath__35[18], inst_cellmath__35[17], inst_cellmath__35[16], inst_cellmath__35[15], inst_cellmath__35[14], inst_cellmath__35[13], inst_cellmath__35[12], inst_cellmath__35[11], inst_cellmath__35[10], inst_cellmath__35[9], inst_cellmath__35[8], inst_cellmath__35[7], inst_cellmath__35[6], inst_cellmath__35[5], inst_cellmath__35[4], inst_cellmath__35[3], inst_cellmath__35[2]}), .inst_fa_1033_10_in3({inst_cellmath__34[25], inst_cellmath__34[24], inst_cellmath__34[23], inst_cellmath__34[22], inst_cellmath__34[21], inst_cellmath__34[20], inst_cellmath__34[19], inst_cellmath__34[18], inst_cellmath__34[17], inst_cellmath__34[16], inst_cellmath__34[15], inst_cellmath__34[14], inst_cellmath__34[13], inst_cellmath__34[12], inst_cellmath__34[11], inst_cellmath__34[10], inst_cellmath__34[9], inst_cellmath__34[8], inst_cellmath__34[7], inst_cellmath__34[6], inst_cellmath__34[5], inst_cellmath__34[4], inst_cellmath__34[3], inst_cellmath__34[2]}));
cynw_cm_float_div_ieee_inst_cellmath__31_2mx_bdw410776230_bdw cynw_cm_float_div_ieee_I162 (.inst_cellmath__31_2mx_out0({inst_cellmath__31[25], inst_cellmath__31[24], inst_cellmath__31[23], inst_cellmath__31[22], inst_cellmath__31[21], inst_cellmath__31[20], inst_cellmath__31[19], inst_cellmath__31[18], inst_cellmath__31[17], inst_cellmath__31[16], inst_cellmath__31[15], inst_cellmath__31[14], inst_cellmath__31[13], inst_cellmath__31[12], inst_cellmath__31[11], inst_cellmath__31[10], inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__31_2mx_in0({inst_lookup0_cellmath__29[2]}), .inst_cellmath__31_2mx_in1({N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150}));
cynw_cm_float_div_ieee_inst_fa_1052_10_bdw410776230_bdw cynw_cm_float_div_ieee_I163 (.inst_fa_1052_10_out0({inst_cellmath__39__W1[25], inst_cellmath__39__W1[24], inst_it2_cellmath__61[25], inst_it2_cellmath__61[24], inst_it2_cellmath__61[23], inst_it2_cellmath__61[22], inst_it2_cellmath__61[21], inst_it2_cellmath__61[20], inst_it2_cellmath__61[19], inst_it2_cellmath__61[18], inst_it2_cellmath__61[17], inst_it2_cellmath__61[16], inst_it2_cellmath__61[15], inst_it2_cellmath__61[14], inst_it2_cellmath__61[13], inst_it2_cellmath__61[12], inst_it2_cellmath__61[11], inst_it2_cellmath__61[10], inst_it2_cellmath__61[9], inst_it2_cellmath__61[8], inst_it2_cellmath__61[7], inst_it2_cellmath__61[6], inst_it2_cellmath__61[5], inst_it2_cellmath__61[4], inst_it2_cellmath__61[3], inst_it2_cellmath__61[2]}), .inst_fa_1052_10_out1({inst_cellmath__39__W0[24], inst_cellmath__39__W0[23], inst_it2_cellmath__60[25], inst_it2_cellmath__60[24], inst_it2_cellmath__60[23], inst_it2_cellmath__60[22], inst_it2_cellmath__60[21], inst_it2_cellmath__60[20], inst_it2_cellmath__60[19], inst_it2_cellmath__60[18], inst_it2_cellmath__60[17], inst_it2_cellmath__60[16], inst_it2_cellmath__60[15], inst_it2_cellmath__60[14], inst_it2_cellmath__60[13], inst_it2_cellmath__60[12], inst_it2_cellmath__60[11], inst_it2_cellmath__60[10], inst_it2_cellmath__60[9], inst_it2_cellmath__60[8], inst_it2_cellmath__60[7], inst_it2_cellmath__60[6], inst_it2_cellmath__60[5], inst_it2_cellmath__60[4], inst_it2_cellmath__60[3]}), .inst_fa_1052_10_in0({inst_cellmath__38__W1[25], inst_cellmath__38__W1[24], inst_cellmath__38__W1[23], inst_cellmath__38__W1[22], inst_cellmath__38__W1[21], inst_cellmath__38__W1[20], inst_cellmath__38__W1[19], inst_cellmath__38__W1[18], inst_cellmath__38__W1[17], inst_cellmath__38__W1[16], inst_cellmath__38__W1[15], inst_cellmath__38__W1[14], inst_cellmath__38__W1[13], inst_cellmath__38__W1[12], inst_cellmath__38__W1[11], inst_cellmath__38__W1[10], inst_cellmath__38__W1[9], inst_cellmath__38__W1[8], inst_cellmath__38__W1[7], inst_cellmath__38__W1[6], inst_cellmath__38__W1[5], inst_cellmath__38__W1[4], inst_cellmath__38__W1[3], inst_cellmath__38__W1[2], inst_cellmath__38__W1[1], inst_cellmath__38__W1[0]}), .inst_fa_1052_10_in1({inst_cellmath__38__W0[24], inst_cellmath__38__W0[23], inst_cellmath__38__W0[22], inst_cellmath__38__W0[21], inst_cellmath__38__W0[20], inst_cellmath__38__W0[19], inst_cellmath__38__W0[18], inst_cellmath__38__W0[17], inst_cellmath__38__W0[16], inst_cellmath__38__W0[15], inst_cellmath__38__W0[14], inst_cellmath__38__W0[13], inst_cellmath__38__W0[12], inst_cellmath__38__W0[11], inst_cellmath__38__W0[10], inst_cellmath__38__W0[9], inst_cellmath__38__W0[8], inst_cellmath__38__W0[7], inst_cellmath__38__W0[6], inst_cellmath__38__W0[5], inst_cellmath__38__W0[4], inst_cellmath__38__W0[3], inst_cellmath__38__W0[2], inst_cellmath__38__W0[1], inst_cellmath__38__W0[0]}), .inst_fa_1052_10_in2({inst_cellmath__31[25], inst_cellmath__31[24], inst_cellmath__31[23], inst_cellmath__31[22], inst_cellmath__31[21], inst_cellmath__31[20], inst_cellmath__31[19], inst_cellmath__31[18], inst_cellmath__31[17], inst_cellmath__31[16], inst_cellmath__31[15], inst_cellmath__31[14], inst_cellmath__31[13], inst_cellmath__31[12], inst_cellmath__31[11], inst_cellmath__31[10], inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}));
cynw_cm_float_div_ieee_inst_it2_cellmath__51_0_bdw410776230_bdw cynw_cm_float_div_ieee_I164 (.inst_it2_cellmath__51_0_out0({inst_it2_lookup1_cellmath__53[6], inst_it2_lookup1_cellmath__53[5], inst_it2_lookup1_cellmath__53[4], inst_it2_lookup1_cellmath__53[3], inst_it2_lookup1_cellmath__53[2]}), .inst_it2_cellmath__51_0_in0({inst_cellmath__39__W1[25], inst_cellmath__39__W1[24], inst_it2_cellmath__61[25], inst_it2_cellmath__61[24], inst_it2_cellmath__61[23]}), .inst_it2_cellmath__51_0_in1({inst_cellmath__39__W0[24], inst_cellmath__39__W0[23], inst_it2_cellmath__60[25], inst_it2_cellmath__60[24], inst_it2_cellmath__60[23]}));
cynw_cm_float_div_ieee_inst_it2_lookup1_cellmath__55_0_bdw410776230_bdw cynw_cm_float_div_ieee_I165 (.inst_it2_lookup1_cellmath__55_0_out0({inst_it2_lookup1_cellmath__55[2], inst_it2_lookup1_cellmath__55[1], inst_it2_lookup1_cellmath__55[0]}), .inst_it2_lookup1_cellmath__55_0_in0({inst_it2_lookup1_cellmath__53[6], inst_it2_lookup1_cellmath__53[5], inst_it2_lookup1_cellmath__53[4], inst_it2_lookup1_cellmath__53[3], inst_it2_lookup1_cellmath__53[2]}), .inst_it2_lookup1_cellmath__55_0_in1({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0]}));
cynw_cm_float_div_ieee_inst_it2_cellmath__56__57__bdw410776230_bdw cynw_cm_float_div_ieee_I166 (.inst_it2_cellmath__56__57__out0({N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N1719}), .inst_it2_cellmath__56__57__in0({inst_it2_lookup1_cellmath__55[0]}), .inst_it2_cellmath__56__57__in1({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}));
cynw_cm_float_div_ieee_inst_it2_cellmath__57__61__bdw410776230_bdw cynw_cm_float_div_ieee_I167 (.inst_it2_cellmath__57__61__out0({N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N1874, N1873}), .inst_it2_cellmath__57__61__in0({inst_it2_lookup1_cellmath__55[1]}), .inst_it2_cellmath__57__61__in1({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}));
DFFQXL inst_cellmath__112_0_0__I168 (.Q(inst_cellmath__112[0]), .D(N1751), .CK(clk));
DFFQXL inst_cellmath__112_0_1__I169 (.Q(inst_cellmath__112[1]), .D(N1752), .CK(clk));
DFFQXL inst_cellmath__112_0_2__I170 (.Q(inst_cellmath__112[2]), .D(N1753), .CK(clk));
DFFQXL inst_cellmath__112_0_3__I171 (.Q(inst_cellmath__112[3]), .D(N1754), .CK(clk));
DFFQXL inst_cellmath__112_0_4__I172 (.Q(inst_cellmath__112[4]), .D(N1755), .CK(clk));
DFFQXL inst_cellmath__112_0_5__I173 (.Q(inst_cellmath__112[5]), .D(N1756), .CK(clk));
DFFQXL inst_cellmath__112_0_6__I174 (.Q(inst_cellmath__112[6]), .D(N1757), .CK(clk));
DFFQXL inst_cellmath__112_0_7__I175 (.Q(inst_cellmath__112[7]), .D(N1758), .CK(clk));
DFFQXL inst_cellmath__112_0_8__I176 (.Q(inst_cellmath__112[8]), .D(N1759), .CK(clk));
DFFQXL inst_cellmath__112_0_9__I177 (.Q(inst_cellmath__112[9]), .D(N1760), .CK(clk));
DFFQXL inst_cellmath__112_0_10__I178 (.Q(inst_cellmath__112[10]), .D(N1761), .CK(clk));
DFFQXL inst_cellmath__112_0_11__I179 (.Q(inst_cellmath__112[11]), .D(N1762), .CK(clk));
DFFQXL inst_cellmath__112_0_12__I180 (.Q(inst_cellmath__112[12]), .D(N1763), .CK(clk));
DFFQXL inst_cellmath__112_0_13__I181 (.Q(inst_cellmath__112[13]), .D(N1764), .CK(clk));
DFFQXL inst_cellmath__112_0_14__I182 (.Q(inst_cellmath__112[14]), .D(N1765), .CK(clk));
DFFQXL inst_cellmath__112_0_15__I183 (.Q(inst_cellmath__112[15]), .D(N1766), .CK(clk));
DFFQXL inst_cellmath__112_0_16__I184 (.Q(inst_cellmath__112[16]), .D(N1767), .CK(clk));
DFFQXL inst_cellmath__112_0_17__I185 (.Q(inst_cellmath__112[17]), .D(N1768), .CK(clk));
DFFQXL inst_cellmath__112_0_18__I186 (.Q(inst_cellmath__112[18]), .D(N1769), .CK(clk));
DFFQXL inst_cellmath__112_0_19__I187 (.Q(inst_cellmath__112[19]), .D(N1770), .CK(clk));
DFFQXL inst_cellmath__112_0_20__I188 (.Q(inst_cellmath__112[20]), .D(N1771), .CK(clk));
DFFQXL inst_cellmath__112_0_21__I189 (.Q(inst_cellmath__112[21]), .D(N1772), .CK(clk));
cynw_cm_float_div_ieee_inst_cellmath__120_0_bdw410776230_bdw cynw_cm_float_div_ieee_I190 (.inst_cellmath__120_0_out0({inst_cellmath__120[25], inst_cellmath__120[24], inst_cellmath__120[23], inst_cellmath__120[22], inst_cellmath__120[21], inst_cellmath__120[20], inst_cellmath__120[19], inst_cellmath__120[18], inst_cellmath__120[17], inst_cellmath__120[16], inst_cellmath__120[15], inst_cellmath__120[14], inst_cellmath__120[13], inst_cellmath__120[12], inst_cellmath__120[11], inst_cellmath__120[10], inst_cellmath__120[9], inst_cellmath__120[8], inst_cellmath__120[7], inst_cellmath__120[6], inst_cellmath__120[5], inst_cellmath__120[4], inst_cellmath__120[3], inst_cellmath__120[2], inst_cellmath__120[1], inst_cellmath__120[0]}), .inst_cellmath__120_0_in0({inst_cellmath__17[25], inst_cellmath__17[24], inst_cellmath__17[23], inst_cellmath__17[22], inst_cellmath__17[21], inst_cellmath__17[20], inst_cellmath__17[19], inst_cellmath__17[18], inst_cellmath__17[17], inst_cellmath__17[16], inst_cellmath__17[15], inst_cellmath__17[14], inst_cellmath__17[13], inst_cellmath__17[12], inst_cellmath__17[11], inst_cellmath__17[10], inst_cellmath__17[9], inst_cellmath__17[8], inst_cellmath__17[7], inst_cellmath__17[6], inst_cellmath__17[5], inst_cellmath__17[4], inst_cellmath__17[3], inst_cellmath__17[2], inst_cellmath__17[1], inst_cellmath__17[0]}), .inst_cellmath__120_0_in1({inst_cellmath__16[25], inst_cellmath__16[24], inst_cellmath__16[23], inst_cellmath__16[22], inst_cellmath__16[21], inst_cellmath__16[20], inst_cellmath__16[19], inst_cellmath__16[18], inst_cellmath__16[17], inst_cellmath__16[16], inst_cellmath__16[15], inst_cellmath__16[14], inst_cellmath__16[13], inst_cellmath__16[12], inst_cellmath__16[11], inst_cellmath__16[10], inst_cellmath__16[9], inst_cellmath__16[8], inst_cellmath__16[7], inst_cellmath__16[6], inst_cellmath__16[5], inst_cellmath__16[4], inst_cellmath__16[3], inst_cellmath__16[2], inst_cellmath__16[1], 1'B0}));
DFFQXL inst_cellmath__44_0_0__I191 (.Q(inst_cellmath__44[0]), .D(inst_cellmath__40[0]), .CK(clk));
DFFQXL inst_cellmath__44_0_1__I192 (.Q(inst_cellmath__44[1]), .D(inst_cellmath__40[1]), .CK(clk));
DFFQXL inst_cellmath__44_0_2__I193 (.Q(inst_cellmath__44[2]), .D(inst_cellmath__40[2]), .CK(clk));
DFFQXL inst_cellmath__44_0_3__I194 (.Q(inst_cellmath__44[3]), .D(inst_cellmath__40[3]), .CK(clk));
DFFQXL inst_cellmath__44_0_4__I195 (.Q(inst_cellmath__44[4]), .D(inst_cellmath__40[4]), .CK(clk));
DFFQXL inst_cellmath__44_0_5__I196 (.Q(inst_cellmath__44[5]), .D(inst_cellmath__40[5]), .CK(clk));
DFFQXL inst_cellmath__44_0_6__I197 (.Q(inst_cellmath__44[6]), .D(inst_cellmath__40[6]), .CK(clk));
DFFQXL inst_cellmath__44_0_7__I198 (.Q(inst_cellmath__44[7]), .D(inst_cellmath__40[7]), .CK(clk));
DFFQXL inst_cellmath__44_0_8__I199 (.Q(inst_cellmath__44[8]), .D(inst_cellmath__40[8]), .CK(clk));
DFFQXL inst_cellmath__44_0_9__I200 (.Q(inst_cellmath__44[9]), .D(inst_cellmath__40[9]), .CK(clk));
DFFQXL inst_cellmath__44_0_10__I201 (.Q(inst_cellmath__44[10]), .D(inst_cellmath__40[10]), .CK(clk));
DFFQXL inst_cellmath__44_0_11__I202 (.Q(inst_cellmath__44[11]), .D(inst_cellmath__40[11]), .CK(clk));
DFFQXL inst_cellmath__44_0_12__I203 (.Q(inst_cellmath__44[12]), .D(inst_cellmath__40[12]), .CK(clk));
DFFQXL inst_cellmath__44_0_13__I204 (.Q(inst_cellmath__44[13]), .D(inst_cellmath__40[13]), .CK(clk));
DFFQXL inst_cellmath__44_0_14__I205 (.Q(inst_cellmath__44[14]), .D(inst_cellmath__40[14]), .CK(clk));
DFFQXL inst_cellmath__44_0_15__I206 (.Q(inst_cellmath__44[15]), .D(inst_cellmath__40[15]), .CK(clk));
DFFQXL inst_cellmath__44_0_16__I207 (.Q(inst_cellmath__44[16]), .D(inst_cellmath__40[16]), .CK(clk));
DFFQXL inst_cellmath__44_0_17__I208 (.Q(inst_cellmath__44[17]), .D(inst_cellmath__40[17]), .CK(clk));
DFFQXL inst_cellmath__44_0_18__I209 (.Q(inst_cellmath__44[18]), .D(inst_cellmath__40[18]), .CK(clk));
DFFQXL inst_cellmath__44_0_19__I210 (.Q(inst_cellmath__44[19]), .D(inst_cellmath__40[19]), .CK(clk));
DFFQXL inst_cellmath__44_0_20__I211 (.Q(inst_cellmath__44[20]), .D(inst_cellmath__40[20]), .CK(clk));
DFFQXL inst_cellmath__44_0_21__I212 (.Q(inst_cellmath__44[21]), .D(inst_cellmath__40[21]), .CK(clk));
DFFQXL inst_cellmath__44_0_22__I213 (.Q(inst_cellmath__44[22]), .D(inst_cellmath__40[22]), .CK(clk));
DFFQXL inst_cellmath__44_0_23__I214 (.Q(inst_cellmath__44[23]), .D(inst_cellmath__40[23]), .CK(clk));
DFFQXL inst_cellmath__44_0_24__I215 (.Q(inst_cellmath__44[24]), .D(inst_cellmath__40[24]), .CK(clk));
DFFQXL inst_cellmath__44_0_25__I216 (.Q(inst_cellmath__44[25]), .D(inst_cellmath__40[25]), .CK(clk));
DFFQXL inst_cellmath__44_0_26__I217 (.Q(inst_cellmath__44[26]), .D(inst_cellmath__40[26]), .CK(clk));
DFFQXL inst_cellmath__44_0_27__I218 (.Q(inst_cellmath__44[27]), .D(inst_cellmath__40[27]), .CK(clk));
DFFQXL inst_cellmath__44_0_28__I219 (.Q(inst_cellmath__44[28]), .D(inst_cellmath__40[28]), .CK(clk));
DFFQXL inst_cellmath__45_0_0__I220 (.Q(inst_cellmath__45[0]), .D(inst_cellmath__41[0]), .CK(clk));
DFFQXL inst_cellmath__45_0_1__I221 (.Q(inst_cellmath__45[1]), .D(inst_cellmath__41[1]), .CK(clk));
DFFQXL inst_cellmath__45_0_2__I222 (.Q(inst_cellmath__45[2]), .D(inst_cellmath__41[2]), .CK(clk));
DFFQXL inst_cellmath__45_0_3__I223 (.Q(inst_cellmath__45[3]), .D(inst_cellmath__41[3]), .CK(clk));
DFFQXL inst_cellmath__45_0_4__I224 (.Q(inst_cellmath__45[4]), .D(inst_cellmath__41[4]), .CK(clk));
DFFQXL inst_cellmath__45_0_5__I225 (.Q(inst_cellmath__45[5]), .D(inst_cellmath__41[5]), .CK(clk));
DFFQXL inst_cellmath__45_0_6__I226 (.Q(inst_cellmath__45[6]), .D(inst_cellmath__41[6]), .CK(clk));
DFFQXL inst_cellmath__45_0_7__I227 (.Q(inst_cellmath__45[7]), .D(inst_cellmath__41[7]), .CK(clk));
DFFQXL inst_cellmath__45_0_8__I228 (.Q(inst_cellmath__45[8]), .D(inst_cellmath__41[8]), .CK(clk));
DFFQXL inst_cellmath__45_0_9__I229 (.Q(inst_cellmath__45[9]), .D(inst_cellmath__41[9]), .CK(clk));
DFFQXL inst_cellmath__45_0_10__I230 (.Q(inst_cellmath__45[10]), .D(inst_cellmath__41[10]), .CK(clk));
DFFQXL inst_cellmath__45_0_11__I231 (.Q(inst_cellmath__45[11]), .D(inst_cellmath__41[11]), .CK(clk));
DFFQXL inst_cellmath__45_0_12__I232 (.Q(inst_cellmath__45[12]), .D(inst_cellmath__41[12]), .CK(clk));
DFFQXL inst_cellmath__45_0_13__I233 (.Q(inst_cellmath__45[13]), .D(inst_cellmath__41[13]), .CK(clk));
DFFQXL inst_cellmath__45_0_14__I234 (.Q(inst_cellmath__45[14]), .D(inst_cellmath__41[14]), .CK(clk));
DFFQXL inst_cellmath__45_0_15__I235 (.Q(inst_cellmath__45[15]), .D(inst_cellmath__41[15]), .CK(clk));
DFFQXL inst_cellmath__45_0_16__I236 (.Q(inst_cellmath__45[16]), .D(inst_cellmath__41[16]), .CK(clk));
DFFQXL inst_cellmath__45_0_17__I237 (.Q(inst_cellmath__45[17]), .D(inst_cellmath__41[17]), .CK(clk));
DFFQXL inst_cellmath__45_0_18__I238 (.Q(inst_cellmath__45[18]), .D(inst_cellmath__41[18]), .CK(clk));
DFFQXL inst_cellmath__45_0_19__I239 (.Q(inst_cellmath__45[19]), .D(inst_cellmath__41[19]), .CK(clk));
DFFQXL inst_cellmath__45_0_20__I240 (.Q(inst_cellmath__45[20]), .D(inst_cellmath__41[20]), .CK(clk));
DFFQXL inst_cellmath__45_0_21__I241 (.Q(inst_cellmath__45[21]), .D(inst_cellmath__41[21]), .CK(clk));
DFFQXL inst_cellmath__45_0_22__I242 (.Q(inst_cellmath__45[22]), .D(inst_cellmath__41[22]), .CK(clk));
DFFQXL inst_cellmath__45_0_23__I243 (.Q(inst_cellmath__45[23]), .D(inst_cellmath__41[23]), .CK(clk));
DFFQXL inst_cellmath__45_0_24__I244 (.Q(inst_cellmath__45[24]), .D(inst_cellmath__41[24]), .CK(clk));
DFFQXL inst_cellmath__45_0_25__I245 (.Q(inst_cellmath__45[25]), .D(inst_cellmath__41[25]), .CK(clk));
DFFQXL inst_cellmath__45_0_26__I246 (.Q(inst_cellmath__45[26]), .D(inst_cellmath__41[26]), .CK(clk));
DFFQXL inst_cellmath__45_0_27__I247 (.Q(inst_cellmath__45[27]), .D(inst_cellmath__41[27]), .CK(clk));
DFFQXL inst_cellmath__45_0_28__I248 (.Q(inst_cellmath__45[28]), .D(inst_cellmath__41[28]), .CK(clk));
cynw_cm_float_div_ieee_inst_cellmath__124_0_bdw410776230_bdw cynw_cm_float_div_ieee_I249 (.inst_cellmath__124_0_out0({inst_cellmath__124[28], inst_cellmath__124[27], inst_cellmath__124[26], inst_cellmath__124[25], inst_cellmath__124[24], inst_cellmath__124[23], inst_cellmath__124[22], inst_cellmath__124[21], inst_cellmath__124[20], inst_cellmath__124[19], inst_cellmath__124[18], inst_cellmath__124[17], inst_cellmath__124[16], inst_cellmath__124[15], inst_cellmath__124[14], inst_cellmath__124[13], inst_cellmath__124[12], inst_cellmath__124[11], inst_cellmath__124[10], inst_cellmath__124[9], inst_cellmath__124[8], inst_cellmath__124[7], inst_cellmath__124[6], inst_cellmath__124[5], inst_cellmath__124[4], inst_cellmath__124[3], inst_cellmath__124[2], inst_cellmath__124[1], inst_cellmath__124[0]}), .inst_cellmath__124_0_in0({inst_cellmath__45[28], inst_cellmath__45[27], inst_cellmath__45[26], inst_cellmath__45[25], inst_cellmath__45[24], inst_cellmath__45[23], inst_cellmath__45[22], inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__124_0_in1({inst_cellmath__44[28], inst_cellmath__44[27], inst_cellmath__44[26], inst_cellmath__44[25], inst_cellmath__44[24], inst_cellmath__44[23], inst_cellmath__44[22], inst_cellmath__44[21], inst_cellmath__44[20], inst_cellmath__44[19], inst_cellmath__44[18], inst_cellmath__44[17], inst_cellmath__44[16], inst_cellmath__44[15], inst_cellmath__44[14], inst_cellmath__44[13], inst_cellmath__44[12], inst_cellmath__44[11], inst_cellmath__44[10], inst_cellmath__44[9], inst_cellmath__44[8], inst_cellmath__44[7], inst_cellmath__44[6], inst_cellmath__44[5], inst_cellmath__44[4], inst_cellmath__44[3], inst_cellmath__44[2], inst_cellmath__44[1], inst_cellmath__44[0]}), .inst_cellmath__124_0_in2({inst_cellmath__120[25]}));
INVXL cynw_cm_float_div_ieee_I250 (.Y(inst_cellmath__122), .A(inst_cellmath__124[28]));
cynw_cm_float_div_ieee_inst_cellmath__125_0_bdw410776230_bdw cynw_cm_float_div_ieee_I251 (.inst_cellmath__125_0_out0({inst_cellmath__125[22], inst_cellmath__125[21], inst_cellmath__125[20], inst_cellmath__125[19], inst_cellmath__125[18], inst_cellmath__125[17], inst_cellmath__125[16], inst_cellmath__125[15], inst_cellmath__125[14], inst_cellmath__125[13], inst_cellmath__125[12], inst_cellmath__125[11], inst_cellmath__125[10], inst_cellmath__125[9], inst_cellmath__125[8], inst_cellmath__125[7], inst_cellmath__125[6], inst_cellmath__125[5], inst_cellmath__125[4], inst_cellmath__125[3], inst_cellmath__125[2], inst_cellmath__125[1], inst_cellmath__125[0]}), .inst_cellmath__125_0_in0({inst_cellmath__124[27], inst_cellmath__124[26], inst_cellmath__124[25], inst_cellmath__124[24], inst_cellmath__124[23], inst_cellmath__124[22], inst_cellmath__124[21], inst_cellmath__124[20], inst_cellmath__124[19], inst_cellmath__124[18], inst_cellmath__124[17], inst_cellmath__124[16], inst_cellmath__124[15], inst_cellmath__124[14], inst_cellmath__124[13], inst_cellmath__124[12], inst_cellmath__124[11], inst_cellmath__124[10], inst_cellmath__124[9], inst_cellmath__124[8], inst_cellmath__124[7], inst_cellmath__124[6], inst_cellmath__124[5], inst_cellmath__124[4]}), .inst_cellmath__125_0_in1(inst_cellmath__122));
cynw_cm_float_div_ieee_inst_cellmath__126_0_bdw410776230_bdw cynw_cm_float_div_ieee_I252 (.inst_cellmath__126_0_out0(inst_cellmath__126), .inst_cellmath__126_0_in0({inst_cellmath__124[4], inst_cellmath__124[3]}), .inst_cellmath__126_0_in1(inst_cellmath__122));
cynw_cm_float_div_ieee_inst_cellmath__129_0_bdw410776230_bdw cynw_cm_float_div_ieee_I253 (.inst_cellmath__129_0_out0({inst_cellmath__129[22], inst_cellmath__129[21], inst_cellmath__129[20], inst_cellmath__129[19], inst_cellmath__129[18], inst_cellmath__129[17], inst_cellmath__129[16], inst_cellmath__129[15], inst_cellmath__129[14], inst_cellmath__129[13], inst_cellmath__129[12], inst_cellmath__129[11], inst_cellmath__129[10], inst_cellmath__129[9], inst_cellmath__129[8], inst_cellmath__129[7], inst_cellmath__129[6], inst_cellmath__129[5], inst_cellmath__129[4], inst_cellmath__129[3], inst_cellmath__129[2], inst_cellmath__129[1], inst_cellmath__129[0]}), .inst_cellmath__129_0_in0(inst_cellmath__126), .inst_cellmath__129_0_in1({inst_cellmath__125[22], inst_cellmath__125[21], inst_cellmath__125[20], inst_cellmath__125[19], inst_cellmath__125[18], inst_cellmath__125[17], inst_cellmath__125[16], inst_cellmath__125[15], inst_cellmath__125[14], inst_cellmath__125[13], inst_cellmath__125[12], inst_cellmath__125[11], inst_cellmath__125[10], inst_cellmath__125[9], inst_cellmath__125[8], inst_cellmath__125[7], inst_cellmath__125[6], inst_cellmath__125[5], inst_cellmath__125[4], inst_cellmath__125[3], inst_cellmath__125[2], inst_cellmath__125[1], inst_cellmath__125[0]}));
cynw_cm_float_div_ieee_inst_cellmath__127__104__bdw410776230_bdw cynw_cm_float_div_ieee_I254 (.inst_cellmath__127__104__out0({N1682}), .inst_cellmath__127__104__in0({inst_cellmath__124[3], inst_cellmath__124[2], inst_cellmath__124[1], inst_cellmath__124[0]}));
cynw_cm_float_div_ieee_inst_cellmath__127__103__bdw410776230_bdw cynw_cm_float_div_ieee_I255 (.inst_cellmath__127__103__out0({N1681}), .inst_cellmath__127__103__in0({inst_cellmath__124[2], inst_cellmath__124[1], inst_cellmath__124[0]}));
cynw_cm_float_div_ieee_inst_cellmath__127_0_bdw410776230_bdw cynw_cm_float_div_ieee_I256 (.inst_cellmath__127_0_out0(inst_cellmath__127), .inst_cellmath__127_0_in0({N1682}), .inst_cellmath__127_0_in1({N1681}), .inst_cellmath__127_0_in2(inst_cellmath__122));
cynw_cm_float_div_ieee_inst_cellmath__130__105__bdw410776230_bdw cynw_cm_float_div_ieee_I257 (.inst_cellmath__130__105__out0({N1683}), .inst_cellmath__130__105__in0(inst_cellmath__127), .inst_cellmath__130__105__in1({inst_cellmath__125[0]}), .inst_cellmath__130__105__in2({inst_cellmath__120[25], inst_cellmath__120[24], inst_cellmath__120[23], inst_cellmath__120[22], inst_cellmath__120[21], inst_cellmath__120[20], inst_cellmath__120[19], inst_cellmath__120[18], inst_cellmath__120[17], inst_cellmath__120[16], inst_cellmath__120[15], inst_cellmath__120[14], inst_cellmath__120[13], inst_cellmath__120[12], inst_cellmath__120[11], inst_cellmath__120[10], inst_cellmath__120[9], inst_cellmath__120[8], inst_cellmath__120[7], inst_cellmath__120[6], inst_cellmath__120[5], inst_cellmath__120[4], inst_cellmath__120[3], inst_cellmath__120[2], inst_cellmath__120[1], inst_cellmath__120[0]}));
cynw_cm_float_div_ieee_inst_cellmath__121__106__bdw410776230_bdw cynw_cm_float_div_ieee_I258 (.inst_cellmath__121__106__out0({N1922}), .inst_cellmath__121__106__in0({N1683}), .inst_cellmath__121__106__in1({inst_cellmath__129[0]}));
INVXL cynw_cm_float_div_ieee_I259 (.Y(N1322), .A(accept));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_0__I260 (.q(inst_cellmath__13[0]), .r(N1322), .d(inst_cellmath__12[0]), .clk(clk));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_1__I261 (.q(inst_cellmath__13[1]), .r(N1322), .d(inst_cellmath__12[1]), .clk(clk));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_2__I262 (.q(inst_cellmath__13[2]), .r(N1322), .d(inst_cellmath__12[2]), .clk(clk));
arith_fdrq_A_bdw410776230_bdw inst_cellmath__13_0_3__I263 (.q(inst_cellmath__13[3]), .r(N1322), .d(inst_cellmath__12[3]), .clk(clk));
cynw_cm_float_div_ieee_inst_cellmath__12__18__bdw410776230_bdw cynw_cm_float_div_ieee_I264 (.inst_cellmath__12__18__out0({N1326, N1325, N1324, N1323}), .inst_cellmath__12__18__in0({inst_cellmath__13[3], inst_cellmath__13[2], inst_cellmath__13[1], inst_cellmath__13[0]}));
cynw_cm_float_div_ieee_inst_cellmath__12__19__bdw410776230_bdw cynw_cm_float_div_ieee_I265 (.inst_cellmath__12__19__out0({N1327}), .inst_cellmath__12__19__in0({inst_cellmath__13[3], inst_cellmath__13[2], inst_cellmath__13[1], inst_cellmath__13[0]}));
cynw_cm_float_div_ieee_inst_cellmath__12_0_bdw410776230_bdw cynw_cm_float_div_ieee_I266 (.inst_cellmath__12_0_out0({inst_cellmath__12[3], inst_cellmath__12[2], inst_cellmath__12[1], inst_cellmath__12[0]}), .inst_cellmath__12_0_in0({N1327}), .inst_cellmath__12_0_in1({N1326, N1325, N1324, N1323}));
cynw_cm_float_div_ieee_inst_cellmath__46_0_bdw410776230_bdw cynw_cm_float_div_ieee_I267 (.inst_cellmath__46_0_out0({inst_cellmath__46[24], inst_cellmath__46[23], inst_cellmath__46[22], inst_cellmath__46[21], inst_cellmath__46[20], inst_cellmath__46[19], inst_cellmath__46[18], inst_cellmath__46[17], inst_cellmath__46[16], inst_cellmath__46[15], inst_cellmath__46[14], inst_cellmath__46[13], inst_cellmath__46[12], inst_cellmath__46[11], inst_cellmath__46[10], inst_cellmath__46[9], inst_cellmath__46[8], inst_cellmath__46[7], inst_cellmath__46[6], inst_cellmath__46[5], inst_cellmath__46[4], inst_cellmath__46[3], inst_cellmath__46[2], inst_cellmath__46[1], inst_cellmath__46[0]}), .inst_cellmath__46_0_in0({inst_cellmath__44[24], inst_cellmath__44[23], inst_cellmath__44[22], inst_cellmath__44[21], inst_cellmath__44[20], inst_cellmath__44[19], inst_cellmath__44[18], inst_cellmath__44[17], inst_cellmath__44[16], inst_cellmath__44[15], inst_cellmath__44[14], inst_cellmath__44[13], inst_cellmath__44[12], inst_cellmath__44[11], inst_cellmath__44[10], inst_cellmath__44[9], inst_cellmath__44[8], inst_cellmath__44[7], inst_cellmath__44[6], inst_cellmath__44[5], inst_cellmath__44[4], inst_cellmath__44[3], inst_cellmath__44[2], inst_cellmath__44[1], inst_cellmath__44[0]}), .inst_cellmath__46_0_in1(inst_cellmath__11));
cynw_cm_float_div_ieee_inst_cellmath__47_0_bdw410776230_bdw cynw_cm_float_div_ieee_I268 (.inst_cellmath__47_0_out0({inst_cellmath__47[24], inst_cellmath__47[23], inst_cellmath__47[22], inst_cellmath__47[21], inst_cellmath__47[20], inst_cellmath__47[19], inst_cellmath__47[18], inst_cellmath__47[17], inst_cellmath__47[16], inst_cellmath__47[15], inst_cellmath__47[14], inst_cellmath__47[13], inst_cellmath__47[12], inst_cellmath__47[11], inst_cellmath__47[10], inst_cellmath__47[9], inst_cellmath__47[8], inst_cellmath__47[7], inst_cellmath__47[6], inst_cellmath__47[5], inst_cellmath__47[4], inst_cellmath__47[3], inst_cellmath__47[2], inst_cellmath__47[1], inst_cellmath__47[0]}), .inst_cellmath__47_0_in0({inst_cellmath__45[24], inst_cellmath__45[23], inst_cellmath__45[22], inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__47_0_in1(inst_cellmath__11));
cynw_cm_float_div_ieee_inst_cellmath__48__47__bdw410776230_bdw cynw_cm_float_div_ieee_I269 (.inst_cellmath__48__47__out0({N1417}), .inst_cellmath__48__47__in0({inst_lookup0_cellmath__29[1], inst_lookup0_cellmath__29[0]}));
cynw_cm_float_div_ieee_inst_cellmath__48__44__bdw410776230_bdw cynw_cm_float_div_ieee_I270 (.inst_cellmath__48__44__out0({N1447}), .inst_cellmath__48__44__in0({inst_lookup0_cellmath__29[2], inst_lookup0_cellmath__29[1]}), .inst_cellmath__48__44__in1({N1417}));
cynw_cm_float_div_ieee_inst_cellmath__42_0_bdw410776230_bdw cynw_cm_float_div_ieee_I271 (.inst_cellmath__42_0_out0({inst_cellmath__42[26], inst_cellmath__42[25], inst_cellmath__42[24], inst_cellmath__42[23], inst_cellmath__42[22], inst_cellmath__42[21], inst_cellmath__42[20], inst_cellmath__42[19], inst_cellmath__42[18], inst_cellmath__42[17], inst_cellmath__42[16], inst_cellmath__42[15], inst_cellmath__42[14], inst_cellmath__42[13], inst_cellmath__42[12], inst_cellmath__42[11], inst_cellmath__42[10], inst_cellmath__42[9], inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6], inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__42_0_in0({inst_lookup0_cellmath__29[0]}), .inst_cellmath__42_0_in1({N1447}), .inst_cellmath__42_0_in2({inst_cellmath__47[24], inst_cellmath__47[23], inst_cellmath__47[22], inst_cellmath__47[21], inst_cellmath__47[20], inst_cellmath__47[19], inst_cellmath__47[18], inst_cellmath__47[17], inst_cellmath__47[16], inst_cellmath__47[15], inst_cellmath__47[14], inst_cellmath__47[13], inst_cellmath__47[12], inst_cellmath__47[11], inst_cellmath__47[10], inst_cellmath__47[9], inst_cellmath__47[8], inst_cellmath__47[7], inst_cellmath__47[6], inst_cellmath__47[5], inst_cellmath__47[4], inst_cellmath__47[3], inst_cellmath__47[2], inst_cellmath__47[1], inst_cellmath__47[0]}), .inst_cellmath__42_0_in3({inst_cellmath__46[24], inst_cellmath__46[23], inst_cellmath__46[22], inst_cellmath__46[21], inst_cellmath__46[20], inst_cellmath__46[19], inst_cellmath__46[18], inst_cellmath__46[17], inst_cellmath__46[16], inst_cellmath__46[15], inst_cellmath__46[14], inst_cellmath__46[13], inst_cellmath__46[12], inst_cellmath__46[11], inst_cellmath__46[10], inst_cellmath__46[9], inst_cellmath__46[8], inst_cellmath__46[7], inst_cellmath__46[6], inst_cellmath__46[5], inst_cellmath__46[4], inst_cellmath__46[3], inst_cellmath__46[2], inst_cellmath__46[1], inst_cellmath__46[0]}), .inst_cellmath__42_0_in4(inst_cellmath__35[0]));
cynw_cm_float_div_ieee_inst_cellmath__50_0_bdw410776230_bdw cynw_cm_float_div_ieee_I272 (.inst_cellmath__50_0_out0({inst_cellmath__50[1], inst_cellmath__50[0]}), .inst_cellmath__50_0_in0({inst_lookup0_cellmath__29[0]}), .inst_cellmath__50_0_in1({N1447}));
cynw_cm_float_div_ieee_inst_cellmath__43__56__bdw410776230_bdw cynw_cm_float_div_ieee_I273 (.inst_cellmath__43__56__out0({N1527}), .inst_cellmath__43__56__in0({inst_lookup0_cellmath__29[0]}), .inst_cellmath__43__56__in1({N1447}));
cynw_cm_float_div_ieee_inst_cellmath__43__55__bdw410776230_bdw cynw_cm_float_div_ieee_I274 (.inst_cellmath__43__55__out0({N1528}), .inst_cellmath__43__55__in0({inst_lookup0_cellmath__29[2]}), .inst_cellmath__43__55__in1({N1527}));
cynw_cm_float_div_ieee_inst_cellmath__43_0_bdw410776230_bdw cynw_cm_float_div_ieee_I275 (.inst_cellmath__43_0_out0({inst_cellmath__43[26], inst_cellmath__43[25], inst_cellmath__43[24], inst_cellmath__43[23], inst_cellmath__43[22], inst_cellmath__43[21], inst_cellmath__43[20], inst_cellmath__43[19], inst_cellmath__43[18], inst_cellmath__43[17], inst_cellmath__43[16], inst_cellmath__43[15], inst_cellmath__43[14], inst_cellmath__43[13], inst_cellmath__43[12], inst_cellmath__43[11], inst_cellmath__43[10], inst_cellmath__43[9], inst_cellmath__43[8], inst_cellmath__43[7], inst_cellmath__43[6], inst_cellmath__43[5], inst_cellmath__43[4], inst_cellmath__43[3], inst_cellmath__43[2], inst_cellmath__43[1], inst_cellmath__43[0]}), .inst_cellmath__43_0_in0({inst_cellmath__50[1], inst_cellmath__50[0]}), .inst_cellmath__43_0_in1({inst_cellmath__47[24], inst_cellmath__47[23], inst_cellmath__47[22], inst_cellmath__47[21], inst_cellmath__47[20], inst_cellmath__47[19], inst_cellmath__47[18], inst_cellmath__47[17], inst_cellmath__47[16], inst_cellmath__47[15], inst_cellmath__47[14], inst_cellmath__47[13], inst_cellmath__47[12], inst_cellmath__47[11], inst_cellmath__47[10], inst_cellmath__47[9], inst_cellmath__47[8], inst_cellmath__47[7], inst_cellmath__47[6], inst_cellmath__47[5], inst_cellmath__47[4], inst_cellmath__47[3], inst_cellmath__47[2], inst_cellmath__47[1], inst_cellmath__47[0]}), .inst_cellmath__43_0_in2({inst_cellmath__46[24], inst_cellmath__46[23], inst_cellmath__46[22], inst_cellmath__46[21], inst_cellmath__46[20], inst_cellmath__46[19], inst_cellmath__46[18], inst_cellmath__46[17], inst_cellmath__46[16], inst_cellmath__46[15], inst_cellmath__46[14], inst_cellmath__46[13], inst_cellmath__46[12], inst_cellmath__46[11], inst_cellmath__46[10], inst_cellmath__46[9], inst_cellmath__46[8], inst_cellmath__46[7], inst_cellmath__46[6], inst_cellmath__46[5], inst_cellmath__46[4], inst_cellmath__46[3], inst_cellmath__46[2], inst_cellmath__46[1], inst_cellmath__46[0]}), .inst_cellmath__43_0_in3({N1528}));
cynw_cm_float_div_ieee_inst_it2_cellmath__56_2mx_bdw410776230_bdw cynw_cm_float_div_ieee_I276 (.inst_it2_cellmath__56_2mx_out0({inst_it2_cellmath__56[25], inst_it2_cellmath__56[24], inst_it2_cellmath__56[23], inst_it2_cellmath__56[22], inst_it2_cellmath__56[21], inst_it2_cellmath__56[20], inst_it2_cellmath__56[19], inst_it2_cellmath__56[18], inst_it2_cellmath__56[17], inst_it2_cellmath__56[16], inst_it2_cellmath__56[15], inst_it2_cellmath__56[14], inst_it2_cellmath__56[13], inst_it2_cellmath__56[12], inst_it2_cellmath__56[11], inst_it2_cellmath__56[10], inst_it2_cellmath__56[9], inst_it2_cellmath__56[8], inst_it2_cellmath__56[7], inst_it2_cellmath__56[6], inst_it2_cellmath__56[5], inst_it2_cellmath__56[4], inst_it2_cellmath__56[3], inst_it2_cellmath__56[2], inst_it2_cellmath__56[1], inst_it2_cellmath__56[0]}), .inst_it2_cellmath__56_2mx_in0({inst_it2_lookup1_cellmath__55[2]}), .inst_it2_cellmath__56_2mx_in1({N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201}));
cynw_cm_float_div_ieee_inst_it2_cellmath__57_2mx_bdw410776230_bdw cynw_cm_float_div_ieee_I277 (.inst_it2_cellmath__57_2mx_out0({inst_it2_cellmath__57[25], inst_it2_cellmath__57[24], inst_it2_cellmath__57[23], inst_it2_cellmath__57[22], inst_it2_cellmath__57[21], inst_it2_cellmath__57[20], inst_it2_cellmath__57[19], inst_it2_cellmath__57[18], inst_it2_cellmath__57[17], inst_it2_cellmath__57[16], inst_it2_cellmath__57[15], inst_it2_cellmath__57[14], inst_it2_cellmath__57[13], inst_it2_cellmath__57[12], inst_it2_cellmath__57[11], inst_it2_cellmath__57[10], inst_it2_cellmath__57[9], inst_it2_cellmath__57[8], inst_it2_cellmath__57[7], inst_it2_cellmath__57[6], inst_it2_cellmath__57[5], inst_it2_cellmath__57[4], inst_it2_cellmath__57[3], inst_it2_cellmath__57[2], inst_it2_cellmath__57[1], inst_it2_cellmath__57[0]}), .inst_it2_cellmath__57_2mx_in0({inst_it2_lookup1_cellmath__55[2]}), .inst_it2_cellmath__57_2mx_in1({N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254}));
INVXL cynw_cm_float_div_ieee_I278 (.Y(inst_it2_cellmath__61[0]), .A(inst_it2_lookup1_cellmath__55[2]));
cynw_cm_float_div_ieee_inst_fa_1820_10_bdw410776230_bdw cynw_cm_float_div_ieee_I279 (.inst_fa_1820_10_out0({inst_it2_cellmath__62__W1[25], inst_it2_cellmath__62__W1[24], inst_it2_cellmath__62__W1[23], inst_it2_cellmath__62__W1[22], inst_it2_cellmath__62__W1[21], inst_it2_cellmath__62__W1[20], inst_it2_cellmath__62__W1[19], inst_it2_cellmath__62__W1[18], inst_it2_cellmath__62__W1[17], inst_it2_cellmath__62__W1[16], inst_it2_cellmath__62__W1[15], inst_it2_cellmath__62__W1[14], inst_it2_cellmath__62__W1[13], inst_it2_cellmath__62__W1[12], inst_it2_cellmath__62__W1[11], inst_it2_cellmath__62__W1[10], inst_it2_cellmath__62__W1[9], inst_it2_cellmath__62__W1[8], inst_it2_cellmath__62__W1[7], inst_it2_cellmath__62__W1[6], inst_it2_cellmath__62__W1[5], inst_it2_cellmath__62__W1[4], inst_it2_cellmath__62__W1[3], inst_it2_cellmath__62__W1[2], inst_it2_cellmath__62__W1[1], inst_it2_cellmath__62__W1[0]}), .inst_fa_1820_10_out1({inst_it2_cellmath__62__W0[24], inst_it2_cellmath__62__W0[23], inst_it2_cellmath__62__W0[22], inst_it2_cellmath__62__W0[21], inst_it2_cellmath__62__W0[20], inst_it2_cellmath__62__W0[19], inst_it2_cellmath__62__W0[18], inst_it2_cellmath__62__W0[17], inst_it2_cellmath__62__W0[16], inst_it2_cellmath__62__W0[15], inst_it2_cellmath__62__W0[14], inst_it2_cellmath__62__W0[13], inst_it2_cellmath__62__W0[12], inst_it2_cellmath__62__W0[11], inst_it2_cellmath__62__W0[10], inst_it2_cellmath__62__W0[9], inst_it2_cellmath__62__W0[8], inst_it2_cellmath__62__W0[7], inst_it2_cellmath__62__W0[6], inst_it2_cellmath__62__W0[5], inst_it2_cellmath__62__W0[4], inst_it2_cellmath__62__W0[3], inst_it2_cellmath__62__W0[2], inst_it2_cellmath__62__W0[1], inst_it2_cellmath__62__W0[0]}), .inst_fa_1820_10_in0(inst_it2_cellmath__61[0]), .inst_fa_1820_10_in1({inst_it2_cellmath__56[25], inst_it2_cellmath__56[24], inst_it2_cellmath__56[23], inst_it2_cellmath__56[22], inst_it2_cellmath__56[21], inst_it2_cellmath__56[20], inst_it2_cellmath__56[19], inst_it2_cellmath__56[18], inst_it2_cellmath__56[17], inst_it2_cellmath__56[16], inst_it2_cellmath__56[15], inst_it2_cellmath__56[14], inst_it2_cellmath__56[13], inst_it2_cellmath__56[12], inst_it2_cellmath__56[11], inst_it2_cellmath__56[10], inst_it2_cellmath__56[9], inst_it2_cellmath__56[8], inst_it2_cellmath__56[7], inst_it2_cellmath__56[6], inst_it2_cellmath__56[5], inst_it2_cellmath__56[4], inst_it2_cellmath__56[3], inst_it2_cellmath__56[2], inst_it2_cellmath__56[1], inst_it2_cellmath__56[0]}), .inst_fa_1820_10_in2({inst_it2_cellmath__61[25], inst_it2_cellmath__61[24], inst_it2_cellmath__61[23], inst_it2_cellmath__61[22], inst_it2_cellmath__61[21], inst_it2_cellmath__61[20], inst_it2_cellmath__61[19], inst_it2_cellmath__61[18], inst_it2_cellmath__61[17], inst_it2_cellmath__61[16], inst_it2_cellmath__61[15], inst_it2_cellmath__61[14], inst_it2_cellmath__61[13], inst_it2_cellmath__61[12], inst_it2_cellmath__61[11], inst_it2_cellmath__61[10], inst_it2_cellmath__61[9], inst_it2_cellmath__61[8], inst_it2_cellmath__61[7], inst_it2_cellmath__61[6], inst_it2_cellmath__61[5], inst_it2_cellmath__61[4], inst_it2_cellmath__61[3], inst_it2_cellmath__61[2]}), .inst_fa_1820_10_in3({inst_it2_cellmath__60[25], inst_it2_cellmath__60[24], inst_it2_cellmath__60[23], inst_it2_cellmath__60[22], inst_it2_cellmath__60[21], inst_it2_cellmath__60[20], inst_it2_cellmath__60[19], inst_it2_cellmath__60[18], inst_it2_cellmath__60[17], inst_it2_cellmath__60[16], inst_it2_cellmath__60[15], inst_it2_cellmath__60[14], inst_it2_cellmath__60[13], inst_it2_cellmath__60[12], inst_it2_cellmath__60[11], inst_it2_cellmath__60[10], inst_it2_cellmath__60[9], inst_it2_cellmath__60[8], inst_it2_cellmath__60[7], inst_it2_cellmath__60[6], inst_it2_cellmath__60[5], inst_it2_cellmath__60[4], inst_it2_cellmath__60[3]}));
cynw_cm_float_div_ieee_inst_fa_1839_10_bdw410776230_bdw cynw_cm_float_div_ieee_I280 (.inst_fa_1839_10_out0({inst_it2_cellmath__63__W1[25], inst_it2_cellmath__63__W1[24], inst_it2_cellmath__63__W1[23], inst_it2_cellmath__63__W1[22], inst_it2_cellmath__63__W1[21], inst_it2_cellmath__63__W1[20], inst_it2_cellmath__63__W1[19], inst_it2_cellmath__63__W1[18], inst_it2_cellmath__63__W1[17], inst_it2_cellmath__63__W1[16], inst_it2_cellmath__63__W1[15], inst_it2_cellmath__63__W1[14], inst_it2_cellmath__63__W1[13], inst_it2_cellmath__63__W1[12], inst_it2_cellmath__63__W1[11], inst_it2_cellmath__63__W1[10], inst_it2_cellmath__63__W1[9], inst_it2_cellmath__63__W1[8], inst_it2_cellmath__63__W1[7], inst_it2_cellmath__63__W1[6], inst_it2_cellmath__63__W1[5], inst_it2_cellmath__63__W1[4], inst_it2_cellmath__63__W1[3], inst_it2_cellmath__63__W1[2], inst_it2_cellmath__63__W1[1], inst_it2_cellmath__63__W1[0]}), .inst_fa_1839_10_out1({inst_cellmath__14[25], inst_cellmath__14[24], inst_cellmath__14[23], inst_cellmath__14[22], inst_cellmath__14[21], inst_cellmath__14[20], inst_cellmath__14[19], inst_cellmath__14[18], inst_cellmath__14[17], inst_cellmath__14[16], inst_cellmath__14[15], inst_cellmath__14[14], inst_cellmath__14[13], inst_cellmath__14[12], inst_cellmath__14[11], inst_cellmath__14[10], inst_cellmath__14[9], inst_cellmath__14[8], inst_cellmath__14[7], inst_cellmath__14[6], inst_cellmath__14[5], inst_cellmath__14[4], inst_cellmath__14[3], inst_cellmath__14[2], inst_cellmath__14[1]}), .inst_fa_1839_10_in0({inst_it2_cellmath__62__W1[25], inst_it2_cellmath__62__W1[24], inst_it2_cellmath__62__W1[23], inst_it2_cellmath__62__W1[22], inst_it2_cellmath__62__W1[21], inst_it2_cellmath__62__W1[20], inst_it2_cellmath__62__W1[19], inst_it2_cellmath__62__W1[18], inst_it2_cellmath__62__W1[17], inst_it2_cellmath__62__W1[16], inst_it2_cellmath__62__W1[15], inst_it2_cellmath__62__W1[14], inst_it2_cellmath__62__W1[13], inst_it2_cellmath__62__W1[12], inst_it2_cellmath__62__W1[11], inst_it2_cellmath__62__W1[10], inst_it2_cellmath__62__W1[9], inst_it2_cellmath__62__W1[8], inst_it2_cellmath__62__W1[7], inst_it2_cellmath__62__W1[6], inst_it2_cellmath__62__W1[5], inst_it2_cellmath__62__W1[4], inst_it2_cellmath__62__W1[3], inst_it2_cellmath__62__W1[2], inst_it2_cellmath__62__W1[1], inst_it2_cellmath__62__W1[0]}), .inst_fa_1839_10_in1({inst_it2_cellmath__62__W0[24], inst_it2_cellmath__62__W0[23], inst_it2_cellmath__62__W0[22], inst_it2_cellmath__62__W0[21], inst_it2_cellmath__62__W0[20], inst_it2_cellmath__62__W0[19], inst_it2_cellmath__62__W0[18], inst_it2_cellmath__62__W0[17], inst_it2_cellmath__62__W0[16], inst_it2_cellmath__62__W0[15], inst_it2_cellmath__62__W0[14], inst_it2_cellmath__62__W0[13], inst_it2_cellmath__62__W0[12], inst_it2_cellmath__62__W0[11], inst_it2_cellmath__62__W0[10], inst_it2_cellmath__62__W0[9], inst_it2_cellmath__62__W0[8], inst_it2_cellmath__62__W0[7], inst_it2_cellmath__62__W0[6], inst_it2_cellmath__62__W0[5], inst_it2_cellmath__62__W0[4], inst_it2_cellmath__62__W0[3], inst_it2_cellmath__62__W0[2], inst_it2_cellmath__62__W0[1], inst_it2_cellmath__62__W0[0]}), .inst_fa_1839_10_in2({inst_it2_cellmath__57[25], inst_it2_cellmath__57[24], inst_it2_cellmath__57[23], inst_it2_cellmath__57[22], inst_it2_cellmath__57[21], inst_it2_cellmath__57[20], inst_it2_cellmath__57[19], inst_it2_cellmath__57[18], inst_it2_cellmath__57[17], inst_it2_cellmath__57[16], inst_it2_cellmath__57[15], inst_it2_cellmath__57[14], inst_it2_cellmath__57[13], inst_it2_cellmath__57[12], inst_it2_cellmath__57[11], inst_it2_cellmath__57[10], inst_it2_cellmath__57[9], inst_it2_cellmath__57[8], inst_it2_cellmath__57[7], inst_it2_cellmath__57[6], inst_it2_cellmath__57[5], inst_it2_cellmath__57[4], inst_it2_cellmath__57[3], inst_it2_cellmath__57[2], inst_it2_cellmath__57[1], inst_it2_cellmath__57[0]}));
cynw_cm_float_div_ieee_inst_it2_cellmath__64__71__bdw410776230_bdw cynw_cm_float_div_ieee_I281 (.inst_it2_cellmath__64__71__out0({N1555}), .inst_it2_cellmath__64__71__in0({inst_it2_lookup1_cellmath__55[1], inst_it2_lookup1_cellmath__55[0]}));
cynw_cm_float_div_ieee_inst_it2_cellmath__64__68__bdw410776230_bdw cynw_cm_float_div_ieee_I282 (.inst_it2_cellmath__64__68__out0({N1587}), .inst_it2_cellmath__64__68__in0({inst_it2_lookup1_cellmath__55[2], inst_it2_lookup1_cellmath__55[1]}), .inst_it2_cellmath__64__68__in1({N1555}));
cynw_cm_float_div_ieee_inst_cellmath__40_0_bdw410776230_bdw cynw_cm_float_div_ieee_I283 (.inst_cellmath__40_0_out0({inst_cellmath__40[28], inst_cellmath__40[27], inst_cellmath__40[26], inst_cellmath__40[25], inst_cellmath__40[24], inst_cellmath__40[23], inst_cellmath__40[22], inst_cellmath__40[21], inst_cellmath__40[20], inst_cellmath__40[19], inst_cellmath__40[18], inst_cellmath__40[17], inst_cellmath__40[16], inst_cellmath__40[15], inst_cellmath__40[14], inst_cellmath__40[13], inst_cellmath__40[12], inst_cellmath__40[11], inst_cellmath__40[10], inst_cellmath__40[9], inst_cellmath__40[8], inst_cellmath__40[7], inst_cellmath__40[6], inst_cellmath__40[5], inst_cellmath__40[4], inst_cellmath__40[3], inst_cellmath__40[2], inst_cellmath__40[1], inst_cellmath__40[0]}), .inst_cellmath__40_0_in0({inst_it2_lookup1_cellmath__55[0]}), .inst_cellmath__40_0_in1({N1587}), .inst_cellmath__40_0_in2(inst_it2_cellmath__61[0]), .inst_cellmath__40_0_in3({inst_cellmath__43[26], inst_cellmath__43[25], inst_cellmath__43[24], inst_cellmath__43[23], inst_cellmath__43[22], inst_cellmath__43[21], inst_cellmath__43[20], inst_cellmath__43[19], inst_cellmath__43[18], inst_cellmath__43[17], inst_cellmath__43[16], inst_cellmath__43[15], inst_cellmath__43[14], inst_cellmath__43[13], inst_cellmath__43[12], inst_cellmath__43[11], inst_cellmath__43[10], inst_cellmath__43[9], inst_cellmath__43[8], inst_cellmath__43[7], inst_cellmath__43[6], inst_cellmath__43[5], inst_cellmath__43[4], inst_cellmath__43[3], inst_cellmath__43[2], inst_cellmath__43[1], inst_cellmath__43[0]}), .inst_cellmath__40_0_in4({inst_cellmath__42[26], inst_cellmath__42[25], inst_cellmath__42[24], inst_cellmath__42[23], inst_cellmath__42[22], inst_cellmath__42[21], inst_cellmath__42[20], inst_cellmath__42[19], inst_cellmath__42[18], inst_cellmath__42[17], inst_cellmath__42[16], inst_cellmath__42[15], inst_cellmath__42[14], inst_cellmath__42[13], inst_cellmath__42[12], inst_cellmath__42[11], inst_cellmath__42[10], inst_cellmath__42[9], inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6], inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}));
cynw_cm_float_div_ieee_inst_it2_cellmath__66_0_bdw410776230_bdw cynw_cm_float_div_ieee_I284 (.inst_it2_cellmath__66_0_out0({inst_it2_cellmath__66[1], inst_it2_cellmath__66[0]}), .inst_it2_cellmath__66_0_in0({inst_it2_lookup1_cellmath__55[0]}), .inst_it2_cellmath__66_0_in1({N1587}));
cynw_cm_float_div_ieee_inst_cellmath__41__80__bdw410776230_bdw cynw_cm_float_div_ieee_I285 (.inst_cellmath__41__80__out0({N1673}), .inst_cellmath__41__80__in0({inst_it2_lookup1_cellmath__55[0]}), .inst_cellmath__41__80__in1({N1587}));
cynw_cm_float_div_ieee_inst_cellmath__41__79__bdw410776230_bdw cynw_cm_float_div_ieee_I286 (.inst_cellmath__41__79__out0({N1674}), .inst_cellmath__41__79__in0({inst_it2_lookup1_cellmath__55[2]}), .inst_cellmath__41__79__in1({N1673}));
cynw_cm_float_div_ieee_inst_cellmath__41_0_bdw410776230_bdw cynw_cm_float_div_ieee_I287 (.inst_cellmath__41_0_out0({inst_cellmath__41[28], inst_cellmath__41[27], inst_cellmath__41[26], inst_cellmath__41[25], inst_cellmath__41[24], inst_cellmath__41[23], inst_cellmath__41[22], inst_cellmath__41[21], inst_cellmath__41[20], inst_cellmath__41[19], inst_cellmath__41[18], inst_cellmath__41[17], inst_cellmath__41[16], inst_cellmath__41[15], inst_cellmath__41[14], inst_cellmath__41[13], inst_cellmath__41[12], inst_cellmath__41[11], inst_cellmath__41[10], inst_cellmath__41[9], inst_cellmath__41[8], inst_cellmath__41[7], inst_cellmath__41[6], inst_cellmath__41[5], inst_cellmath__41[4], inst_cellmath__41[3], inst_cellmath__41[2], inst_cellmath__41[1], inst_cellmath__41[0]}), .inst_cellmath__41_0_in0({inst_it2_cellmath__66[1], inst_it2_cellmath__66[0]}), .inst_cellmath__41_0_in1({inst_cellmath__43[26], inst_cellmath__43[25], inst_cellmath__43[24], inst_cellmath__43[23], inst_cellmath__43[22], inst_cellmath__43[21], inst_cellmath__43[20], inst_cellmath__43[19], inst_cellmath__43[18], inst_cellmath__43[17], inst_cellmath__43[16], inst_cellmath__43[15], inst_cellmath__43[14], inst_cellmath__43[13], inst_cellmath__43[12], inst_cellmath__43[11], inst_cellmath__43[10], inst_cellmath__43[9], inst_cellmath__43[8], inst_cellmath__43[7], inst_cellmath__43[6], inst_cellmath__43[5], inst_cellmath__43[4], inst_cellmath__43[3], inst_cellmath__43[2], inst_cellmath__43[1], inst_cellmath__43[0]}), .inst_cellmath__41_0_in2({inst_cellmath__42[26], inst_cellmath__42[25], inst_cellmath__42[24], inst_cellmath__42[23], inst_cellmath__42[22], inst_cellmath__42[21], inst_cellmath__42[20], inst_cellmath__42[19], inst_cellmath__42[18], inst_cellmath__42[17], inst_cellmath__42[16], inst_cellmath__42[15], inst_cellmath__42[14], inst_cellmath__42[13], inst_cellmath__42[12], inst_cellmath__42[11], inst_cellmath__42[10], inst_cellmath__42[9], inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6], inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__41_0_in3({N1674}));
cynw_cm_float_div_ieee_inst_cellmath__67_0_bdw410776230_bdw cynw_cm_float_div_ieee_I288 (.inst_cellmath__67_0_out0({inst_cellmath__67[7], inst_cellmath__67[6], inst_cellmath__67[5], inst_cellmath__67[4], inst_cellmath__67[3], inst_cellmath__67[2], inst_cellmath__67[1], inst_cellmath__67[0]}), .inst_cellmath__67_0_in0({inst_cellmath__9[30], inst_cellmath__9[29], inst_cellmath__9[28], inst_cellmath__9[27], inst_cellmath__9[26], inst_cellmath__9[25], inst_cellmath__9[24], inst_cellmath__9[23]}), .inst_cellmath__67_0_in1({inst_cellmath__8[30], inst_cellmath__8[29], inst_cellmath__8[28], inst_cellmath__8[27], inst_cellmath__8[26], inst_cellmath__8[25], inst_cellmath__8[24], inst_cellmath__8[23]}));
cynw_cm_float_div_ieee_inst_cellmath__68_0_bdw410776230_bdw cynw_cm_float_div_ieee_I289 (.inst_cellmath__68_0_out0({inst_cellmath__68[9], inst_cellmath__68[8], inst_cellmath__68[7], inst_cellmath__68[6], inst_cellmath__68[5], inst_cellmath__68[4], inst_cellmath__68[3], inst_cellmath__68[2], inst_cellmath__68[1], inst_cellmath__68[0]}), .inst_cellmath__68_0_in0({inst_cellmath__9[30], inst_cellmath__9[29], inst_cellmath__9[28], inst_cellmath__9[27], inst_cellmath__9[26], inst_cellmath__9[25], inst_cellmath__9[24], inst_cellmath__9[23]}), .inst_cellmath__68_0_in1({inst_cellmath__8[30], inst_cellmath__8[29], inst_cellmath__8[28], inst_cellmath__8[27], inst_cellmath__8[26], inst_cellmath__8[25], inst_cellmath__8[24], inst_cellmath__8[23]}));
cynw_cm_float_div_ieee_inst_cellmath__69__82__bdw410776230_bdw cynw_cm_float_div_ieee_I290 (.inst_cellmath__69__82__out0({N1675}), .inst_cellmath__69__82__in0({inst_cellmath__68[7], inst_cellmath__68[6], inst_cellmath__68[5], inst_cellmath__68[4], inst_cellmath__68[3], inst_cellmath__68[2], inst_cellmath__68[1], inst_cellmath__68[0]}));
cynw_cm_float_div_ieee_inst_cellmath__69__81__bdw410776230_bdw cynw_cm_float_div_ieee_I291 (.inst_cellmath__69__81__out0({N1676}), .inst_cellmath__69__81__in0({N1675}), .inst_cellmath__69__81__in1({inst_cellmath__68[8]}));
cynw_cm_float_div_ieee_inst_cellmath__69_0_bdw410776230_bdw cynw_cm_float_div_ieee_I292 (.inst_cellmath__69_0_out0(inst_cellmath__69), .inst_cellmath__69_0_in0({N1676}), .inst_cellmath__69_0_in1({inst_cellmath__68[9]}));
cynw_cm_float_div_ieee_inst_cellmath__70__83__bdw410776230_bdw cynw_cm_float_div_ieee_I293 (.inst_cellmath__70__83__out0({N1677}), .inst_cellmath__70__83__in0({inst_cellmath__68[8], inst_cellmath__68[7], inst_cellmath__68[6], inst_cellmath__68[5], inst_cellmath__68[4], inst_cellmath__68[3], inst_cellmath__68[2], inst_cellmath__68[1], inst_cellmath__68[0]}));
cynw_cm_float_div_ieee_inst_cellmath__70_0_bdw410776230_bdw cynw_cm_float_div_ieee_I294 (.inst_cellmath__70_0_out0(inst_cellmath__70), .inst_cellmath__70_0_in0({N1677}), .inst_cellmath__70_0_in1({inst_cellmath__68[9]}));
cynw_cm_float_div_ieee_inst_cellmath__71_0_bdw410776230_bdw cynw_cm_float_div_ieee_I295 (.inst_cellmath__71_0_out0(inst_cellmath__71), .inst_cellmath__71_0_in0({inst_cellmath__68[9], inst_cellmath__68[8], inst_cellmath__68[7], inst_cellmath__68[6], inst_cellmath__68[5], inst_cellmath__68[4], inst_cellmath__68[3], inst_cellmath__68[2], inst_cellmath__68[1], inst_cellmath__68[0]}));
cynw_cm_float_div_ieee_inst_cellmath__72_0_bdw410776230_bdw cynw_cm_float_div_ieee_I296 (.inst_cellmath__72_0_out0(inst_cellmath__72), .inst_cellmath__72_0_in0({inst_cellmath__68[8], inst_cellmath__68[7], inst_cellmath__68[6], inst_cellmath__68[5], inst_cellmath__68[4], inst_cellmath__68[3], inst_cellmath__68[2], inst_cellmath__68[1], inst_cellmath__68[0]}));
cynw_cm_float_div_ieee_inst_cellmath__73_0_bdw410776230_bdw cynw_cm_float_div_ieee_I297 (.inst_cellmath__73_0_out0(inst_cellmath__73), .inst_cellmath__73_0_in0(inst_cellmath__71), .inst_cellmath__73_0_in1(inst_cellmath__69));
cynw_cm_float_div_ieee_inst_cellmath__74_0_bdw410776230_bdw cynw_cm_float_div_ieee_I298 (.inst_cellmath__74_0_out0(inst_cellmath__74), .inst_cellmath__74_0_in0(inst_cellmath__72), .inst_cellmath__74_0_in1(inst_cellmath__70));
cynw_cm_float_div_ieee_inst_cellmath__75_0_bdw410776230_bdw cynw_cm_float_div_ieee_I299 (.inst_cellmath__75_0_out0(inst_cellmath__75), .inst_cellmath__75_0_in0({inst_cellmath__8[30], inst_cellmath__8[29], inst_cellmath__8[28], inst_cellmath__8[27], inst_cellmath__8[26], inst_cellmath__8[25], inst_cellmath__8[24], inst_cellmath__8[23]}));
cynw_cm_float_div_ieee_inst_cellmath__76_0_bdw410776230_bdw cynw_cm_float_div_ieee_I300 (.inst_cellmath__76_0_out0(inst_cellmath__76), .inst_cellmath__76_0_in0({inst_cellmath__9[30], inst_cellmath__9[29], inst_cellmath__9[28], inst_cellmath__9[27], inst_cellmath__9[26], inst_cellmath__9[25], inst_cellmath__9[24], inst_cellmath__9[23]}));
cynw_cm_float_div_ieee_inst_cellmath__77_0_bdw410776230_bdw cynw_cm_float_div_ieee_I301 (.inst_cellmath__77_0_out0(inst_cellmath__77), .inst_cellmath__77_0_in0({inst_cellmath__8[22], inst_cellmath__8[21], inst_cellmath__8[20], inst_cellmath__8[19], inst_cellmath__8[18], inst_cellmath__8[17], inst_cellmath__8[16], inst_cellmath__8[15], inst_cellmath__8[14], inst_cellmath__8[13], inst_cellmath__8[12], inst_cellmath__8[11], inst_cellmath__8[10], inst_cellmath__8[9], inst_cellmath__8[8], inst_cellmath__8[7], inst_cellmath__8[6], inst_cellmath__8[5], inst_cellmath__8[4], inst_cellmath__8[3], inst_cellmath__8[2], inst_cellmath__8[1], inst_cellmath__8[0]}));
cynw_cm_float_div_ieee_inst_cellmath__78_0_bdw410776230_bdw cynw_cm_float_div_ieee_I302 (.inst_cellmath__78_0_out0(inst_cellmath__78), .inst_cellmath__78_0_in0({inst_it2_lookup1_cellmath__53[1], inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}));
cynw_cm_float_div_ieee_inst_cellmath__79_1_bdw410776230_bdw cynw_cm_float_div_ieee_I303 (.inst_cellmath__79_1_out0(inst_cellmath__79), .inst_cellmath__79_1_in0(inst_cellmath__77), .inst_cellmath__79_1_in1(inst_cellmath__75));
cynw_cm_float_div_ieee_inst_cellmath__80_0_bdw410776230_bdw cynw_cm_float_div_ieee_I304 (.inst_cellmath__80_0_out0(inst_cellmath__80), .inst_cellmath__80_0_in0(inst_cellmath__78), .inst_cellmath__80_0_in1(inst_cellmath__76));
cynw_cm_float_div_ieee_inst_cellmath__83_0_bdw410776230_bdw cynw_cm_float_div_ieee_I305 (.inst_cellmath__83_0_out0(inst_cellmath__83), .inst_cellmath__83_0_in0(inst_cellmath__77), .inst_cellmath__83_0_in1(inst_cellmath__75));
cynw_cm_float_div_ieee_inst_cellmath__84_0_bdw410776230_bdw cynw_cm_float_div_ieee_I306 (.inst_cellmath__84_0_out0(inst_cellmath__84), .inst_cellmath__84_0_in0(inst_cellmath__78), .inst_cellmath__84_0_in1(inst_cellmath__76));
cynw_cm_float_div_ieee_inst_cellmath__85__85__bdw410776230_bdw cynw_cm_float_div_ieee_I307 (.inst_cellmath__85__85__out0(inst_cellmath__85), .inst_cellmath__85__85__in0({inst_cellmath__8[30], inst_cellmath__8[29], inst_cellmath__8[28], inst_cellmath__8[27], inst_cellmath__8[26], inst_cellmath__8[25], inst_cellmath__8[24], inst_cellmath__8[23]}));
cynw_cm_float_div_ieee_inst_cellmath__86__86__bdw410776230_bdw cynw_cm_float_div_ieee_I308 (.inst_cellmath__86__86__out0(inst_cellmath__86), .inst_cellmath__86__86__in0({inst_cellmath__9[30], inst_cellmath__9[29], inst_cellmath__9[28], inst_cellmath__9[27], inst_cellmath__9[26], inst_cellmath__9[25], inst_cellmath__9[24], inst_cellmath__9[23]}));
cynw_cm_float_div_ieee_inst_cellmath__87__87__bdw410776230_bdw cynw_cm_float_div_ieee_I309 (.inst_cellmath__87__87__out0({N1678}), .inst_cellmath__87__87__in0(inst_cellmath__84), .inst_cellmath__87__87__in1(inst_cellmath__83));
cynw_cm_float_div_ieee_inst_cellmath__87__88__bdw410776230_bdw cynw_cm_float_div_ieee_I310 (.inst_cellmath__87__88__out0({N1679}), .inst_cellmath__87__88__in0(inst_cellmath__86), .inst_cellmath__87__88__in1(inst_cellmath__85));
cynw_cm_float_div_ieee_inst_cellmath__87_0_bdw410776230_bdw cynw_cm_float_div_ieee_I311 (.inst_cellmath__87_0_out0(inst_cellmath__87), .inst_cellmath__87_0_in0({N1679}), .inst_cellmath__87_0_in1({N1678}), .inst_cellmath__87_0_in2(inst_cellmath__80), .inst_cellmath__87_0_in3(inst_cellmath__79));
cynw_cm_float_div_ieee_inst_cellmath__88_0_bdw410776230_bdw cynw_cm_float_div_ieee_I312 (.inst_cellmath__88_0_out0(inst_cellmath__88), .inst_cellmath__88_0_in0(inst_cellmath__86), .inst_cellmath__88_0_in1(inst_cellmath__83));
cynw_cm_float_div_ieee_inst_cellmath__89_0_bdw410776230_bdw cynw_cm_float_div_ieee_I313 (.inst_cellmath__89_0_out0(inst_cellmath__89), .inst_cellmath__89_0_in0(inst_cellmath__85), .inst_cellmath__89_0_in1(inst_cellmath__84));
cynw_cm_float_div_ieee_inst_cellmath__91_0_bdw410776230_bdw cynw_cm_float_div_ieee_I314 (.inst_cellmath__91_0_out0(inst_cellmath__91), .inst_cellmath__91_0_in0({inst_cellmath__9[31]}), .inst_cellmath__91_0_in1({inst_cellmath__8[31]}));
cynw_cm_float_div_ieee_inst_cellmath__92__95__bdw410776230_bdw cynw_cm_float_div_ieee_I315 (.inst_cellmath__92__95__out0({N1680}), .inst_cellmath__92__95__in0(inst_cellmath__91), .inst_cellmath__92__95__in1(inst_cellmath__87));
cynw_cm_float_div_ieee_inst_cellmath__90_2WWMM_bdw410776230_bdw cynw_cm_float_div_ieee_I316 (.inst_cellmath__90_2WWMM_out0({N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750}), .inst_cellmath__90_2WWMM_in0({inst_cellmath__9[31]}), .inst_cellmath__90_2WWMM_in1({inst_it2_lookup1_cellmath__53[0], inst_cellmath__9[20], inst_cellmath__9[19], inst_cellmath__9[18], inst_cellmath__9[17], inst_cellmath__9[16], inst_cellmath__9[15], inst_cellmath__9[14], inst_cellmath__9[13], inst_cellmath__9[12], inst_cellmath__9[11], inst_cellmath__9[10], inst_cellmath__9[9], inst_cellmath__9[8], inst_cellmath__9[7], inst_cellmath__9[6], inst_cellmath__9[5], inst_cellmath__9[4], inst_cellmath__9[3], inst_cellmath__9[2], inst_cellmath__9[1], inst_cellmath__9[0]}), .inst_cellmath__90_2WWMM_in2({N1680}), .inst_cellmath__90_2WWMM_in3({inst_cellmath__8[31]}), .inst_cellmath__90_2WWMM_in4({inst_cellmath__8[21], inst_cellmath__8[20], inst_cellmath__8[19], inst_cellmath__8[18], inst_cellmath__8[17], inst_cellmath__8[16], inst_cellmath__8[15], inst_cellmath__8[14], inst_cellmath__8[13], inst_cellmath__8[12], inst_cellmath__8[11], inst_cellmath__8[10], inst_cellmath__8[9], inst_cellmath__8[8], inst_cellmath__8[7], inst_cellmath__8[6], inst_cellmath__8[5], inst_cellmath__8[4], inst_cellmath__8[3], inst_cellmath__8[2], inst_cellmath__8[1], inst_cellmath__8[0]}), .inst_cellmath__90_2WWMM_in5(inst_cellmath__80), .inst_cellmath__90_2WWMM_in6(inst_cellmath__79));
cynw_cm_float_div_ieee_inst_cellmath__96_0_bdw410776230_bdw cynw_cm_float_div_ieee_I317 (.inst_cellmath__96_0_out0(inst_cellmath__96), .inst_cellmath__96_0_in0({inst_cellmath__12[3], inst_cellmath__12[2], inst_cellmath__12[1], inst_cellmath__12[0]}));
DFFQXL inst_cellmath__98_0_I318 (.Q(inst_cellmath__113[31]), .D(N1750), .CK(clk));
DFFQXL inst_cellmath__100_0_I319 (.Q(inst_cellmath__100), .D(inst_cellmath__87), .CK(clk));
DFFQXL inst_cellmath__101_0_I320 (.Q(inst_cellmath__101), .D(inst_cellmath__88), .CK(clk));
DFFQXL inst_cellmath__102_0_I321 (.Q(inst_cellmath__102), .D(inst_cellmath__89), .CK(clk));
DFFQXL inst_cellmath__103_0_I322 (.Q(inst_cellmath__103), .D(inst_cellmath__69), .CK(clk));
DFFQXL inst_cellmath__104_0_I323 (.Q(inst_cellmath__104), .D(inst_cellmath__73), .CK(clk));
DFFQXL inst_cellmath__105_0_I324 (.Q(inst_cellmath__105), .D(inst_cellmath__70), .CK(clk));
DFFQXL inst_cellmath__106_0_I325 (.Q(inst_cellmath__106), .D(inst_cellmath__74), .CK(clk));
DFFQXL inst_cellmath__110_0_0__I326 (.Q(inst_cellmath__110[0]), .D(inst_cellmath__67[0]), .CK(clk));
DFFQXL inst_cellmath__110_0_1__I327 (.Q(inst_cellmath__110[1]), .D(inst_cellmath__67[1]), .CK(clk));
DFFQXL inst_cellmath__110_0_2__I328 (.Q(inst_cellmath__110[2]), .D(inst_cellmath__67[2]), .CK(clk));
DFFQXL inst_cellmath__110_0_3__I329 (.Q(inst_cellmath__110[3]), .D(inst_cellmath__67[3]), .CK(clk));
DFFQXL inst_cellmath__110_0_4__I330 (.Q(inst_cellmath__110[4]), .D(inst_cellmath__67[4]), .CK(clk));
DFFQXL inst_cellmath__110_0_5__I331 (.Q(inst_cellmath__110[5]), .D(inst_cellmath__67[5]), .CK(clk));
DFFQXL inst_cellmath__110_0_6__I332 (.Q(inst_cellmath__110[6]), .D(inst_cellmath__67[6]), .CK(clk));
DFFQXL inst_cellmath__110_0_7__I333 (.Q(inst_cellmath__110[7]), .D(inst_cellmath__67[7]), .CK(clk));
DFFQXL inst_cellmath__111_0_0__I334 (.Q(inst_cellmath__111[0]), .D(inst_cellmath__68[0]), .CK(clk));
DFFQXL inst_cellmath__111_0_1__I335 (.Q(inst_cellmath__111[1]), .D(inst_cellmath__68[1]), .CK(clk));
DFFQXL inst_cellmath__111_0_2__I336 (.Q(inst_cellmath__111[2]), .D(inst_cellmath__68[2]), .CK(clk));
DFFQXL inst_cellmath__111_0_3__I337 (.Q(inst_cellmath__111[3]), .D(inst_cellmath__68[3]), .CK(clk));
DFFQXL inst_cellmath__111_0_4__I338 (.Q(inst_cellmath__111[4]), .D(inst_cellmath__68[4]), .CK(clk));
DFFQXL inst_cellmath__111_0_5__I339 (.Q(inst_cellmath__111[5]), .D(inst_cellmath__68[5]), .CK(clk));
DFFQXL inst_cellmath__111_0_6__I340 (.Q(inst_cellmath__111[6]), .D(inst_cellmath__68[6]), .CK(clk));
DFFQXL inst_cellmath__111_0_7__I341 (.Q(inst_cellmath__111[7]), .D(inst_cellmath__68[7]), .CK(clk));
DFFQXL inst_cellmath__109_0_I342 (.Q(inst_cellmath__109), .D(inst_cellmath__96), .CK(clk));
INVXL cynw_cm_float_div_ieee_I362 (.Y(N4587), .A(inst_cellmath__109));
INVX2 cynw_cm_float_div_ieee_I369 (.Y(N4594), .A(N4587));
cynw_cm_float_div_ieee_inst_cellmath__133__109__bdw410776230_bdw cynw_cm_float_div_ieee_I343 (.inst_cellmath__133__109__out0({N1685}), .inst_cellmath__133__109__in0(inst_cellmath__103), .inst_cellmath__133__109__in1(inst_cellmath__101), .inst_cellmath__133__109__in2(inst_cellmath__100));
cynw_cm_float_div_ieee_inst_cellmath__135_0_bdw410776230_bdw cynw_cm_float_div_ieee_I344 (.inst_cellmath__135_0_out0(inst_cellmath__135), .inst_cellmath__135_0_in0(inst_cellmath__105), .inst_cellmath__135_0_in1(inst_cellmath__103), .inst_cellmath__135_0_in2(inst_cellmath__102), .inst_cellmath__135_0_in3(inst_cellmath__101), .inst_cellmath__135_0_in4(inst_cellmath__100));
cynw_cm_float_div_ieee_inst_cellmath__136_0_bdw410776230_bdw cynw_cm_float_div_ieee_I345 (.inst_cellmath__136_0_out0(inst_cellmath__136), .inst_cellmath__136_0_in0(inst_cellmath__106), .inst_cellmath__136_0_in1(inst_cellmath__104), .inst_cellmath__136_0_in2(inst_cellmath__102), .inst_cellmath__136_0_in3(inst_cellmath__101), .inst_cellmath__136_0_in4(inst_cellmath__100));
cynw_cm_float_div_ieee_inst_cellmath__137_2_bdw410776230_bdw cynw_cm_float_div_ieee_I346 (.inst_cellmath__137_2_out0(inst_cellmath__137), .inst_cellmath__137_2_in0(inst_cellmath__136), .inst_cellmath__137_2_in1(inst_cellmath__135), .inst_cellmath__137_2_in2(inst_cellmath__122));
cynw_cm_float_div_ieee_inst_cellmath__113__113__bdw410776230_bdw cynw_cm_float_div_ieee_I347 (.inst_cellmath__113__113__out0({inst_cellmath__113[30], inst_cellmath__113[29], inst_cellmath__113[28], inst_cellmath__113[27], inst_cellmath__113[26], inst_cellmath__113[25], inst_cellmath__113[24], inst_cellmath__113[23]}), .inst_cellmath__113__113__in0(inst_cellmath__137), .inst_cellmath__113__113__in1({N1685}), .inst_cellmath__113__113__in2(inst_cellmath__122), .inst_cellmath__113__113__in3({inst_cellmath__111[7], inst_cellmath__111[6], inst_cellmath__111[5], inst_cellmath__111[4], inst_cellmath__111[3], inst_cellmath__111[2], inst_cellmath__111[1], inst_cellmath__111[0]}), .inst_cellmath__113__113__in4({inst_cellmath__110[7], inst_cellmath__110[6], inst_cellmath__110[5], inst_cellmath__110[4], inst_cellmath__110[3], inst_cellmath__110[2], inst_cellmath__110[1], inst_cellmath__110[0]}));
cynw_cm_float_div_ieee_inst_cellmath__113__115__U_2WWMM_bdw410776230_bdw cynw_cm_float_div_ieee_I348 (.inst_cellmath__113__115__U_2WWMM_out0({inst_cellmath__113[22], inst_cellmath__113[21], inst_cellmath__113[20], inst_cellmath__113[19], inst_cellmath__113[18], inst_cellmath__113[17], inst_cellmath__113[16], inst_cellmath__113[15], inst_cellmath__113[14], inst_cellmath__113[13], inst_cellmath__113[12], inst_cellmath__113[11], inst_cellmath__113[10], inst_cellmath__113[9], inst_cellmath__113[8], inst_cellmath__113[7], inst_cellmath__113[6], inst_cellmath__113[5], inst_cellmath__113[4], inst_cellmath__113[3], inst_cellmath__113[2], inst_cellmath__113[1], inst_cellmath__113[0]}), .inst_cellmath__113__115__U_2WWMM_in0(inst_cellmath__137), .inst_cellmath__113__115__U_2WWMM_in1({inst_cellmath__129[22], inst_cellmath__129[21], inst_cellmath__129[20], inst_cellmath__129[19], inst_cellmath__129[18], inst_cellmath__129[17], inst_cellmath__129[16], inst_cellmath__129[15], inst_cellmath__129[14], inst_cellmath__129[13], inst_cellmath__129[12], inst_cellmath__129[11], inst_cellmath__129[10], inst_cellmath__129[9], inst_cellmath__129[8], inst_cellmath__129[7], inst_cellmath__129[6], inst_cellmath__129[5], inst_cellmath__129[4], inst_cellmath__129[3], inst_cellmath__129[2], inst_cellmath__129[1]}), .inst_cellmath__113__115__U_2WWMM_in2({N1922}), .inst_cellmath__113__115__U_2WWMM_in3({inst_cellmath__112[21], inst_cellmath__112[20], inst_cellmath__112[19], inst_cellmath__112[18], inst_cellmath__112[17], inst_cellmath__112[16], inst_cellmath__112[15], inst_cellmath__112[14], inst_cellmath__112[13], inst_cellmath__112[12], inst_cellmath__112[11], inst_cellmath__112[10], inst_cellmath__112[9], inst_cellmath__112[8], inst_cellmath__112[7], inst_cellmath__112[6], inst_cellmath__112[5], inst_cellmath__112[4], inst_cellmath__112[3], inst_cellmath__112[2], inst_cellmath__112[1], inst_cellmath__112[0]}), .inst_cellmath__113__115__U_2WWMM_in4(inst_cellmath__100));
assign inst_cellmath__9[21] = inst_it2_lookup1_cellmath__53[0];
assign inst_cellmath__9[22] = inst_it2_lookup1_cellmath__53[1];
assign inst_cellmath__14[0] = 1'B0;
assign inst_cellmath__16[0] = 1'B0;
assign inst_lookup0_cellmath__27[0] = inst_it2_lookup1_cellmath__53[0];
assign inst_lookup0_cellmath__27[1] = inst_it2_lookup1_cellmath__53[1];
assign inst_cellmath__34[0] = inst_cellmath__35[0];
assign inst_cellmath__34[1] = 1'B0;
assign inst_cellmath__35[1] = 1'B0;
assign inst_cellmath__38__W0[25] = 1'B0;
assign inst_cellmath__39__W0[0] = inst_it2_cellmath__60[3];
assign inst_cellmath__39__W0[1] = inst_it2_cellmath__60[4];
assign inst_cellmath__39__W0[2] = inst_it2_cellmath__60[5];
assign inst_cellmath__39__W0[3] = inst_it2_cellmath__60[6];
assign inst_cellmath__39__W0[4] = inst_it2_cellmath__60[7];
assign inst_cellmath__39__W0[5] = inst_it2_cellmath__60[8];
assign inst_cellmath__39__W0[6] = inst_it2_cellmath__60[9];
assign inst_cellmath__39__W0[7] = inst_it2_cellmath__60[10];
assign inst_cellmath__39__W0[8] = inst_it2_cellmath__60[11];
assign inst_cellmath__39__W0[9] = inst_it2_cellmath__60[12];
assign inst_cellmath__39__W0[10] = inst_it2_cellmath__60[13];
assign inst_cellmath__39__W0[11] = inst_it2_cellmath__60[14];
assign inst_cellmath__39__W0[12] = inst_it2_cellmath__60[15];
assign inst_cellmath__39__W0[13] = inst_it2_cellmath__60[16];
assign inst_cellmath__39__W0[14] = inst_it2_cellmath__60[17];
assign inst_cellmath__39__W0[15] = inst_it2_cellmath__60[18];
assign inst_cellmath__39__W0[16] = inst_it2_cellmath__60[19];
assign inst_cellmath__39__W0[17] = inst_it2_cellmath__60[20];
assign inst_cellmath__39__W0[18] = inst_it2_cellmath__60[21];
assign inst_cellmath__39__W0[19] = inst_it2_cellmath__60[22];
assign inst_cellmath__39__W0[20] = inst_it2_cellmath__60[23];
assign inst_cellmath__39__W0[21] = inst_it2_cellmath__60[24];
assign inst_cellmath__39__W0[22] = inst_it2_cellmath__60[25];
assign inst_cellmath__39__W0[25] = 1'B0;
assign inst_cellmath__39__W1[0] = inst_it2_cellmath__61[2];
assign inst_cellmath__39__W1[1] = inst_it2_cellmath__61[3];
assign inst_cellmath__39__W1[2] = inst_it2_cellmath__61[4];
assign inst_cellmath__39__W1[3] = inst_it2_cellmath__61[5];
assign inst_cellmath__39__W1[4] = inst_it2_cellmath__61[6];
assign inst_cellmath__39__W1[5] = inst_it2_cellmath__61[7];
assign inst_cellmath__39__W1[6] = inst_it2_cellmath__61[8];
assign inst_cellmath__39__W1[7] = inst_it2_cellmath__61[9];
assign inst_cellmath__39__W1[8] = inst_it2_cellmath__61[10];
assign inst_cellmath__39__W1[9] = inst_it2_cellmath__61[11];
assign inst_cellmath__39__W1[10] = inst_it2_cellmath__61[12];
assign inst_cellmath__39__W1[11] = inst_it2_cellmath__61[13];
assign inst_cellmath__39__W1[12] = inst_it2_cellmath__61[14];
assign inst_cellmath__39__W1[13] = inst_it2_cellmath__61[15];
assign inst_cellmath__39__W1[14] = inst_it2_cellmath__61[16];
assign inst_cellmath__39__W1[15] = inst_it2_cellmath__61[17];
assign inst_cellmath__39__W1[16] = inst_it2_cellmath__61[18];
assign inst_cellmath__39__W1[17] = inst_it2_cellmath__61[19];
assign inst_cellmath__39__W1[18] = inst_it2_cellmath__61[20];
assign inst_cellmath__39__W1[19] = inst_it2_cellmath__61[21];
assign inst_cellmath__39__W1[20] = inst_it2_cellmath__61[22];
assign inst_cellmath__39__W1[21] = inst_it2_cellmath__61[23];
assign inst_cellmath__39__W1[22] = inst_it2_cellmath__61[24];
assign inst_cellmath__39__W1[23] = inst_it2_cellmath__61[25];
assign inst_cellmath__42[27] = 1'B0;
assign inst_cellmath__42[28] = 1'B0;
assign inst_cellmath__43[27] = 1'B0;
assign inst_cellmath__43[28] = 1'B0;
assign inst_cellmath__46[25] = 1'B0;
assign inst_cellmath__46[26] = 1'B0;
assign inst_cellmath__46[27] = 1'B0;
assign inst_cellmath__46[28] = 1'B0;
assign inst_cellmath__47[25] = 1'B0;
assign inst_cellmath__47[26] = 1'B0;
assign inst_cellmath__47[27] = 1'B0;
assign inst_cellmath__47[28] = 1'B0;
assign inst_it2_cellmath__60[0] = inst_it2_cellmath__61[0];
assign inst_it2_cellmath__60[1] = 1'B0;
assign inst_it2_cellmath__60[2] = 1'B0;
assign inst_it2_cellmath__61[1] = 1'B0;
assign inst_it2_cellmath__62__W0[25] = 1'B0;
assign inst_cellmath__67[8] = 1'B0;
assign inst_cellmath__67[9] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__23_0_bdw410776230_bdw (
	inst_cellmath__23_0_out0,
	inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__23_0_out0;
input [25:21] inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1;
wire N62,N66,N68,N70,N72;
ADDHX1 inst_cellmath__23_0_I20 (.CO(N62), .S(inst_cellmath__23_0_out0[0]), .A(inst_cellmath__23_0_in0[21]), .B(inst_cellmath__23_0_in1[21]));
ADDFX1 inst_cellmath__23_0_I21 (.CO(N66), .S(inst_cellmath__23_0_out0[1]), .A(inst_cellmath__23_0_in1[22]), .B(inst_cellmath__23_0_in0[22]), .CI(N62));
ADDFX1 inst_cellmath__23_0_I22 (.CO(N68), .S(inst_cellmath__23_0_out0[2]), .A(inst_cellmath__23_0_in1[23]), .B(inst_cellmath__23_0_in0[23]), .CI(N66));
ADDFX1 inst_cellmath__23_0_I23 (.CO(N70), .S(inst_cellmath__23_0_out0[3]), .A(inst_cellmath__23_0_in1[24]), .B(inst_cellmath__23_0_in0[24]), .CI(N68));
ADDFX1 inst_cellmath__23_0_I24 (.CO(N72), .S(inst_cellmath__23_0_out0[4]), .A(inst_cellmath__23_0_in1[25]), .B(inst_cellmath__23_0_in0[25]), .CI(N70));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__22_0_bdw410776230_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__22_0_out0;
input [22:20] inst_cellmath__22_0_in0;
input [2:0] inst_cellmath__22_0_in1;
wire N58,N59,N60,N61,N62,N65,N78 
	,N81;
NAND2XL inst_cellmath__22_0_I19 (.Y(N58), .A(inst_cellmath__22_0_in0[20]), .B(inst_cellmath__22_0_in1[0]));
NOR2XL inst_cellmath__22_0_I20 (.Y(N59), .A(inst_cellmath__22_0_in0[21]), .B(inst_cellmath__22_0_in1[1]));
NAND2XL inst_cellmath__22_0_I21 (.Y(N60), .A(inst_cellmath__22_0_in0[21]), .B(inst_cellmath__22_0_in1[1]));
NOR2XL inst_cellmath__22_0_I22 (.Y(N61), .A(inst_cellmath__22_0_in0[22]), .B(inst_cellmath__22_0_in1[2]));
NAND2XL inst_cellmath__22_0_I23 (.Y(N62), .A(inst_cellmath__22_0_in0[22]), .B(inst_cellmath__22_0_in1[2]));
AO21XL inst_cellmath__22_0_I26 (.Y(N65), .A0(N60), .A1(N58), .B0(N59));
AO21XL inst_cellmath__22_0_I32 (.Y(inst_cellmath__22_0_out0[4]), .A0(N62), .A1(N65), .B0(N61));
NAND2BXL inst_cellmath__22_0_I39 (.Y(N78), .AN(N59), .B(N60));
NAND2BXL inst_cellmath__22_0_I42 (.Y(N81), .AN(N61), .B(N62));
XOR2XL inst_cellmath__22_0_I43 (.Y(inst_cellmath__22_0_out0[0]), .A(inst_cellmath__22_0_in0[20]), .B(inst_cellmath__22_0_in1[0]));
XOR2XL inst_cellmath__22_0_I50 (.Y(inst_cellmath__22_0_out0[1]), .A(N58), .B(N78));
XOR2XL inst_cellmath__22_0_I51 (.Y(inst_cellmath__22_0_out0[2]), .A(N65), .B(N81));
assign inst_cellmath__22_0_out0[3] = inst_cellmath__22_0_out0[4];
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__24_0_bdw410776230_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1,
	inst_cellmath__24_0_in2
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__24_0_out0;
input [4:0] inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1;
input  inst_cellmath__24_0_in2;
MX2XL inst_cellmath__24_0_I10 (.Y(inst_cellmath__24_0_out0[0]), .A(inst_cellmath__24_0_in0[0]), .B(inst_cellmath__24_0_in1[0]), .S0(inst_cellmath__24_0_in2));
MX2XL inst_cellmath__24_0_I11 (.Y(inst_cellmath__24_0_out0[1]), .A(inst_cellmath__24_0_in0[1]), .B(inst_cellmath__24_0_in1[1]), .S0(inst_cellmath__24_0_in2));
MX2XL inst_cellmath__24_0_I12 (.Y(inst_cellmath__24_0_out0[2]), .A(inst_cellmath__24_0_in0[2]), .B(inst_cellmath__24_0_in1[2]), .S0(inst_cellmath__24_0_in2));
MX2XL inst_cellmath__24_0_I13 (.Y(inst_cellmath__24_0_out0[3]), .A(inst_cellmath__24_0_in0[3]), .B(inst_cellmath__24_0_in1[3]), .S0(inst_cellmath__24_0_in2));
MX2XL inst_cellmath__24_0_I14 (.Y(inst_cellmath__24_0_out0[4]), .A(inst_cellmath__24_0_in0[4]), .B(inst_cellmath__24_0_in1[4]), .S0(inst_cellmath__24_0_in2));
endmodule

module cynw_cm_float_div_ieee_inst_lookup0_cellmath__29_0_bdw410776230_bdw (
	inst_lookup0_cellmath__29_0_out0,
	inst_lookup0_cellmath__29_0_in0,
	inst_lookup0_cellmath__29_0_in1
	); /* architecture "gate_level" */ 
output [2:0] inst_lookup0_cellmath__29_0_out0;
input [22:21] inst_lookup0_cellmath__29_0_in0;
input [4:0] inst_lookup0_cellmath__29_0_in1;
wire N41,N116,N183,N212,N248,N252,N253 
	,N259,N263,N287,N379,N393,N457,N514,N519 
	,N525,N527,N530,N532,N533,N536,N798,N895 
	,N933,N934,N938,N939,N1005,N1007,N1038,N1046 
	,N1047,N1051,N1052,N1056,N1057,N1061,N1084,N1089 
	,N1093,N1096,N1099,N1119,N1126,N1133;
INVXL inst_lookup0_cellmath__29_0_I848 (.Y(N1084), .A(inst_lookup0_cellmath__29_0_in0[22]));
INVXL inst_lookup0_cellmath__29_0_I20 (.Y(N41), .A(inst_lookup0_cellmath__29_0_in0[21]));
INVXL inst_lookup0_cellmath__29_0_I853 (.Y(N1089), .A(inst_lookup0_cellmath__29_0_in1[0]));
INVXL inst_lookup0_cellmath__29_0_I857 (.Y(N1093), .A(inst_lookup0_cellmath__29_0_in1[1]));
NOR2XL inst_lookup0_cellmath__29_0_I81 (.Y(N116), .A(N1093), .B(N1089));
NOR2XL inst_lookup0_cellmath__29_0_I133 (.Y(N183), .A(N1089), .B(N1084));
NAND2XL inst_lookup0_cellmath__29_0_I157 (.Y(N212), .A(N41), .B(N1084));
AOI22XL inst_lookup0_cellmath__29_0_I185 (.Y(N248), .A0(N1089), .A1(inst_lookup0_cellmath__29_0_in0[22]), .B0(N212), .B1(inst_lookup0_cellmath__29_0_in1[0]));
AOI22XL inst_lookup0_cellmath__29_0_I189 (.Y(N252), .A0(N1093), .A1(N248), .B0(N183), .B1(inst_lookup0_cellmath__29_0_in1[1]));
NAND2XL hyperpropagate_3_1_A_I899 (.Y(N1119), .A(inst_lookup0_cellmath__29_0_in0[22]), .B(inst_lookup0_cellmath__29_0_in1[0]));
NOR2XL hyperpropagate_3_1_A_I900 (.Y(N253), .A(N1093), .B(N1119));
INVXL inst_lookup0_cellmath__29_0_I860 (.Y(N1096), .A(inst_lookup0_cellmath__29_0_in1[2]));
AOI22XL inst_lookup0_cellmath__29_0_I193 (.Y(N259), .A0(N1096), .A1(N252), .B0(N116), .B1(inst_lookup0_cellmath__29_0_in1[2]));
NAND2XL inst_lookup0_cellmath__29_0_I195 (.Y(N263), .A(N116), .B(inst_lookup0_cellmath__29_0_in1[2]));
NOR2XL inst_lookup0_cellmath__29_0_I217 (.Y(N287), .A(N41), .B(N1084));
NOR2XL inst_lookup0_cellmath__29_0_I295 (.Y(N379), .A(inst_lookup0_cellmath__29_0_in0[21]), .B(inst_lookup0_cellmath__29_0_in0[22]));
NAND2XL hyperpropagate_3_1_A_I901 (.Y(N1126), .A(N1089), .B(N379));
NOR2XL hyperpropagate_3_1_A_I902 (.Y(N393), .A(inst_lookup0_cellmath__29_0_in1[1]), .B(N1126));
AOI22XL inst_lookup0_cellmath__29_0_I355 (.Y(N457), .A0(N1089), .A1(N1084), .B0(N379), .B1(inst_lookup0_cellmath__29_0_in1[0]));
NAND2XL inst_lookup0_cellmath__29_0_I403 (.Y(N514), .A(inst_lookup0_cellmath__29_0_in0[22]), .B(inst_lookup0_cellmath__29_0_in0[21]));
AOI22XL inst_lookup0_cellmath__29_0_I407 (.Y(N519), .A0(N1089), .A1(N514), .B0(N1084), .B1(inst_lookup0_cellmath__29_0_in1[0]));
AOI22XL inst_lookup0_cellmath__29_0_I411 (.Y(N525), .A0(N1093), .A1(N519), .B0(N457), .B1(inst_lookup0_cellmath__29_0_in1[1]));
NAND4BXL inst_lookup0_cellmath__29_0_I885 (.Y(N527), .AN(N1093), .B(inst_lookup0_cellmath__29_0_in1[0]), .C(inst_lookup0_cellmath__29_0_in1[2]), .D(N287));
AOI22XL inst_lookup0_cellmath__29_0_I415 (.Y(N530), .A0(N1096), .A1(N525), .B0(N393), .B1(inst_lookup0_cellmath__29_0_in1[2]));
INVXL inst_lookup0_cellmath__29_0_I863 (.Y(N1099), .A(inst_lookup0_cellmath__29_0_in1[3]));
AOI22XL inst_lookup0_cellmath__29_0_I417 (.Y(N532), .A0(N1099), .A1(N527), .B0(N259), .B1(inst_lookup0_cellmath__29_0_in1[3]));
NOR2XL andori2bb1_A_I903 (.Y(N1133), .A(inst_lookup0_cellmath__29_0_in1[2]), .B(N253));
NOR2XL andori2bb1_A_I904 (.Y(N533), .A(N1133), .B(N1099));
AOI22XL inst_lookup0_cellmath__29_0_I419 (.Y(N536), .A0(N1099), .A1(N530), .B0(N263), .B1(inst_lookup0_cellmath__29_0_in1[3]));
NAND4BXL inst_lookup0_cellmath__29_0_I888 (.Y(N798), .AN(inst_lookup0_cellmath__29_0_in1[1]), .B(N287), .C(N1096), .D(N1089));
AOI22XL inst_lookup0_cellmath__29_0_I713 (.Y(N895), .A0(N41), .A1(N1084), .B0(inst_lookup0_cellmath__29_0_in0[22]), .B1(inst_lookup0_cellmath__29_0_in0[21]));
AOI22XL inst_lookup0_cellmath__29_0_I741 (.Y(N933), .A0(N1089), .A1(N1084), .B0(N895), .B1(inst_lookup0_cellmath__29_0_in1[0]));
AOI22XL inst_lookup0_cellmath__29_0_I742 (.Y(N934), .A0(N1089), .A1(inst_lookup0_cellmath__29_0_in0[22]), .B0(N287), .B1(inst_lookup0_cellmath__29_0_in1[0]));
AOI22XL inst_lookup0_cellmath__29_0_I745 (.Y(N938), .A0(N1093), .A1(N933), .B0(N1084), .B1(inst_lookup0_cellmath__29_0_in1[1]));
NOR2XL inst_lookup0_cellmath__29_0_I746 (.Y(N939), .A(inst_lookup0_cellmath__29_0_in1[1]), .B(N934));
NAND2XL inst_lookup0_cellmath__29_0_I797 (.Y(N1005), .A(N379), .B(inst_lookup0_cellmath__29_0_in1[0]));
NOR2XL inst_lookup0_cellmath__29_0_I798 (.Y(N1007), .A(N1089), .B(N212));
NOR2XL inst_lookup0_cellmath__29_0_I819 (.Y(N1038), .A(N1089), .B(inst_lookup0_cellmath__29_0_in0[22]));
AOI22XL inst_lookup0_cellmath__29_0_I823 (.Y(N1046), .A0(N1093), .A1(N1038), .B0(N1005), .B1(inst_lookup0_cellmath__29_0_in1[1]));
NAND2XL inst_lookup0_cellmath__29_0_I824 (.Y(N1047), .A(N1007), .B(inst_lookup0_cellmath__29_0_in1[1]));
AOI22XL inst_lookup0_cellmath__29_0_I827 (.Y(N1051), .A0(N1096), .A1(N1046), .B0(N938), .B1(inst_lookup0_cellmath__29_0_in1[2]));
AOI22XL inst_lookup0_cellmath__29_0_I828 (.Y(N1052), .A0(N1096), .A1(N1047), .B0(N939), .B1(inst_lookup0_cellmath__29_0_in1[2]));
AOI22XL inst_lookup0_cellmath__29_0_I831 (.Y(N1056), .A0(N1099), .A1(N1051), .B0(N798), .B1(inst_lookup0_cellmath__29_0_in1[3]));
NOR2XL inst_lookup0_cellmath__29_0_I832 (.Y(N1057), .A(inst_lookup0_cellmath__29_0_in1[3]), .B(N1052));
INVXL inst_lookup0_cellmath__29_0_I834 (.Y(N1061), .A(inst_lookup0_cellmath__29_0_in1[4]));
AOI22XL inst_lookup0_cellmath__29_0_I1039 (.Y(inst_lookup0_cellmath__29_0_out0[0]), .A0(inst_lookup0_cellmath__29_0_in1[4]), .A1(N532), .B0(N1061), .B1(N1056));
AOI22XL inst_lookup0_cellmath__29_0_I836 (.Y(inst_lookup0_cellmath__29_0_out0[1]), .A0(N1061), .A1(N1057), .B0(N533), .B1(inst_lookup0_cellmath__29_0_in1[4]));
NOR2XL inst_lookup0_cellmath__29_0_I837 (.Y(inst_lookup0_cellmath__29_0_out0[2]), .A(N1061), .B(N536));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__30__31__bdw410776230_bdw (
	inst_cellmath__30__31__out0,
	inst_cellmath__30__31__in0,
	inst_cellmath__30__31__in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__30__31__out0;
input [0:0] inst_cellmath__30__31__in0;
input [22:0] inst_cellmath__30__31__in1;
wire N351;
INVXL buf1_A_I102 (.Y(N351), .A(inst_cellmath__30__31__in0[0]));
INVXL buf1_A_I103 (.Y(inst_cellmath__30__31__out0[24]), .A(N351));
AND2XL inst_cellmath__30__31__I27 (.Y(inst_cellmath__30__31__out0[1]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[0]));
AND2XL inst_cellmath__30__31__I28 (.Y(inst_cellmath__30__31__out0[2]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[1]));
AND2XL inst_cellmath__30__31__I29 (.Y(inst_cellmath__30__31__out0[3]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[2]));
AND2XL inst_cellmath__30__31__I30 (.Y(inst_cellmath__30__31__out0[4]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[3]));
AND2XL inst_cellmath__30__31__I31 (.Y(inst_cellmath__30__31__out0[5]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[4]));
AND2XL inst_cellmath__30__31__I32 (.Y(inst_cellmath__30__31__out0[6]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[5]));
AND2XL inst_cellmath__30__31__I33 (.Y(inst_cellmath__30__31__out0[7]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[6]));
AND2XL inst_cellmath__30__31__I34 (.Y(inst_cellmath__30__31__out0[8]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[7]));
AND2XL inst_cellmath__30__31__I35 (.Y(inst_cellmath__30__31__out0[9]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[8]));
AND2XL inst_cellmath__30__31__I36 (.Y(inst_cellmath__30__31__out0[10]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[9]));
AND2XL inst_cellmath__30__31__I37 (.Y(inst_cellmath__30__31__out0[11]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[10]));
AND2XL inst_cellmath__30__31__I38 (.Y(inst_cellmath__30__31__out0[12]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[11]));
AND2XL inst_cellmath__30__31__I39 (.Y(inst_cellmath__30__31__out0[13]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[12]));
AND2XL inst_cellmath__30__31__I40 (.Y(inst_cellmath__30__31__out0[14]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[13]));
AND2XL inst_cellmath__30__31__I41 (.Y(inst_cellmath__30__31__out0[15]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[14]));
AND2XL inst_cellmath__30__31__I42 (.Y(inst_cellmath__30__31__out0[16]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[15]));
AND2XL inst_cellmath__30__31__I43 (.Y(inst_cellmath__30__31__out0[17]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[16]));
AND2XL inst_cellmath__30__31__I44 (.Y(inst_cellmath__30__31__out0[18]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[17]));
AND2XL inst_cellmath__30__31__I45 (.Y(inst_cellmath__30__31__out0[19]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[18]));
AND2XL inst_cellmath__30__31__I46 (.Y(inst_cellmath__30__31__out0[20]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[19]));
AND2XL inst_cellmath__30__31__I47 (.Y(inst_cellmath__30__31__out0[21]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[20]));
AND2XL inst_cellmath__30__31__I48 (.Y(inst_cellmath__30__31__out0[22]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[21]));
AND2XL inst_cellmath__30__31__I49 (.Y(inst_cellmath__30__31__out0[23]), .A(inst_cellmath__30__31__out0[24]), .B(inst_cellmath__30__31__in1[22]));
assign inst_cellmath__30__31__out0[0] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__31__35__bdw410776230_bdw (
	inst_cellmath__31__35__out0,
	inst_cellmath__31__35__in0,
	inst_cellmath__31__35__in1
	); /* architecture "gate_level" */ 
output [25:0] inst_cellmath__31__35__out0;
input [1:1] inst_cellmath__31__35__in0;
input [22:0] inst_cellmath__31__35__in1;
wire N356;
INVXL buf1_A_I104 (.Y(N356), .A(inst_cellmath__31__35__in0[1]));
INVXL buf1_A_I105 (.Y(inst_cellmath__31__35__out0[25]), .A(N356));
AND2XL inst_cellmath__31__35__I29 (.Y(inst_cellmath__31__35__out0[2]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[0]));
AND2XL inst_cellmath__31__35__I30 (.Y(inst_cellmath__31__35__out0[3]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[1]));
AND2XL inst_cellmath__31__35__I31 (.Y(inst_cellmath__31__35__out0[4]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[2]));
AND2XL inst_cellmath__31__35__I32 (.Y(inst_cellmath__31__35__out0[5]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[3]));
AND2XL inst_cellmath__31__35__I33 (.Y(inst_cellmath__31__35__out0[6]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[4]));
AND2XL inst_cellmath__31__35__I34 (.Y(inst_cellmath__31__35__out0[7]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[5]));
AND2XL inst_cellmath__31__35__I35 (.Y(inst_cellmath__31__35__out0[8]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[6]));
AND2XL inst_cellmath__31__35__I36 (.Y(inst_cellmath__31__35__out0[9]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[7]));
AND2XL inst_cellmath__31__35__I37 (.Y(inst_cellmath__31__35__out0[10]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[8]));
AND2XL inst_cellmath__31__35__I38 (.Y(inst_cellmath__31__35__out0[11]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[9]));
AND2XL inst_cellmath__31__35__I39 (.Y(inst_cellmath__31__35__out0[12]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[10]));
AND2XL inst_cellmath__31__35__I40 (.Y(inst_cellmath__31__35__out0[13]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[11]));
AND2XL inst_cellmath__31__35__I41 (.Y(inst_cellmath__31__35__out0[14]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[12]));
AND2XL inst_cellmath__31__35__I42 (.Y(inst_cellmath__31__35__out0[15]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[13]));
AND2XL inst_cellmath__31__35__I43 (.Y(inst_cellmath__31__35__out0[16]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[14]));
AND2XL inst_cellmath__31__35__I44 (.Y(inst_cellmath__31__35__out0[17]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[15]));
AND2XL inst_cellmath__31__35__I45 (.Y(inst_cellmath__31__35__out0[18]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[16]));
AND2XL inst_cellmath__31__35__I46 (.Y(inst_cellmath__31__35__out0[19]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[17]));
AND2XL inst_cellmath__31__35__I47 (.Y(inst_cellmath__31__35__out0[20]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[18]));
AND2XL inst_cellmath__31__35__I48 (.Y(inst_cellmath__31__35__out0[21]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[19]));
AND2XL inst_cellmath__31__35__I49 (.Y(inst_cellmath__31__35__out0[22]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[20]));
AND2XL inst_cellmath__31__35__I50 (.Y(inst_cellmath__31__35__out0[23]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[21]));
AND2XL inst_cellmath__31__35__I51 (.Y(inst_cellmath__31__35__out0[24]), .A(inst_cellmath__31__35__out0[25]), .B(inst_cellmath__31__35__in1[22]));
assign inst_cellmath__31__35__out0[0] = 1'B0;
assign inst_cellmath__31__35__out0[1] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__20_0_bdw410776230_bdw (
	inst_cellmath__20_0_out0,
	inst_cellmath__20_0_in0,
	inst_cellmath__20_0_in1,
	inst_cellmath__20_0_in2
	); /* architecture "gate_level" */ 
output [23:0] inst_cellmath__20_0_out0;
input [22:0] inst_cellmath__20_0_in0;
input [23:0] inst_cellmath__20_0_in1;
input  inst_cellmath__20_0_in2;
wire N325,N328;
INVXL buf1_A_I85 (.Y(N328), .A(inst_cellmath__20_0_in2));
INVXL buf1_A_I86 (.Y(N325), .A(N328));
OR2XL inst_cellmath__20_0_I83 (.Y(inst_cellmath__20_0_out0[0]), .A(N325), .B(inst_cellmath__20_0_in1[0]));
MX2XL inst_cellmath__20_0_I49 (.Y(inst_cellmath__20_0_out0[1]), .A(inst_cellmath__20_0_in1[1]), .B(inst_cellmath__20_0_in0[0]), .S0(N325));
MX2XL inst_cellmath__20_0_I50 (.Y(inst_cellmath__20_0_out0[2]), .A(inst_cellmath__20_0_in1[2]), .B(inst_cellmath__20_0_in0[1]), .S0(N325));
MX2XL inst_cellmath__20_0_I51 (.Y(inst_cellmath__20_0_out0[3]), .A(inst_cellmath__20_0_in1[3]), .B(inst_cellmath__20_0_in0[2]), .S0(N325));
MX2XL inst_cellmath__20_0_I52 (.Y(inst_cellmath__20_0_out0[4]), .A(inst_cellmath__20_0_in1[4]), .B(inst_cellmath__20_0_in0[3]), .S0(N325));
MX2XL inst_cellmath__20_0_I53 (.Y(inst_cellmath__20_0_out0[5]), .A(inst_cellmath__20_0_in1[5]), .B(inst_cellmath__20_0_in0[4]), .S0(N325));
MX2XL inst_cellmath__20_0_I54 (.Y(inst_cellmath__20_0_out0[6]), .A(inst_cellmath__20_0_in1[6]), .B(inst_cellmath__20_0_in0[5]), .S0(N325));
MX2XL inst_cellmath__20_0_I55 (.Y(inst_cellmath__20_0_out0[7]), .A(inst_cellmath__20_0_in1[7]), .B(inst_cellmath__20_0_in0[6]), .S0(N325));
MX2XL inst_cellmath__20_0_I56 (.Y(inst_cellmath__20_0_out0[8]), .A(inst_cellmath__20_0_in1[8]), .B(inst_cellmath__20_0_in0[7]), .S0(N325));
MX2XL inst_cellmath__20_0_I57 (.Y(inst_cellmath__20_0_out0[9]), .A(inst_cellmath__20_0_in1[9]), .B(inst_cellmath__20_0_in0[8]), .S0(N325));
MX2XL inst_cellmath__20_0_I58 (.Y(inst_cellmath__20_0_out0[10]), .A(inst_cellmath__20_0_in1[10]), .B(inst_cellmath__20_0_in0[9]), .S0(N325));
MX2XL inst_cellmath__20_0_I59 (.Y(inst_cellmath__20_0_out0[11]), .A(inst_cellmath__20_0_in1[11]), .B(inst_cellmath__20_0_in0[10]), .S0(N325));
MX2XL inst_cellmath__20_0_I60 (.Y(inst_cellmath__20_0_out0[12]), .A(inst_cellmath__20_0_in1[12]), .B(inst_cellmath__20_0_in0[11]), .S0(N325));
MX2XL inst_cellmath__20_0_I61 (.Y(inst_cellmath__20_0_out0[13]), .A(inst_cellmath__20_0_in1[13]), .B(inst_cellmath__20_0_in0[12]), .S0(N325));
MX2XL inst_cellmath__20_0_I62 (.Y(inst_cellmath__20_0_out0[14]), .A(inst_cellmath__20_0_in1[14]), .B(inst_cellmath__20_0_in0[13]), .S0(N325));
MX2XL inst_cellmath__20_0_I63 (.Y(inst_cellmath__20_0_out0[15]), .A(inst_cellmath__20_0_in1[15]), .B(inst_cellmath__20_0_in0[14]), .S0(N325));
MX2XL inst_cellmath__20_0_I64 (.Y(inst_cellmath__20_0_out0[16]), .A(inst_cellmath__20_0_in1[16]), .B(inst_cellmath__20_0_in0[15]), .S0(N325));
MX2XL inst_cellmath__20_0_I65 (.Y(inst_cellmath__20_0_out0[17]), .A(inst_cellmath__20_0_in1[17]), .B(inst_cellmath__20_0_in0[16]), .S0(N325));
MX2XL inst_cellmath__20_0_I66 (.Y(inst_cellmath__20_0_out0[18]), .A(inst_cellmath__20_0_in1[18]), .B(inst_cellmath__20_0_in0[17]), .S0(N325));
MX2XL inst_cellmath__20_0_I67 (.Y(inst_cellmath__20_0_out0[19]), .A(inst_cellmath__20_0_in1[19]), .B(inst_cellmath__20_0_in0[18]), .S0(N325));
MX2XL inst_cellmath__20_0_I68 (.Y(inst_cellmath__20_0_out0[20]), .A(inst_cellmath__20_0_in1[20]), .B(inst_cellmath__20_0_in0[19]), .S0(N325));
MX2XL inst_cellmath__20_0_I69 (.Y(inst_cellmath__20_0_out0[21]), .A(inst_cellmath__20_0_in1[21]), .B(inst_cellmath__20_0_in0[20]), .S0(N325));
MX2XL inst_cellmath__20_0_I70 (.Y(inst_cellmath__20_0_out0[22]), .A(inst_cellmath__20_0_in1[22]), .B(inst_cellmath__20_0_in0[21]), .S0(N325));
MX2XL inst_cellmath__20_0_I71 (.Y(inst_cellmath__20_0_out0[23]), .A(inst_cellmath__20_0_in1[23]), .B(inst_cellmath__20_0_in0[22]), .S0(N325));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__21_0_bdw410776230_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1,
	inst_cellmath__21_0_in2
	); /* architecture "gate_level" */ 
output [23:0] inst_cellmath__21_0_out0;
input [22:0] inst_cellmath__21_0_in0;
input [23:0] inst_cellmath__21_0_in1;
input  inst_cellmath__21_0_in2;
wire N146,N147,N148,N149,N150,N151,N152 
	,N153,N154,N155,N156,N157,N158,N159,N160 
	,N161,N162,N163,N164,N165,N166,N217,N220 
	,N221;
INVXL inst_cellmath__21_0_I48 (.Y(N146), .A(inst_cellmath__21_0_in1[1]));
INVXL inst_cellmath__21_0_I49 (.Y(N147), .A(inst_cellmath__21_0_in1[2]));
INVXL inst_cellmath__21_0_I50 (.Y(N148), .A(inst_cellmath__21_0_in1[3]));
INVXL inst_cellmath__21_0_I51 (.Y(N149), .A(inst_cellmath__21_0_in1[4]));
INVXL inst_cellmath__21_0_I52 (.Y(N150), .A(inst_cellmath__21_0_in1[5]));
INVXL inst_cellmath__21_0_I53 (.Y(N151), .A(inst_cellmath__21_0_in1[6]));
INVXL inst_cellmath__21_0_I54 (.Y(N152), .A(inst_cellmath__21_0_in1[7]));
INVXL inst_cellmath__21_0_I55 (.Y(N153), .A(inst_cellmath__21_0_in1[8]));
INVXL inst_cellmath__21_0_I56 (.Y(N154), .A(inst_cellmath__21_0_in1[9]));
INVXL inst_cellmath__21_0_I57 (.Y(N155), .A(inst_cellmath__21_0_in1[10]));
INVXL inst_cellmath__21_0_I58 (.Y(N156), .A(inst_cellmath__21_0_in1[11]));
INVXL inst_cellmath__21_0_I59 (.Y(N157), .A(inst_cellmath__21_0_in1[12]));
INVXL inst_cellmath__21_0_I60 (.Y(N158), .A(inst_cellmath__21_0_in1[13]));
INVXL inst_cellmath__21_0_I61 (.Y(N159), .A(inst_cellmath__21_0_in1[14]));
INVXL inst_cellmath__21_0_I62 (.Y(N160), .A(inst_cellmath__21_0_in1[15]));
INVXL inst_cellmath__21_0_I63 (.Y(N161), .A(inst_cellmath__21_0_in1[16]));
INVXL inst_cellmath__21_0_I64 (.Y(N162), .A(inst_cellmath__21_0_in1[17]));
INVXL inst_cellmath__21_0_I65 (.Y(N163), .A(inst_cellmath__21_0_in1[18]));
INVXL inst_cellmath__21_0_I66 (.Y(N164), .A(inst_cellmath__21_0_in1[19]));
INVXL inst_cellmath__21_0_I67 (.Y(N165), .A(inst_cellmath__21_0_in1[20]));
INVXL inst_cellmath__21_0_I68 (.Y(N166), .A(inst_cellmath__21_0_in1[21]));
INVXL inst_cellmath__21_0_I107 (.Y(N217), .A(inst_cellmath__21_0_in2));
NAND2BXL inst_cellmath__21_0_I112 (.Y(inst_cellmath__21_0_out0[0]), .AN(inst_cellmath__21_0_in1[0]), .B(N217));
AOI22XL inst_cellmath__21_0_I73 (.Y(inst_cellmath__21_0_out0[1]), .A0(N217), .A1(N146), .B0(inst_cellmath__21_0_in0[0]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I74 (.Y(inst_cellmath__21_0_out0[2]), .A0(N217), .A1(N147), .B0(inst_cellmath__21_0_in0[1]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I75 (.Y(inst_cellmath__21_0_out0[3]), .A0(N217), .A1(N148), .B0(inst_cellmath__21_0_in0[2]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I76 (.Y(inst_cellmath__21_0_out0[4]), .A0(N217), .A1(N149), .B0(inst_cellmath__21_0_in0[3]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I77 (.Y(inst_cellmath__21_0_out0[5]), .A0(N217), .A1(N150), .B0(inst_cellmath__21_0_in0[4]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I78 (.Y(inst_cellmath__21_0_out0[6]), .A0(N217), .A1(N151), .B0(inst_cellmath__21_0_in0[5]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I79 (.Y(inst_cellmath__21_0_out0[7]), .A0(N217), .A1(N152), .B0(inst_cellmath__21_0_in0[6]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I80 (.Y(inst_cellmath__21_0_out0[8]), .A0(N217), .A1(N153), .B0(inst_cellmath__21_0_in0[7]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I81 (.Y(inst_cellmath__21_0_out0[9]), .A0(N217), .A1(N154), .B0(inst_cellmath__21_0_in0[8]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I82 (.Y(inst_cellmath__21_0_out0[10]), .A0(N217), .A1(N155), .B0(inst_cellmath__21_0_in0[9]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I83 (.Y(inst_cellmath__21_0_out0[11]), .A0(N217), .A1(N156), .B0(inst_cellmath__21_0_in0[10]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I84 (.Y(inst_cellmath__21_0_out0[12]), .A0(N217), .A1(N157), .B0(inst_cellmath__21_0_in0[11]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I85 (.Y(inst_cellmath__21_0_out0[13]), .A0(N217), .A1(N158), .B0(inst_cellmath__21_0_in0[12]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I86 (.Y(inst_cellmath__21_0_out0[14]), .A0(N217), .A1(N159), .B0(inst_cellmath__21_0_in0[13]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I87 (.Y(inst_cellmath__21_0_out0[15]), .A0(N217), .A1(N160), .B0(inst_cellmath__21_0_in0[14]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I88 (.Y(inst_cellmath__21_0_out0[16]), .A0(N217), .A1(N161), .B0(inst_cellmath__21_0_in0[15]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I89 (.Y(inst_cellmath__21_0_out0[17]), .A0(N217), .A1(N162), .B0(inst_cellmath__21_0_in0[16]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I90 (.Y(inst_cellmath__21_0_out0[18]), .A0(N217), .A1(N163), .B0(inst_cellmath__21_0_in0[17]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I91 (.Y(inst_cellmath__21_0_out0[19]), .A0(N217), .A1(N164), .B0(inst_cellmath__21_0_in0[18]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I92 (.Y(inst_cellmath__21_0_out0[20]), .A0(N217), .A1(N165), .B0(inst_cellmath__21_0_in0[19]), .B1(inst_cellmath__21_0_in2));
AOI22XL inst_cellmath__21_0_I93 (.Y(inst_cellmath__21_0_out0[21]), .A0(N217), .A1(N166), .B0(inst_cellmath__21_0_in0[20]), .B1(inst_cellmath__21_0_in2));
INVXL inst_cellmath__21_0_I110 (.Y(N220), .A(inst_cellmath__21_0_in1[22]));
AOI22XL inst_cellmath__21_0_I94 (.Y(inst_cellmath__21_0_out0[22]), .A0(N217), .A1(N220), .B0(inst_cellmath__21_0_in0[21]), .B1(inst_cellmath__21_0_in2));
INVXL inst_cellmath__21_0_I111 (.Y(N221), .A(inst_cellmath__21_0_in1[23]));
AOI22XL inst_cellmath__21_0_I95 (.Y(inst_cellmath__21_0_out0[23]), .A0(N217), .A1(N221), .B0(inst_cellmath__21_0_in0[22]), .B1(inst_cellmath__21_0_in2));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__30_2mx_bdw410776230_bdw (
	inst_cellmath__30_2mx_out0,
	inst_cellmath__30_2mx_in0,
	inst_cellmath__30_2mx_in1
	); /* architecture "gate_level" */ 
output [25:0] inst_cellmath__30_2mx_out0;
input [2:2] inst_cellmath__30_2mx_in0;
input [24:1] inst_cellmath__30_2mx_in1;
wire N340;
INVXL inst_cellmath__30_2mx_I92 (.Y(inst_cellmath__30_2mx_out0[0]), .A(inst_cellmath__30_2mx_in0[2]));
INVXL inst_cellmath__30_2mx_I87 (.Y(N340), .A(inst_cellmath__30_2mx_out0[0]));
XNOR2X1 inst_cellmath__30_2mx_I29 (.Y(inst_cellmath__30_2mx_out0[1]), .A(inst_cellmath__30_2mx_in1[1]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I30 (.Y(inst_cellmath__30_2mx_out0[2]), .A(inst_cellmath__30_2mx_in1[2]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I31 (.Y(inst_cellmath__30_2mx_out0[3]), .A(inst_cellmath__30_2mx_in1[3]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I32 (.Y(inst_cellmath__30_2mx_out0[4]), .A(inst_cellmath__30_2mx_in1[4]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I33 (.Y(inst_cellmath__30_2mx_out0[5]), .A(inst_cellmath__30_2mx_in1[5]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I34 (.Y(inst_cellmath__30_2mx_out0[6]), .A(inst_cellmath__30_2mx_in1[6]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I35 (.Y(inst_cellmath__30_2mx_out0[7]), .A(inst_cellmath__30_2mx_in1[7]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I36 (.Y(inst_cellmath__30_2mx_out0[8]), .A(inst_cellmath__30_2mx_in1[8]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I37 (.Y(inst_cellmath__30_2mx_out0[9]), .A(inst_cellmath__30_2mx_in1[9]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I38 (.Y(inst_cellmath__30_2mx_out0[10]), .A(inst_cellmath__30_2mx_in1[10]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I39 (.Y(inst_cellmath__30_2mx_out0[11]), .A(inst_cellmath__30_2mx_in1[11]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I40 (.Y(inst_cellmath__30_2mx_out0[12]), .A(inst_cellmath__30_2mx_in1[12]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I41 (.Y(inst_cellmath__30_2mx_out0[13]), .A(inst_cellmath__30_2mx_in1[13]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I42 (.Y(inst_cellmath__30_2mx_out0[14]), .A(inst_cellmath__30_2mx_in1[14]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I43 (.Y(inst_cellmath__30_2mx_out0[15]), .A(inst_cellmath__30_2mx_in1[15]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I44 (.Y(inst_cellmath__30_2mx_out0[16]), .A(inst_cellmath__30_2mx_in1[16]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I45 (.Y(inst_cellmath__30_2mx_out0[17]), .A(inst_cellmath__30_2mx_in1[17]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I46 (.Y(inst_cellmath__30_2mx_out0[18]), .A(inst_cellmath__30_2mx_in1[18]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I47 (.Y(inst_cellmath__30_2mx_out0[19]), .A(inst_cellmath__30_2mx_in1[19]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I48 (.Y(inst_cellmath__30_2mx_out0[20]), .A(inst_cellmath__30_2mx_in1[20]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I49 (.Y(inst_cellmath__30_2mx_out0[21]), .A(inst_cellmath__30_2mx_in1[21]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I50 (.Y(inst_cellmath__30_2mx_out0[22]), .A(inst_cellmath__30_2mx_in1[22]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I51 (.Y(inst_cellmath__30_2mx_out0[23]), .A(inst_cellmath__30_2mx_in1[23]), .B(N340));
XNOR2X1 inst_cellmath__30_2mx_I52 (.Y(inst_cellmath__30_2mx_out0[24]), .A(inst_cellmath__30_2mx_in1[24]), .B(N340));
assign inst_cellmath__30_2mx_out0[25] = inst_cellmath__30_2mx_out0[0];
endmodule

module cynw_cm_float_div_ieee_inst_fa_1033_10_bdw410776230_bdw (
	inst_fa_1033_10_out0,
	inst_fa_1033_10_out1,
	inst_fa_1033_10_in0,
	inst_fa_1033_10_in1,
	inst_fa_1033_10_in2,
	inst_fa_1033_10_in3
	); /* architecture "gate_level" */ 
output [25:0] inst_fa_1033_10_out0;
output [24:0] inst_fa_1033_10_out1;
input  inst_fa_1033_10_in0;
input [25:0] inst_fa_1033_10_in1;
input [23:0] inst_fa_1033_10_in2,
	inst_fa_1033_10_in3;
wire N231;
ADDFX1 inst_fa_1033_10_I2 (.CO(inst_fa_1033_10_out1[2]), .S(inst_fa_1033_10_out0[2]), .A(inst_fa_1033_10_in2[0]), .B(inst_fa_1033_10_in3[0]), .CI(inst_fa_1033_10_in1[2]));
ADDFX1 inst_fa_1033_10_I3 (.CO(inst_fa_1033_10_out1[3]), .S(inst_fa_1033_10_out0[3]), .A(inst_fa_1033_10_in2[1]), .B(inst_fa_1033_10_in3[1]), .CI(inst_fa_1033_10_in1[3]));
ADDFX1 inst_fa_1033_10_I4 (.CO(inst_fa_1033_10_out1[4]), .S(inst_fa_1033_10_out0[4]), .A(inst_fa_1033_10_in2[2]), .B(inst_fa_1033_10_in3[2]), .CI(inst_fa_1033_10_in1[4]));
ADDFX1 inst_fa_1033_10_I5 (.CO(inst_fa_1033_10_out1[5]), .S(inst_fa_1033_10_out0[5]), .A(inst_fa_1033_10_in2[3]), .B(inst_fa_1033_10_in3[3]), .CI(inst_fa_1033_10_in1[5]));
ADDFX1 inst_fa_1033_10_I6 (.CO(inst_fa_1033_10_out1[6]), .S(inst_fa_1033_10_out0[6]), .A(inst_fa_1033_10_in2[4]), .B(inst_fa_1033_10_in3[4]), .CI(inst_fa_1033_10_in1[6]));
ADDFX1 inst_fa_1033_10_I7 (.CO(inst_fa_1033_10_out1[7]), .S(inst_fa_1033_10_out0[7]), .A(inst_fa_1033_10_in2[5]), .B(inst_fa_1033_10_in3[5]), .CI(inst_fa_1033_10_in1[7]));
ADDFX1 inst_fa_1033_10_I8 (.CO(inst_fa_1033_10_out1[8]), .S(inst_fa_1033_10_out0[8]), .A(inst_fa_1033_10_in2[6]), .B(inst_fa_1033_10_in3[6]), .CI(inst_fa_1033_10_in1[8]));
ADDFX1 inst_fa_1033_10_I9 (.CO(inst_fa_1033_10_out1[9]), .S(inst_fa_1033_10_out0[9]), .A(inst_fa_1033_10_in2[7]), .B(inst_fa_1033_10_in3[7]), .CI(inst_fa_1033_10_in1[9]));
ADDFX1 inst_fa_1033_10_I10 (.CO(inst_fa_1033_10_out1[10]), .S(inst_fa_1033_10_out0[10]), .A(inst_fa_1033_10_in2[8]), .B(inst_fa_1033_10_in3[8]), .CI(inst_fa_1033_10_in1[10]));
ADDFX1 inst_fa_1033_10_I11 (.CO(inst_fa_1033_10_out1[11]), .S(inst_fa_1033_10_out0[11]), .A(inst_fa_1033_10_in2[9]), .B(inst_fa_1033_10_in3[9]), .CI(inst_fa_1033_10_in1[11]));
ADDFX1 inst_fa_1033_10_I12 (.CO(inst_fa_1033_10_out1[12]), .S(inst_fa_1033_10_out0[12]), .A(inst_fa_1033_10_in2[10]), .B(inst_fa_1033_10_in3[10]), .CI(inst_fa_1033_10_in1[12]));
ADDFX1 inst_fa_1033_10_I13 (.CO(inst_fa_1033_10_out1[13]), .S(inst_fa_1033_10_out0[13]), .A(inst_fa_1033_10_in2[11]), .B(inst_fa_1033_10_in3[11]), .CI(inst_fa_1033_10_in1[13]));
ADDFX1 inst_fa_1033_10_I14 (.CO(inst_fa_1033_10_out1[14]), .S(inst_fa_1033_10_out0[14]), .A(inst_fa_1033_10_in2[12]), .B(inst_fa_1033_10_in3[12]), .CI(inst_fa_1033_10_in1[14]));
ADDFX1 inst_fa_1033_10_I15 (.CO(inst_fa_1033_10_out1[15]), .S(inst_fa_1033_10_out0[15]), .A(inst_fa_1033_10_in2[13]), .B(inst_fa_1033_10_in3[13]), .CI(inst_fa_1033_10_in1[15]));
ADDFX1 inst_fa_1033_10_I16 (.CO(inst_fa_1033_10_out1[16]), .S(inst_fa_1033_10_out0[16]), .A(inst_fa_1033_10_in2[14]), .B(inst_fa_1033_10_in3[14]), .CI(inst_fa_1033_10_in1[16]));
ADDFX1 inst_fa_1033_10_I17 (.CO(inst_fa_1033_10_out1[17]), .S(inst_fa_1033_10_out0[17]), .A(inst_fa_1033_10_in2[15]), .B(inst_fa_1033_10_in3[15]), .CI(inst_fa_1033_10_in1[17]));
ADDFX1 inst_fa_1033_10_I18 (.CO(inst_fa_1033_10_out1[18]), .S(inst_fa_1033_10_out0[18]), .A(inst_fa_1033_10_in2[16]), .B(inst_fa_1033_10_in3[16]), .CI(inst_fa_1033_10_in1[18]));
ADDFX1 inst_fa_1033_10_I19 (.CO(inst_fa_1033_10_out1[19]), .S(inst_fa_1033_10_out0[19]), .A(inst_fa_1033_10_in2[17]), .B(inst_fa_1033_10_in3[17]), .CI(inst_fa_1033_10_in1[19]));
ADDFX1 inst_fa_1033_10_I20 (.CO(inst_fa_1033_10_out1[20]), .S(inst_fa_1033_10_out0[20]), .A(inst_fa_1033_10_in2[18]), .B(inst_fa_1033_10_in3[18]), .CI(inst_fa_1033_10_in1[20]));
ADDFX1 inst_fa_1033_10_I21 (.CO(inst_fa_1033_10_out1[21]), .S(inst_fa_1033_10_out0[21]), .A(inst_fa_1033_10_in2[19]), .B(inst_fa_1033_10_in3[19]), .CI(inst_fa_1033_10_in1[21]));
ADDFX1 inst_fa_1033_10_I22 (.CO(inst_fa_1033_10_out1[22]), .S(inst_fa_1033_10_out0[22]), .A(inst_fa_1033_10_in2[20]), .B(inst_fa_1033_10_in3[20]), .CI(inst_fa_1033_10_in1[22]));
ADDFX1 inst_fa_1033_10_I23 (.CO(inst_fa_1033_10_out1[23]), .S(inst_fa_1033_10_out0[23]), .A(inst_fa_1033_10_in2[21]), .B(inst_fa_1033_10_in3[21]), .CI(inst_fa_1033_10_in1[23]));
ADDFX1 inst_fa_1033_10_I24 (.CO(inst_fa_1033_10_out1[24]), .S(inst_fa_1033_10_out0[24]), .A(inst_fa_1033_10_in2[22]), .B(inst_fa_1033_10_in3[22]), .CI(inst_fa_1033_10_in1[24]));
ADDFX1 inst_fa_1033_10_I25 (.CO(N231), .S(inst_fa_1033_10_out0[25]), .A(inst_fa_1033_10_in2[23]), .B(inst_fa_1033_10_in3[23]), .CI(inst_fa_1033_10_in1[25]));
assign inst_fa_1033_10_out0[0] = inst_fa_1033_10_in1[0];
assign inst_fa_1033_10_out0[1] = inst_fa_1033_10_in1[1];
assign inst_fa_1033_10_out1[0] = inst_fa_1033_10_in0;
assign inst_fa_1033_10_out1[1] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__31_2mx_bdw410776230_bdw (
	inst_cellmath__31_2mx_out0,
	inst_cellmath__31_2mx_in0,
	inst_cellmath__31_2mx_in1
	); /* architecture "gate_level" */ 
output [25:0] inst_cellmath__31_2mx_out0;
input [2:2] inst_cellmath__31_2mx_in0;
input [25:2] inst_cellmath__31_2mx_in1;
wire N270,N271;
INVXL inst_cellmath__31_2mx_I112 (.Y(N270), .A(inst_cellmath__31_2mx_in0[2]));
INVXL inst_cellmath__31_2mx_I113 (.Y(N271), .A(N270));
INVXL inst_cellmath__31_2mx_I111 (.Y(inst_cellmath__31_2mx_out0[1]), .A(N271));
MXI2XL inst_cellmath__31_2mx_I114 (.Y(inst_cellmath__31_2mx_out0[2]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[2]));
MXI2XL inst_cellmath__31_2mx_I115 (.Y(inst_cellmath__31_2mx_out0[3]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[3]));
MXI2XL inst_cellmath__31_2mx_I116 (.Y(inst_cellmath__31_2mx_out0[4]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[4]));
MXI2XL inst_cellmath__31_2mx_I117 (.Y(inst_cellmath__31_2mx_out0[5]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[5]));
MXI2XL inst_cellmath__31_2mx_I118 (.Y(inst_cellmath__31_2mx_out0[6]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[6]));
MXI2XL inst_cellmath__31_2mx_I119 (.Y(inst_cellmath__31_2mx_out0[7]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[7]));
MXI2XL inst_cellmath__31_2mx_I120 (.Y(inst_cellmath__31_2mx_out0[8]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[8]));
MXI2XL inst_cellmath__31_2mx_I121 (.Y(inst_cellmath__31_2mx_out0[9]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[9]));
MXI2XL inst_cellmath__31_2mx_I122 (.Y(inst_cellmath__31_2mx_out0[10]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[10]));
MXI2XL inst_cellmath__31_2mx_I123 (.Y(inst_cellmath__31_2mx_out0[11]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[11]));
MXI2XL inst_cellmath__31_2mx_I124 (.Y(inst_cellmath__31_2mx_out0[12]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[12]));
MXI2XL inst_cellmath__31_2mx_I125 (.Y(inst_cellmath__31_2mx_out0[13]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[13]));
MXI2XL inst_cellmath__31_2mx_I126 (.Y(inst_cellmath__31_2mx_out0[14]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[14]));
MXI2XL inst_cellmath__31_2mx_I127 (.Y(inst_cellmath__31_2mx_out0[15]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[15]));
MXI2XL inst_cellmath__31_2mx_I128 (.Y(inst_cellmath__31_2mx_out0[16]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[16]));
MXI2XL inst_cellmath__31_2mx_I129 (.Y(inst_cellmath__31_2mx_out0[17]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[17]));
MXI2XL inst_cellmath__31_2mx_I130 (.Y(inst_cellmath__31_2mx_out0[18]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[18]));
MXI2XL inst_cellmath__31_2mx_I131 (.Y(inst_cellmath__31_2mx_out0[19]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[19]));
MXI2XL inst_cellmath__31_2mx_I132 (.Y(inst_cellmath__31_2mx_out0[20]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[20]));
MXI2XL inst_cellmath__31_2mx_I133 (.Y(inst_cellmath__31_2mx_out0[21]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[21]));
MXI2XL inst_cellmath__31_2mx_I134 (.Y(inst_cellmath__31_2mx_out0[22]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[22]));
MXI2XL inst_cellmath__31_2mx_I135 (.Y(inst_cellmath__31_2mx_out0[23]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[23]));
MXI2XL inst_cellmath__31_2mx_I136 (.Y(inst_cellmath__31_2mx_out0[24]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[24]));
MXI2XL inst_cellmath__31_2mx_I137 (.Y(inst_cellmath__31_2mx_out0[25]), .A(N271), .B(inst_cellmath__31_2mx_out0[1]), .S0(inst_cellmath__31_2mx_in1[25]));
assign inst_cellmath__31_2mx_out0[0] = inst_cellmath__31_2mx_out0[1];
endmodule

module cynw_cm_float_div_ieee_inst_fa_1052_10_bdw410776230_bdw (
	inst_fa_1052_10_out0,
	inst_fa_1052_10_out1,
	inst_fa_1052_10_in0,
	inst_fa_1052_10_in1,
	inst_fa_1052_10_in2
	); /* architecture "gate_level" */ 
output [25:0] inst_fa_1052_10_out0;
output [24:0] inst_fa_1052_10_out1;
input [25:0] inst_fa_1052_10_in0;
input [24:0] inst_fa_1052_10_in1;
input [25:0] inst_fa_1052_10_in2;
wire N207;
ADDHX1 inst_fa_1052_10_I0 (.CO(inst_fa_1052_10_out1[0]), .S(inst_fa_1052_10_out0[0]), .A(inst_fa_1052_10_in0[0]), .B(inst_fa_1052_10_in2[0]));
ADDFX1 inst_fa_1052_10_I1 (.CO(inst_fa_1052_10_out1[1]), .S(inst_fa_1052_10_out0[1]), .A(inst_fa_1052_10_in1[0]), .B(inst_fa_1052_10_in0[1]), .CI(inst_fa_1052_10_in2[1]));
ADDFX1 inst_fa_1052_10_I2 (.CO(inst_fa_1052_10_out1[2]), .S(inst_fa_1052_10_out0[2]), .A(inst_fa_1052_10_in1[1]), .B(inst_fa_1052_10_in0[2]), .CI(inst_fa_1052_10_in2[2]));
ADDFX1 inst_fa_1052_10_I3 (.CO(inst_fa_1052_10_out1[3]), .S(inst_fa_1052_10_out0[3]), .A(inst_fa_1052_10_in1[2]), .B(inst_fa_1052_10_in0[3]), .CI(inst_fa_1052_10_in2[3]));
ADDFX1 inst_fa_1052_10_I4 (.CO(inst_fa_1052_10_out1[4]), .S(inst_fa_1052_10_out0[4]), .A(inst_fa_1052_10_in1[3]), .B(inst_fa_1052_10_in0[4]), .CI(inst_fa_1052_10_in2[4]));
ADDFX1 inst_fa_1052_10_I5 (.CO(inst_fa_1052_10_out1[5]), .S(inst_fa_1052_10_out0[5]), .A(inst_fa_1052_10_in1[4]), .B(inst_fa_1052_10_in0[5]), .CI(inst_fa_1052_10_in2[5]));
ADDFX1 inst_fa_1052_10_I6 (.CO(inst_fa_1052_10_out1[6]), .S(inst_fa_1052_10_out0[6]), .A(inst_fa_1052_10_in1[5]), .B(inst_fa_1052_10_in0[6]), .CI(inst_fa_1052_10_in2[6]));
ADDFX1 inst_fa_1052_10_I7 (.CO(inst_fa_1052_10_out1[7]), .S(inst_fa_1052_10_out0[7]), .A(inst_fa_1052_10_in1[6]), .B(inst_fa_1052_10_in0[7]), .CI(inst_fa_1052_10_in2[7]));
ADDFX1 inst_fa_1052_10_I8 (.CO(inst_fa_1052_10_out1[8]), .S(inst_fa_1052_10_out0[8]), .A(inst_fa_1052_10_in1[7]), .B(inst_fa_1052_10_in0[8]), .CI(inst_fa_1052_10_in2[8]));
ADDFX1 inst_fa_1052_10_I9 (.CO(inst_fa_1052_10_out1[9]), .S(inst_fa_1052_10_out0[9]), .A(inst_fa_1052_10_in1[8]), .B(inst_fa_1052_10_in0[9]), .CI(inst_fa_1052_10_in2[9]));
ADDFX1 inst_fa_1052_10_I10 (.CO(inst_fa_1052_10_out1[10]), .S(inst_fa_1052_10_out0[10]), .A(inst_fa_1052_10_in1[9]), .B(inst_fa_1052_10_in0[10]), .CI(inst_fa_1052_10_in2[10]));
ADDFX1 inst_fa_1052_10_I11 (.CO(inst_fa_1052_10_out1[11]), .S(inst_fa_1052_10_out0[11]), .A(inst_fa_1052_10_in1[10]), .B(inst_fa_1052_10_in0[11]), .CI(inst_fa_1052_10_in2[11]));
ADDFX1 inst_fa_1052_10_I12 (.CO(inst_fa_1052_10_out1[12]), .S(inst_fa_1052_10_out0[12]), .A(inst_fa_1052_10_in1[11]), .B(inst_fa_1052_10_in0[12]), .CI(inst_fa_1052_10_in2[12]));
ADDFX1 inst_fa_1052_10_I13 (.CO(inst_fa_1052_10_out1[13]), .S(inst_fa_1052_10_out0[13]), .A(inst_fa_1052_10_in1[12]), .B(inst_fa_1052_10_in0[13]), .CI(inst_fa_1052_10_in2[13]));
ADDFX1 inst_fa_1052_10_I14 (.CO(inst_fa_1052_10_out1[14]), .S(inst_fa_1052_10_out0[14]), .A(inst_fa_1052_10_in1[13]), .B(inst_fa_1052_10_in0[14]), .CI(inst_fa_1052_10_in2[14]));
ADDFX1 inst_fa_1052_10_I15 (.CO(inst_fa_1052_10_out1[15]), .S(inst_fa_1052_10_out0[15]), .A(inst_fa_1052_10_in1[14]), .B(inst_fa_1052_10_in0[15]), .CI(inst_fa_1052_10_in2[15]));
ADDFX1 inst_fa_1052_10_I16 (.CO(inst_fa_1052_10_out1[16]), .S(inst_fa_1052_10_out0[16]), .A(inst_fa_1052_10_in1[15]), .B(inst_fa_1052_10_in0[16]), .CI(inst_fa_1052_10_in2[16]));
ADDFX1 inst_fa_1052_10_I17 (.CO(inst_fa_1052_10_out1[17]), .S(inst_fa_1052_10_out0[17]), .A(inst_fa_1052_10_in1[16]), .B(inst_fa_1052_10_in0[17]), .CI(inst_fa_1052_10_in2[17]));
ADDFX1 inst_fa_1052_10_I18 (.CO(inst_fa_1052_10_out1[18]), .S(inst_fa_1052_10_out0[18]), .A(inst_fa_1052_10_in1[17]), .B(inst_fa_1052_10_in0[18]), .CI(inst_fa_1052_10_in2[18]));
ADDFX1 inst_fa_1052_10_I19 (.CO(inst_fa_1052_10_out1[19]), .S(inst_fa_1052_10_out0[19]), .A(inst_fa_1052_10_in1[18]), .B(inst_fa_1052_10_in0[19]), .CI(inst_fa_1052_10_in2[19]));
ADDFX1 inst_fa_1052_10_I20 (.CO(inst_fa_1052_10_out1[20]), .S(inst_fa_1052_10_out0[20]), .A(inst_fa_1052_10_in1[19]), .B(inst_fa_1052_10_in0[20]), .CI(inst_fa_1052_10_in2[20]));
ADDFX1 inst_fa_1052_10_I21 (.CO(inst_fa_1052_10_out1[21]), .S(inst_fa_1052_10_out0[21]), .A(inst_fa_1052_10_in1[20]), .B(inst_fa_1052_10_in0[21]), .CI(inst_fa_1052_10_in2[21]));
ADDFX1 inst_fa_1052_10_I22 (.CO(inst_fa_1052_10_out1[22]), .S(inst_fa_1052_10_out0[22]), .A(inst_fa_1052_10_in1[21]), .B(inst_fa_1052_10_in0[22]), .CI(inst_fa_1052_10_in2[22]));
ADDFX1 inst_fa_1052_10_I23 (.CO(inst_fa_1052_10_out1[23]), .S(inst_fa_1052_10_out0[23]), .A(inst_fa_1052_10_in1[22]), .B(inst_fa_1052_10_in0[23]), .CI(inst_fa_1052_10_in2[23]));
ADDFX1 inst_fa_1052_10_I24 (.CO(inst_fa_1052_10_out1[24]), .S(inst_fa_1052_10_out0[24]), .A(inst_fa_1052_10_in1[23]), .B(inst_fa_1052_10_in0[24]), .CI(inst_fa_1052_10_in2[24]));
ADDFX1 inst_fa_1052_10_I25 (.CO(N207), .S(inst_fa_1052_10_out0[25]), .A(inst_fa_1052_10_in1[24]), .B(inst_fa_1052_10_in0[25]), .CI(inst_fa_1052_10_in2[25]));
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__51_0_bdw410776230_bdw (
	inst_it2_cellmath__51_0_out0,
	inst_it2_cellmath__51_0_in0,
	inst_it2_cellmath__51_0_in1
	); /* architecture "gate_level" */ 
output [4:0] inst_it2_cellmath__51_0_out0;
input [25:21] inst_it2_cellmath__51_0_in0;
input [24:20] inst_it2_cellmath__51_0_in1;
wire N62,N66,N68,N70,N72;
ADDHX1 inst_it2_cellmath__51_0_I20 (.CO(N62), .S(inst_it2_cellmath__51_0_out0[0]), .A(inst_it2_cellmath__51_0_in1[20]), .B(inst_it2_cellmath__51_0_in0[21]));
ADDFX1 inst_it2_cellmath__51_0_I21 (.CO(N66), .S(inst_it2_cellmath__51_0_out0[1]), .A(inst_it2_cellmath__51_0_in0[22]), .B(inst_it2_cellmath__51_0_in1[21]), .CI(N62));
ADDFX1 inst_it2_cellmath__51_0_I22 (.CO(N68), .S(inst_it2_cellmath__51_0_out0[2]), .A(inst_it2_cellmath__51_0_in0[23]), .B(inst_it2_cellmath__51_0_in1[22]), .CI(N66));
ADDFX1 inst_it2_cellmath__51_0_I23 (.CO(N70), .S(inst_it2_cellmath__51_0_out0[3]), .A(inst_it2_cellmath__51_0_in0[24]), .B(inst_it2_cellmath__51_0_in1[23]), .CI(N68));
ADDFX1 inst_it2_cellmath__51_0_I24 (.CO(N72), .S(inst_it2_cellmath__51_0_out0[4]), .A(inst_it2_cellmath__51_0_in1[24]), .B(inst_it2_cellmath__51_0_in0[25]), .CI(N70));
endmodule

module cynw_cm_float_div_ieee_inst_it2_lookup1_cellmath__55_0_bdw410776230_bdw (
	inst_it2_lookup1_cellmath__55_0_out0,
	inst_it2_lookup1_cellmath__55_0_in0,
	inst_it2_lookup1_cellmath__55_0_in1
	); /* architecture "gate_level" */ 
output [2:0] inst_it2_lookup1_cellmath__55_0_out0;
input [4:0] inst_it2_lookup1_cellmath__55_0_in0;
input [22:21] inst_it2_lookup1_cellmath__55_0_in1;
wire N41,N116,N183,N212,N248,N252,N253 
	,N259,N263,N287,N379,N393,N457,N514,N519 
	,N525,N527,N530,N532,N533,N536,N798,N895 
	,N933,N934,N938,N939,N1005,N1007,N1038,N1046 
	,N1047,N1051,N1052,N1056,N1057,N1061,N1084,N1089 
	,N1093,N1096,N1099,N1119,N1126,N1133;
INVXL inst_it2_lookup1_cellmath__55_0_I848 (.Y(N1084), .A(inst_it2_lookup1_cellmath__55_0_in1[22]));
INVXL inst_it2_lookup1_cellmath__55_0_I20 (.Y(N41), .A(inst_it2_lookup1_cellmath__55_0_in1[21]));
INVXL inst_it2_lookup1_cellmath__55_0_I853 (.Y(N1089), .A(inst_it2_lookup1_cellmath__55_0_in0[0]));
INVXL inst_it2_lookup1_cellmath__55_0_I857 (.Y(N1093), .A(inst_it2_lookup1_cellmath__55_0_in0[1]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I81 (.Y(N116), .A(N1093), .B(N1089));
NOR2XL inst_it2_lookup1_cellmath__55_0_I133 (.Y(N183), .A(N1089), .B(N1084));
NAND2XL inst_it2_lookup1_cellmath__55_0_I157 (.Y(N212), .A(N41), .B(N1084));
AOI22XL inst_it2_lookup1_cellmath__55_0_I185 (.Y(N248), .A0(N1089), .A1(inst_it2_lookup1_cellmath__55_0_in1[22]), .B0(N212), .B1(inst_it2_lookup1_cellmath__55_0_in0[0]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I189 (.Y(N252), .A0(N1093), .A1(N248), .B0(N183), .B1(inst_it2_lookup1_cellmath__55_0_in0[1]));
NAND2XL hyperpropagate_3_1_A_I902 (.Y(N1119), .A(inst_it2_lookup1_cellmath__55_0_in1[22]), .B(inst_it2_lookup1_cellmath__55_0_in0[0]));
NOR2XL hyperpropagate_3_1_A_I903 (.Y(N253), .A(N1093), .B(N1119));
INVXL inst_it2_lookup1_cellmath__55_0_I860 (.Y(N1096), .A(inst_it2_lookup1_cellmath__55_0_in0[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I193 (.Y(N259), .A0(N1096), .A1(N252), .B0(N116), .B1(inst_it2_lookup1_cellmath__55_0_in0[2]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I195 (.Y(N263), .A(N116), .B(inst_it2_lookup1_cellmath__55_0_in0[2]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I217 (.Y(N287), .A(N41), .B(N1084));
NOR2XL inst_it2_lookup1_cellmath__55_0_I295 (.Y(N379), .A(inst_it2_lookup1_cellmath__55_0_in1[21]), .B(inst_it2_lookup1_cellmath__55_0_in1[22]));
NAND2XL hyperpropagate_3_1_A_I904 (.Y(N1126), .A(N1089), .B(N379));
NOR2XL hyperpropagate_3_1_A_I905 (.Y(N393), .A(inst_it2_lookup1_cellmath__55_0_in0[1]), .B(N1126));
AOI22XL inst_it2_lookup1_cellmath__55_0_I355 (.Y(N457), .A0(N1089), .A1(N1084), .B0(N379), .B1(inst_it2_lookup1_cellmath__55_0_in0[0]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I403 (.Y(N514), .A(inst_it2_lookup1_cellmath__55_0_in1[22]), .B(inst_it2_lookup1_cellmath__55_0_in1[21]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I407 (.Y(N519), .A0(N1089), .A1(N514), .B0(N1084), .B1(inst_it2_lookup1_cellmath__55_0_in0[0]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I411 (.Y(N525), .A0(N1093), .A1(N519), .B0(N457), .B1(inst_it2_lookup1_cellmath__55_0_in0[1]));
NAND4BXL inst_it2_lookup1_cellmath__55_0_I885 (.Y(N527), .AN(N1093), .B(N287), .C(inst_it2_lookup1_cellmath__55_0_in0[2]), .D(inst_it2_lookup1_cellmath__55_0_in0[0]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I415 (.Y(N530), .A0(N1096), .A1(N525), .B0(N393), .B1(inst_it2_lookup1_cellmath__55_0_in0[2]));
INVXL inst_it2_lookup1_cellmath__55_0_I863 (.Y(N1099), .A(inst_it2_lookup1_cellmath__55_0_in0[3]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I417 (.Y(N532), .A0(N1099), .A1(N527), .B0(N259), .B1(inst_it2_lookup1_cellmath__55_0_in0[3]));
NOR2XL andori2bb1_A_I906 (.Y(N1133), .A(inst_it2_lookup1_cellmath__55_0_in0[2]), .B(N253));
NOR2XL andori2bb1_A_I907 (.Y(N533), .A(N1133), .B(N1099));
AOI22XL inst_it2_lookup1_cellmath__55_0_I419 (.Y(N536), .A0(N1099), .A1(N530), .B0(N263), .B1(inst_it2_lookup1_cellmath__55_0_in0[3]));
NAND4BXL inst_it2_lookup1_cellmath__55_0_I888 (.Y(N798), .AN(inst_it2_lookup1_cellmath__55_0_in0[1]), .B(N287), .C(N1096), .D(N1089));
AOI22XL inst_it2_lookup1_cellmath__55_0_I713 (.Y(N895), .A0(N41), .A1(N1084), .B0(inst_it2_lookup1_cellmath__55_0_in1[22]), .B1(inst_it2_lookup1_cellmath__55_0_in1[21]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I741 (.Y(N933), .A0(N1089), .A1(N1084), .B0(N895), .B1(inst_it2_lookup1_cellmath__55_0_in0[0]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I742 (.Y(N934), .A0(N1089), .A1(inst_it2_lookup1_cellmath__55_0_in1[22]), .B0(N287), .B1(inst_it2_lookup1_cellmath__55_0_in0[0]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I745 (.Y(N938), .A0(N1093), .A1(N933), .B0(N1084), .B1(inst_it2_lookup1_cellmath__55_0_in0[1]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I746 (.Y(N939), .A(inst_it2_lookup1_cellmath__55_0_in0[1]), .B(N934));
NAND2XL inst_it2_lookup1_cellmath__55_0_I797 (.Y(N1005), .A(N379), .B(inst_it2_lookup1_cellmath__55_0_in0[0]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I798 (.Y(N1007), .A(N1089), .B(N212));
NOR2XL inst_it2_lookup1_cellmath__55_0_I819 (.Y(N1038), .A(N1089), .B(inst_it2_lookup1_cellmath__55_0_in1[22]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I823 (.Y(N1046), .A0(N1093), .A1(N1038), .B0(N1005), .B1(inst_it2_lookup1_cellmath__55_0_in0[1]));
NAND2XL inst_it2_lookup1_cellmath__55_0_I824 (.Y(N1047), .A(N1007), .B(inst_it2_lookup1_cellmath__55_0_in0[1]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I827 (.Y(N1051), .A0(N1096), .A1(N1046), .B0(N938), .B1(inst_it2_lookup1_cellmath__55_0_in0[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I828 (.Y(N1052), .A0(N1096), .A1(N1047), .B0(N939), .B1(inst_it2_lookup1_cellmath__55_0_in0[2]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I831 (.Y(N1056), .A0(N1099), .A1(N1051), .B0(N798), .B1(inst_it2_lookup1_cellmath__55_0_in0[3]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I832 (.Y(N1057), .A(inst_it2_lookup1_cellmath__55_0_in0[3]), .B(N1052));
INVXL inst_it2_lookup1_cellmath__55_0_I834 (.Y(N1061), .A(inst_it2_lookup1_cellmath__55_0_in0[4]));
AOI22XL inst_it2_lookup1_cellmath__55_0_I1038 (.Y(inst_it2_lookup1_cellmath__55_0_out0[0]), .A0(inst_it2_lookup1_cellmath__55_0_in0[4]), .A1(N532), .B0(N1061), .B1(N1056));
AOI22XL inst_it2_lookup1_cellmath__55_0_I836 (.Y(inst_it2_lookup1_cellmath__55_0_out0[1]), .A0(N1061), .A1(N1057), .B0(N533), .B1(inst_it2_lookup1_cellmath__55_0_in0[4]));
NOR2XL inst_it2_lookup1_cellmath__55_0_I837 (.Y(inst_it2_lookup1_cellmath__55_0_out0[2]), .A(N1061), .B(N536));
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__56__57__bdw410776230_bdw (
	inst_it2_cellmath__56__57__out0,
	inst_it2_cellmath__56__57__in0,
	inst_it2_cellmath__56__57__in1
	); /* architecture "gate_level" */ 
output [24:0] inst_it2_cellmath__56__57__out0;
input [0:0] inst_it2_cellmath__56__57__in0;
input [22:0] inst_it2_cellmath__56__57__in1;
wire N253;
INVXL inst_it2_cellmath__56__57__I54 (.Y(N253), .A(inst_it2_cellmath__56__57__in0[0]));
INVXL inst_it2_cellmath__56__57__I55 (.Y(inst_it2_cellmath__56__57__out0[24]), .A(N253));
AND2XL inst_it2_cellmath__56__57__I27 (.Y(inst_it2_cellmath__56__57__out0[1]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[0]));
AND2XL inst_it2_cellmath__56__57__I28 (.Y(inst_it2_cellmath__56__57__out0[2]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[1]));
AND2XL inst_it2_cellmath__56__57__I29 (.Y(inst_it2_cellmath__56__57__out0[3]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[2]));
AND2XL inst_it2_cellmath__56__57__I30 (.Y(inst_it2_cellmath__56__57__out0[4]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[3]));
AND2XL inst_it2_cellmath__56__57__I31 (.Y(inst_it2_cellmath__56__57__out0[5]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[4]));
AND2XL inst_it2_cellmath__56__57__I32 (.Y(inst_it2_cellmath__56__57__out0[6]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[5]));
AND2XL inst_it2_cellmath__56__57__I33 (.Y(inst_it2_cellmath__56__57__out0[7]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[6]));
AND2XL inst_it2_cellmath__56__57__I34 (.Y(inst_it2_cellmath__56__57__out0[8]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[7]));
AND2XL inst_it2_cellmath__56__57__I35 (.Y(inst_it2_cellmath__56__57__out0[9]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[8]));
AND2XL inst_it2_cellmath__56__57__I36 (.Y(inst_it2_cellmath__56__57__out0[10]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[9]));
AND2XL inst_it2_cellmath__56__57__I37 (.Y(inst_it2_cellmath__56__57__out0[11]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[10]));
AND2XL inst_it2_cellmath__56__57__I38 (.Y(inst_it2_cellmath__56__57__out0[12]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[11]));
AND2XL inst_it2_cellmath__56__57__I39 (.Y(inst_it2_cellmath__56__57__out0[13]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[12]));
AND2XL inst_it2_cellmath__56__57__I40 (.Y(inst_it2_cellmath__56__57__out0[14]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[13]));
AND2XL inst_it2_cellmath__56__57__I41 (.Y(inst_it2_cellmath__56__57__out0[15]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[14]));
AND2XL inst_it2_cellmath__56__57__I42 (.Y(inst_it2_cellmath__56__57__out0[16]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[15]));
AND2XL inst_it2_cellmath__56__57__I43 (.Y(inst_it2_cellmath__56__57__out0[17]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[16]));
AND2XL inst_it2_cellmath__56__57__I44 (.Y(inst_it2_cellmath__56__57__out0[18]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[17]));
AND2XL inst_it2_cellmath__56__57__I45 (.Y(inst_it2_cellmath__56__57__out0[19]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[18]));
AND2XL inst_it2_cellmath__56__57__I46 (.Y(inst_it2_cellmath__56__57__out0[20]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[19]));
AND2XL inst_it2_cellmath__56__57__I47 (.Y(inst_it2_cellmath__56__57__out0[21]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[20]));
AND2XL inst_it2_cellmath__56__57__I48 (.Y(inst_it2_cellmath__56__57__out0[22]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[21]));
AND2XL inst_it2_cellmath__56__57__I49 (.Y(inst_it2_cellmath__56__57__out0[23]), .A(inst_it2_cellmath__56__57__out0[24]), .B(inst_it2_cellmath__56__57__in1[22]));
assign inst_it2_cellmath__56__57__out0[0] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__57__61__bdw410776230_bdw (
	inst_it2_cellmath__57__61__out0,
	inst_it2_cellmath__57__61__in0,
	inst_it2_cellmath__57__61__in1
	); /* architecture "gate_level" */ 
output [25:0] inst_it2_cellmath__57__61__out0;
input [1:1] inst_it2_cellmath__57__61__in0;
input [22:0] inst_it2_cellmath__57__61__in1;
wire N402;
INVXL buf1_A_I127 (.Y(N402), .A(inst_it2_cellmath__57__61__in0[1]));
INVXL buf1_A_I128 (.Y(inst_it2_cellmath__57__61__out0[25]), .A(N402));
AND2XL inst_it2_cellmath__57__61__I29 (.Y(inst_it2_cellmath__57__61__out0[2]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[0]));
AND2XL inst_it2_cellmath__57__61__I30 (.Y(inst_it2_cellmath__57__61__out0[3]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[1]));
AND2XL inst_it2_cellmath__57__61__I31 (.Y(inst_it2_cellmath__57__61__out0[4]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[2]));
AND2XL inst_it2_cellmath__57__61__I32 (.Y(inst_it2_cellmath__57__61__out0[5]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[3]));
AND2XL inst_it2_cellmath__57__61__I33 (.Y(inst_it2_cellmath__57__61__out0[6]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[4]));
AND2XL inst_it2_cellmath__57__61__I34 (.Y(inst_it2_cellmath__57__61__out0[7]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[5]));
AND2XL inst_it2_cellmath__57__61__I35 (.Y(inst_it2_cellmath__57__61__out0[8]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[6]));
AND2XL inst_it2_cellmath__57__61__I36 (.Y(inst_it2_cellmath__57__61__out0[9]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[7]));
AND2XL inst_it2_cellmath__57__61__I37 (.Y(inst_it2_cellmath__57__61__out0[10]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[8]));
AND2XL inst_it2_cellmath__57__61__I38 (.Y(inst_it2_cellmath__57__61__out0[11]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[9]));
AND2XL inst_it2_cellmath__57__61__I39 (.Y(inst_it2_cellmath__57__61__out0[12]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[10]));
AND2XL inst_it2_cellmath__57__61__I40 (.Y(inst_it2_cellmath__57__61__out0[13]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[11]));
AND2XL inst_it2_cellmath__57__61__I41 (.Y(inst_it2_cellmath__57__61__out0[14]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[12]));
AND2XL inst_it2_cellmath__57__61__I42 (.Y(inst_it2_cellmath__57__61__out0[15]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[13]));
AND2XL inst_it2_cellmath__57__61__I43 (.Y(inst_it2_cellmath__57__61__out0[16]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[14]));
AND2XL inst_it2_cellmath__57__61__I44 (.Y(inst_it2_cellmath__57__61__out0[17]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[15]));
AND2XL inst_it2_cellmath__57__61__I45 (.Y(inst_it2_cellmath__57__61__out0[18]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[16]));
AND2XL inst_it2_cellmath__57__61__I46 (.Y(inst_it2_cellmath__57__61__out0[19]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[17]));
AND2XL inst_it2_cellmath__57__61__I47 (.Y(inst_it2_cellmath__57__61__out0[20]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[18]));
AND2XL inst_it2_cellmath__57__61__I48 (.Y(inst_it2_cellmath__57__61__out0[21]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[19]));
AND2XL inst_it2_cellmath__57__61__I49 (.Y(inst_it2_cellmath__57__61__out0[22]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[20]));
AND2XL inst_it2_cellmath__57__61__I50 (.Y(inst_it2_cellmath__57__61__out0[23]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[21]));
AND2XL inst_it2_cellmath__57__61__I51 (.Y(inst_it2_cellmath__57__61__out0[24]), .A(inst_it2_cellmath__57__61__out0[25]), .B(inst_it2_cellmath__57__61__in1[22]));
assign inst_it2_cellmath__57__61__out0[0] = 1'B0;
assign inst_it2_cellmath__57__61__out0[1] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__120_0_bdw410776230_bdw (
	inst_cellmath__120_0_out0,
	inst_cellmath__120_0_in0,
	inst_cellmath__120_0_in1
	); /* architecture "gate_level" */ 
output [25:0] inst_cellmath__120_0_out0;
input [25:0] inst_cellmath__120_0_in0,
	inst_cellmath__120_0_in1;
wire N251,N255,N257,N259,N261,N263,N265 
	,N267,N269,N271,N273,N275,N277,N279,N281 
	,N283,N285,N287,N289,N291,N293,N295,N297 
	,N299,N301,N303;
ADDHX1 inst_cellmath__120_0_I62 (.CO(N251), .S(inst_cellmath__120_0_out0[0]), .A(inst_cellmath__120_0_in1[0]), .B(inst_cellmath__120_0_in0[0]));
ADDFX1 inst_cellmath__120_0_I63 (.CO(N255), .S(inst_cellmath__120_0_out0[1]), .A(inst_cellmath__120_0_in0[1]), .B(inst_cellmath__120_0_in1[1]), .CI(N251));
ADDFX1 inst_cellmath__120_0_I64 (.CO(N257), .S(inst_cellmath__120_0_out0[2]), .A(inst_cellmath__120_0_in0[2]), .B(inst_cellmath__120_0_in1[2]), .CI(N255));
ADDFX1 inst_cellmath__120_0_I65 (.CO(N259), .S(inst_cellmath__120_0_out0[3]), .A(inst_cellmath__120_0_in0[3]), .B(inst_cellmath__120_0_in1[3]), .CI(N257));
ADDFX1 inst_cellmath__120_0_I66 (.CO(N261), .S(inst_cellmath__120_0_out0[4]), .A(inst_cellmath__120_0_in0[4]), .B(inst_cellmath__120_0_in1[4]), .CI(N259));
ADDFX1 inst_cellmath__120_0_I67 (.CO(N263), .S(inst_cellmath__120_0_out0[5]), .A(inst_cellmath__120_0_in0[5]), .B(inst_cellmath__120_0_in1[5]), .CI(N261));
ADDFX1 inst_cellmath__120_0_I68 (.CO(N265), .S(inst_cellmath__120_0_out0[6]), .A(inst_cellmath__120_0_in0[6]), .B(inst_cellmath__120_0_in1[6]), .CI(N263));
ADDFX1 inst_cellmath__120_0_I69 (.CO(N267), .S(inst_cellmath__120_0_out0[7]), .A(inst_cellmath__120_0_in0[7]), .B(inst_cellmath__120_0_in1[7]), .CI(N265));
ADDFX1 inst_cellmath__120_0_I70 (.CO(N269), .S(inst_cellmath__120_0_out0[8]), .A(inst_cellmath__120_0_in0[8]), .B(inst_cellmath__120_0_in1[8]), .CI(N267));
ADDFX1 inst_cellmath__120_0_I71 (.CO(N271), .S(inst_cellmath__120_0_out0[9]), .A(inst_cellmath__120_0_in0[9]), .B(inst_cellmath__120_0_in1[9]), .CI(N269));
ADDFX1 inst_cellmath__120_0_I72 (.CO(N273), .S(inst_cellmath__120_0_out0[10]), .A(inst_cellmath__120_0_in0[10]), .B(inst_cellmath__120_0_in1[10]), .CI(N271));
ADDFX1 inst_cellmath__120_0_I73 (.CO(N275), .S(inst_cellmath__120_0_out0[11]), .A(inst_cellmath__120_0_in0[11]), .B(inst_cellmath__120_0_in1[11]), .CI(N273));
ADDFX1 inst_cellmath__120_0_I74 (.CO(N277), .S(inst_cellmath__120_0_out0[12]), .A(inst_cellmath__120_0_in0[12]), .B(inst_cellmath__120_0_in1[12]), .CI(N275));
ADDFX1 inst_cellmath__120_0_I75 (.CO(N279), .S(inst_cellmath__120_0_out0[13]), .A(inst_cellmath__120_0_in0[13]), .B(inst_cellmath__120_0_in1[13]), .CI(N277));
ADDFX1 inst_cellmath__120_0_I76 (.CO(N281), .S(inst_cellmath__120_0_out0[14]), .A(inst_cellmath__120_0_in0[14]), .B(inst_cellmath__120_0_in1[14]), .CI(N279));
ADDFX1 inst_cellmath__120_0_I77 (.CO(N283), .S(inst_cellmath__120_0_out0[15]), .A(inst_cellmath__120_0_in0[15]), .B(inst_cellmath__120_0_in1[15]), .CI(N281));
ADDFX1 inst_cellmath__120_0_I78 (.CO(N285), .S(inst_cellmath__120_0_out0[16]), .A(inst_cellmath__120_0_in0[16]), .B(inst_cellmath__120_0_in1[16]), .CI(N283));
ADDFX1 inst_cellmath__120_0_I79 (.CO(N287), .S(inst_cellmath__120_0_out0[17]), .A(inst_cellmath__120_0_in0[17]), .B(inst_cellmath__120_0_in1[17]), .CI(N285));
ADDFX1 inst_cellmath__120_0_I80 (.CO(N289), .S(inst_cellmath__120_0_out0[18]), .A(inst_cellmath__120_0_in0[18]), .B(inst_cellmath__120_0_in1[18]), .CI(N287));
ADDFX1 inst_cellmath__120_0_I81 (.CO(N291), .S(inst_cellmath__120_0_out0[19]), .A(inst_cellmath__120_0_in0[19]), .B(inst_cellmath__120_0_in1[19]), .CI(N289));
ADDFX1 inst_cellmath__120_0_I82 (.CO(N293), .S(inst_cellmath__120_0_out0[20]), .A(inst_cellmath__120_0_in0[20]), .B(inst_cellmath__120_0_in1[20]), .CI(N291));
ADDFX1 inst_cellmath__120_0_I83 (.CO(N295), .S(inst_cellmath__120_0_out0[21]), .A(inst_cellmath__120_0_in1[21]), .B(inst_cellmath__120_0_in0[21]), .CI(N293));
ADDFX1 inst_cellmath__120_0_I84 (.CO(N297), .S(inst_cellmath__120_0_out0[22]), .A(inst_cellmath__120_0_in1[22]), .B(inst_cellmath__120_0_in0[22]), .CI(N295));
ADDFX1 inst_cellmath__120_0_I85 (.CO(N299), .S(inst_cellmath__120_0_out0[23]), .A(inst_cellmath__120_0_in1[23]), .B(inst_cellmath__120_0_in0[23]), .CI(N297));
ADDFX1 inst_cellmath__120_0_I86 (.CO(N301), .S(inst_cellmath__120_0_out0[24]), .A(inst_cellmath__120_0_in1[24]), .B(inst_cellmath__120_0_in0[24]), .CI(N299));
ADDFX1 inst_cellmath__120_0_I87 (.CO(N303), .S(inst_cellmath__120_0_out0[25]), .A(inst_cellmath__120_0_in1[25]), .B(inst_cellmath__120_0_in0[25]), .CI(N301));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__124_0_bdw410776230_bdw (
	inst_cellmath__124_0_out0,
	inst_cellmath__124_0_in0,
	inst_cellmath__124_0_in1,
	inst_cellmath__124_0_in2
	); /* architecture "gate_level" */ 
output [28:0] inst_cellmath__124_0_out0;
input [28:0] inst_cellmath__124_0_in0,
	inst_cellmath__124_0_in1;
input [25:25] inst_cellmath__124_0_in2;
MX2XL inst_cellmath__124_0_I58 (.Y(inst_cellmath__124_0_out0[0]), .A(inst_cellmath__124_0_in1[0]), .B(inst_cellmath__124_0_in0[0]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I59 (.Y(inst_cellmath__124_0_out0[1]), .A(inst_cellmath__124_0_in1[1]), .B(inst_cellmath__124_0_in0[1]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I60 (.Y(inst_cellmath__124_0_out0[2]), .A(inst_cellmath__124_0_in1[2]), .B(inst_cellmath__124_0_in0[2]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I61 (.Y(inst_cellmath__124_0_out0[3]), .A(inst_cellmath__124_0_in1[3]), .B(inst_cellmath__124_0_in0[3]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I62 (.Y(inst_cellmath__124_0_out0[4]), .A(inst_cellmath__124_0_in1[4]), .B(inst_cellmath__124_0_in0[4]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I63 (.Y(inst_cellmath__124_0_out0[5]), .A(inst_cellmath__124_0_in1[5]), .B(inst_cellmath__124_0_in0[5]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I64 (.Y(inst_cellmath__124_0_out0[6]), .A(inst_cellmath__124_0_in1[6]), .B(inst_cellmath__124_0_in0[6]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I65 (.Y(inst_cellmath__124_0_out0[7]), .A(inst_cellmath__124_0_in1[7]), .B(inst_cellmath__124_0_in0[7]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I66 (.Y(inst_cellmath__124_0_out0[8]), .A(inst_cellmath__124_0_in1[8]), .B(inst_cellmath__124_0_in0[8]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I67 (.Y(inst_cellmath__124_0_out0[9]), .A(inst_cellmath__124_0_in1[9]), .B(inst_cellmath__124_0_in0[9]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I68 (.Y(inst_cellmath__124_0_out0[10]), .A(inst_cellmath__124_0_in1[10]), .B(inst_cellmath__124_0_in0[10]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I69 (.Y(inst_cellmath__124_0_out0[11]), .A(inst_cellmath__124_0_in1[11]), .B(inst_cellmath__124_0_in0[11]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I70 (.Y(inst_cellmath__124_0_out0[12]), .A(inst_cellmath__124_0_in1[12]), .B(inst_cellmath__124_0_in0[12]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I71 (.Y(inst_cellmath__124_0_out0[13]), .A(inst_cellmath__124_0_in1[13]), .B(inst_cellmath__124_0_in0[13]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I72 (.Y(inst_cellmath__124_0_out0[14]), .A(inst_cellmath__124_0_in1[14]), .B(inst_cellmath__124_0_in0[14]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I73 (.Y(inst_cellmath__124_0_out0[15]), .A(inst_cellmath__124_0_in1[15]), .B(inst_cellmath__124_0_in0[15]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I74 (.Y(inst_cellmath__124_0_out0[16]), .A(inst_cellmath__124_0_in1[16]), .B(inst_cellmath__124_0_in0[16]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I75 (.Y(inst_cellmath__124_0_out0[17]), .A(inst_cellmath__124_0_in1[17]), .B(inst_cellmath__124_0_in0[17]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I76 (.Y(inst_cellmath__124_0_out0[18]), .A(inst_cellmath__124_0_in1[18]), .B(inst_cellmath__124_0_in0[18]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I77 (.Y(inst_cellmath__124_0_out0[19]), .A(inst_cellmath__124_0_in1[19]), .B(inst_cellmath__124_0_in0[19]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I78 (.Y(inst_cellmath__124_0_out0[20]), .A(inst_cellmath__124_0_in1[20]), .B(inst_cellmath__124_0_in0[20]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I79 (.Y(inst_cellmath__124_0_out0[21]), .A(inst_cellmath__124_0_in1[21]), .B(inst_cellmath__124_0_in0[21]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I80 (.Y(inst_cellmath__124_0_out0[22]), .A(inst_cellmath__124_0_in1[22]), .B(inst_cellmath__124_0_in0[22]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I81 (.Y(inst_cellmath__124_0_out0[23]), .A(inst_cellmath__124_0_in1[23]), .B(inst_cellmath__124_0_in0[23]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I82 (.Y(inst_cellmath__124_0_out0[24]), .A(inst_cellmath__124_0_in1[24]), .B(inst_cellmath__124_0_in0[24]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I83 (.Y(inst_cellmath__124_0_out0[25]), .A(inst_cellmath__124_0_in1[25]), .B(inst_cellmath__124_0_in0[25]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I84 (.Y(inst_cellmath__124_0_out0[26]), .A(inst_cellmath__124_0_in1[26]), .B(inst_cellmath__124_0_in0[26]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I85 (.Y(inst_cellmath__124_0_out0[27]), .A(inst_cellmath__124_0_in1[27]), .B(inst_cellmath__124_0_in0[27]), .S0(inst_cellmath__124_0_in2[25]));
MX2XL inst_cellmath__124_0_I86 (.Y(inst_cellmath__124_0_out0[28]), .A(inst_cellmath__124_0_in1[28]), .B(inst_cellmath__124_0_in0[28]), .S0(inst_cellmath__124_0_in2[25]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__125_0_bdw410776230_bdw (
	inst_cellmath__125_0_out0,
	inst_cellmath__125_0_in0,
	inst_cellmath__125_0_in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__125_0_out0;
input [27:4] inst_cellmath__125_0_in0;
input  inst_cellmath__125_0_in1;
wire N80,N83;
INVXL buf1_A_I31 (.Y(N83), .A(inst_cellmath__125_0_in1));
INVXL buf1_A_I32 (.Y(N80), .A(N83));
MX2XL inst_cellmath__125_0_I0 (.Y(inst_cellmath__125_0_out0[0]), .A(inst_cellmath__125_0_in0[5]), .B(inst_cellmath__125_0_in0[4]), .S0(N80));
MX2XL inst_cellmath__125_0_I1 (.Y(inst_cellmath__125_0_out0[1]), .A(inst_cellmath__125_0_in0[6]), .B(inst_cellmath__125_0_in0[5]), .S0(N80));
MX2XL inst_cellmath__125_0_I2 (.Y(inst_cellmath__125_0_out0[2]), .A(inst_cellmath__125_0_in0[7]), .B(inst_cellmath__125_0_in0[6]), .S0(N80));
MX2XL inst_cellmath__125_0_I3 (.Y(inst_cellmath__125_0_out0[3]), .A(inst_cellmath__125_0_in0[8]), .B(inst_cellmath__125_0_in0[7]), .S0(N80));
MX2XL inst_cellmath__125_0_I4 (.Y(inst_cellmath__125_0_out0[4]), .A(inst_cellmath__125_0_in0[9]), .B(inst_cellmath__125_0_in0[8]), .S0(N80));
MX2XL inst_cellmath__125_0_I5 (.Y(inst_cellmath__125_0_out0[5]), .A(inst_cellmath__125_0_in0[10]), .B(inst_cellmath__125_0_in0[9]), .S0(N80));
MX2XL inst_cellmath__125_0_I6 (.Y(inst_cellmath__125_0_out0[6]), .A(inst_cellmath__125_0_in0[11]), .B(inst_cellmath__125_0_in0[10]), .S0(N80));
MX2XL inst_cellmath__125_0_I7 (.Y(inst_cellmath__125_0_out0[7]), .A(inst_cellmath__125_0_in0[12]), .B(inst_cellmath__125_0_in0[11]), .S0(N80));
MX2XL inst_cellmath__125_0_I8 (.Y(inst_cellmath__125_0_out0[8]), .A(inst_cellmath__125_0_in0[13]), .B(inst_cellmath__125_0_in0[12]), .S0(N80));
MX2XL inst_cellmath__125_0_I9 (.Y(inst_cellmath__125_0_out0[9]), .A(inst_cellmath__125_0_in0[14]), .B(inst_cellmath__125_0_in0[13]), .S0(N80));
MX2XL inst_cellmath__125_0_I10 (.Y(inst_cellmath__125_0_out0[10]), .A(inst_cellmath__125_0_in0[15]), .B(inst_cellmath__125_0_in0[14]), .S0(N80));
MX2XL inst_cellmath__125_0_I11 (.Y(inst_cellmath__125_0_out0[11]), .A(inst_cellmath__125_0_in0[16]), .B(inst_cellmath__125_0_in0[15]), .S0(N80));
MX2XL inst_cellmath__125_0_I12 (.Y(inst_cellmath__125_0_out0[12]), .A(inst_cellmath__125_0_in0[17]), .B(inst_cellmath__125_0_in0[16]), .S0(N80));
MX2XL inst_cellmath__125_0_I13 (.Y(inst_cellmath__125_0_out0[13]), .A(inst_cellmath__125_0_in0[18]), .B(inst_cellmath__125_0_in0[17]), .S0(N80));
MX2XL inst_cellmath__125_0_I14 (.Y(inst_cellmath__125_0_out0[14]), .A(inst_cellmath__125_0_in0[19]), .B(inst_cellmath__125_0_in0[18]), .S0(N80));
MX2XL inst_cellmath__125_0_I15 (.Y(inst_cellmath__125_0_out0[15]), .A(inst_cellmath__125_0_in0[20]), .B(inst_cellmath__125_0_in0[19]), .S0(N80));
MX2XL inst_cellmath__125_0_I16 (.Y(inst_cellmath__125_0_out0[16]), .A(inst_cellmath__125_0_in0[21]), .B(inst_cellmath__125_0_in0[20]), .S0(N80));
MX2XL inst_cellmath__125_0_I17 (.Y(inst_cellmath__125_0_out0[17]), .A(inst_cellmath__125_0_in0[22]), .B(inst_cellmath__125_0_in0[21]), .S0(N80));
MX2XL inst_cellmath__125_0_I18 (.Y(inst_cellmath__125_0_out0[18]), .A(inst_cellmath__125_0_in0[23]), .B(inst_cellmath__125_0_in0[22]), .S0(N80));
MX2XL inst_cellmath__125_0_I19 (.Y(inst_cellmath__125_0_out0[19]), .A(inst_cellmath__125_0_in0[24]), .B(inst_cellmath__125_0_in0[23]), .S0(N80));
MX2XL inst_cellmath__125_0_I20 (.Y(inst_cellmath__125_0_out0[20]), .A(inst_cellmath__125_0_in0[25]), .B(inst_cellmath__125_0_in0[24]), .S0(N80));
MX2XL inst_cellmath__125_0_I21 (.Y(inst_cellmath__125_0_out0[21]), .A(inst_cellmath__125_0_in0[26]), .B(inst_cellmath__125_0_in0[25]), .S0(N80));
MX2XL inst_cellmath__125_0_I22 (.Y(inst_cellmath__125_0_out0[22]), .A(inst_cellmath__125_0_in0[27]), .B(inst_cellmath__125_0_in0[26]), .S0(N80));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__126_0_bdw410776230_bdw (
	inst_cellmath__126_0_out0,
	inst_cellmath__126_0_in0,
	inst_cellmath__126_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__126_0_out0;
input [4:3] inst_cellmath__126_0_in0;
input  inst_cellmath__126_0_in1;
MX2XL inst_cellmath__126_0_I2 (.Y(inst_cellmath__126_0_out0), .A(inst_cellmath__126_0_in0[4]), .B(inst_cellmath__126_0_in0[3]), .S0(inst_cellmath__126_0_in1));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__129_0_bdw410776230_bdw (
	inst_cellmath__129_0_out0,
	inst_cellmath__129_0_in0,
	inst_cellmath__129_0_in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__129_0_out0;
input  inst_cellmath__129_0_in0;
input [22:0] inst_cellmath__129_0_in1;
wire N136,N140,N144,N148,N152,N156,N160 
	,N164,N168,N172,N176,N180,N184,N188,N192 
	,N196,N200,N204,N208,N212,N216,N220;
ADDHX1 inst_cellmath__129_0_I34 (.CO(N136), .S(inst_cellmath__129_0_out0[0]), .A(inst_cellmath__129_0_in0), .B(inst_cellmath__129_0_in1[0]));
ADDHX1 inst_cellmath__129_0_I35 (.CO(N140), .S(inst_cellmath__129_0_out0[1]), .A(inst_cellmath__129_0_in1[1]), .B(N136));
ADDHX1 inst_cellmath__129_0_I36 (.CO(N144), .S(inst_cellmath__129_0_out0[2]), .A(inst_cellmath__129_0_in1[2]), .B(N140));
ADDHX1 inst_cellmath__129_0_I37 (.CO(N148), .S(inst_cellmath__129_0_out0[3]), .A(inst_cellmath__129_0_in1[3]), .B(N144));
ADDHX1 inst_cellmath__129_0_I38 (.CO(N152), .S(inst_cellmath__129_0_out0[4]), .A(inst_cellmath__129_0_in1[4]), .B(N148));
ADDHX1 inst_cellmath__129_0_I39 (.CO(N156), .S(inst_cellmath__129_0_out0[5]), .A(inst_cellmath__129_0_in1[5]), .B(N152));
ADDHX1 inst_cellmath__129_0_I40 (.CO(N160), .S(inst_cellmath__129_0_out0[6]), .A(inst_cellmath__129_0_in1[6]), .B(N156));
ADDHX1 inst_cellmath__129_0_I41 (.CO(N164), .S(inst_cellmath__129_0_out0[7]), .A(inst_cellmath__129_0_in1[7]), .B(N160));
ADDHX1 inst_cellmath__129_0_I42 (.CO(N168), .S(inst_cellmath__129_0_out0[8]), .A(inst_cellmath__129_0_in1[8]), .B(N164));
ADDHX1 inst_cellmath__129_0_I43 (.CO(N172), .S(inst_cellmath__129_0_out0[9]), .A(inst_cellmath__129_0_in1[9]), .B(N168));
ADDHX1 inst_cellmath__129_0_I44 (.CO(N176), .S(inst_cellmath__129_0_out0[10]), .A(inst_cellmath__129_0_in1[10]), .B(N172));
ADDHX1 inst_cellmath__129_0_I45 (.CO(N180), .S(inst_cellmath__129_0_out0[11]), .A(inst_cellmath__129_0_in1[11]), .B(N176));
ADDHX1 inst_cellmath__129_0_I46 (.CO(N184), .S(inst_cellmath__129_0_out0[12]), .A(inst_cellmath__129_0_in1[12]), .B(N180));
ADDHX1 inst_cellmath__129_0_I47 (.CO(N188), .S(inst_cellmath__129_0_out0[13]), .A(inst_cellmath__129_0_in1[13]), .B(N184));
ADDHX1 inst_cellmath__129_0_I48 (.CO(N192), .S(inst_cellmath__129_0_out0[14]), .A(inst_cellmath__129_0_in1[14]), .B(N188));
ADDHX1 inst_cellmath__129_0_I49 (.CO(N196), .S(inst_cellmath__129_0_out0[15]), .A(inst_cellmath__129_0_in1[15]), .B(N192));
ADDHX1 inst_cellmath__129_0_I50 (.CO(N200), .S(inst_cellmath__129_0_out0[16]), .A(inst_cellmath__129_0_in1[16]), .B(N196));
ADDHX1 inst_cellmath__129_0_I51 (.CO(N204), .S(inst_cellmath__129_0_out0[17]), .A(inst_cellmath__129_0_in1[17]), .B(N200));
ADDHX1 inst_cellmath__129_0_I52 (.CO(N208), .S(inst_cellmath__129_0_out0[18]), .A(inst_cellmath__129_0_in1[18]), .B(N204));
ADDHX1 inst_cellmath__129_0_I53 (.CO(N212), .S(inst_cellmath__129_0_out0[19]), .A(inst_cellmath__129_0_in1[19]), .B(N208));
ADDHX1 inst_cellmath__129_0_I54 (.CO(N216), .S(inst_cellmath__129_0_out0[20]), .A(inst_cellmath__129_0_in1[20]), .B(N212));
ADDHX1 inst_cellmath__129_0_I55 (.CO(N220), .S(inst_cellmath__129_0_out0[21]), .A(inst_cellmath__129_0_in1[21]), .B(N216));
XOR2XL inst_cellmath__129_0_I56 (.Y(inst_cellmath__129_0_out0[22]), .A(inst_cellmath__129_0_in1[22]), .B(N220));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__127__104__bdw410776230_bdw (
	inst_cellmath__127__104__out0,
	inst_cellmath__127__104__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__127__104__out0;
input [3:0] inst_cellmath__127__104__in0;
wire N7,N8;
NOR2XL inst_cellmath__127__104__I0 (.Y(N7), .A(inst_cellmath__127__104__in0[0]), .B(inst_cellmath__127__104__in0[1]));
NOR2XL inst_cellmath__127__104__I1 (.Y(N8), .A(inst_cellmath__127__104__in0[3]), .B(inst_cellmath__127__104__in0[2]));
NAND2XL inst_cellmath__127__104__I2 (.Y(inst_cellmath__127__104__out0[0]), .A(N7), .B(N8));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__127__103__bdw410776230_bdw (
	inst_cellmath__127__103__out0,
	inst_cellmath__127__103__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__127__103__out0;
input [2:0] inst_cellmath__127__103__in0;
OR3XL inst_cellmath__127__103__I3 (.Y(inst_cellmath__127__103__out0[0]), .A(inst_cellmath__127__103__in0[0]), .B(inst_cellmath__127__103__in0[1]), .C(inst_cellmath__127__103__in0[2]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__127_0_bdw410776230_bdw (
	inst_cellmath__127_0_out0,
	inst_cellmath__127_0_in0,
	inst_cellmath__127_0_in1,
	inst_cellmath__127_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__127_0_out0;
input [0:0] inst_cellmath__127_0_in0,
	inst_cellmath__127_0_in1;
input  inst_cellmath__127_0_in2;
MX2XL inst_cellmath__127_0_I2 (.Y(inst_cellmath__127_0_out0), .A(inst_cellmath__127_0_in0[0]), .B(inst_cellmath__127_0_in1[0]), .S0(inst_cellmath__127_0_in2));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__130__105__bdw410776230_bdw (
	inst_cellmath__130__105__out0,
	inst_cellmath__130__105__in0,
	inst_cellmath__130__105__in1,
	inst_cellmath__130__105__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__130__105__out0;
input  inst_cellmath__130__105__in0;
input [0:0] inst_cellmath__130__105__in1;
input [25:0] inst_cellmath__130__105__in2;
wire N36,N44,N45,N47,N49,N50,N51 
	,N52,N53,N54,N59,N60,N61,N62,N66 
	;
NOR4X1 inst_cellmath__130__105__I39 (.Y(N36), .A(inst_cellmath__130__105__in2[0]), .B(inst_cellmath__130__105__in2[1]), .C(inst_cellmath__130__105__in2[2]), .D(inst_cellmath__130__105__in2[6]));
NOR3XL inst_cellmath__130__105__I41 (.Y(N44), .A(inst_cellmath__130__105__in2[5]), .B(inst_cellmath__130__105__in2[11]), .C(inst_cellmath__130__105__in2[15]));
NOR3BXL inst_cellmath__130__105__I42 (.Y(N45), .AN(N36), .B(inst_cellmath__130__105__in2[14]), .C(inst_cellmath__130__105__in2[12]));
NOR3XL inst_cellmath__130__105__I43 (.Y(N47), .A(inst_cellmath__130__105__in2[10]), .B(inst_cellmath__130__105__in2[8]), .C(inst_cellmath__130__105__in2[9]));
NOR3XL inst_cellmath__130__105__I44 (.Y(N49), .A(inst_cellmath__130__105__in2[13]), .B(inst_cellmath__130__105__in2[16]), .C(inst_cellmath__130__105__in2[19]));
NOR2XL inst_cellmath__130__105__I19 (.Y(N50), .A(inst_cellmath__130__105__in2[20]), .B(inst_cellmath__130__105__in2[18]));
NOR4X1 inst_cellmath__130__105__I45 (.Y(N51), .A(inst_cellmath__130__105__in2[4]), .B(inst_cellmath__130__105__in2[3]), .C(inst_cellmath__130__105__in2[7]), .D(inst_cellmath__130__105__in2[17]));
NOR2XL inst_cellmath__130__105__I21 (.Y(N52), .A(inst_cellmath__130__105__in2[22]), .B(inst_cellmath__130__105__in2[24]));
NOR2XL inst_cellmath__130__105__I22 (.Y(N53), .A(inst_cellmath__130__105__in2[21]), .B(inst_cellmath__130__105__in2[23]));
NAND2XL inst_cellmath__130__105__I23 (.Y(N54), .A(N45), .B(N44));
NAND2XL inst_cellmath__130__105__I26 (.Y(N61), .A(N53), .B(N49));
NOR2XL inst_cellmath__130__105__I28 (.Y(N59), .A(inst_cellmath__130__105__in2[25]), .B(N54));
NAND4XL inst_cellmath__130__105__I48 (.Y(N60), .A(N47), .B(N50), .C(N51), .D(N52));
NOR2XL inst_cellmath__130__105__I31 (.Y(N62), .A(N61), .B(N60));
NAND3BXL inst_cellmath__130__105__I47 (.Y(N66), .AN(inst_cellmath__130__105__in0), .B(N59), .C(N62));
OR2XL inst_cellmath__130__105__I36 (.Y(inst_cellmath__130__105__out0[0]), .A(N66), .B(inst_cellmath__130__105__in1[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__121__106__bdw410776230_bdw (
	inst_cellmath__121__106__out0,
	inst_cellmath__121__106__in0,
	inst_cellmath__121__106__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__121__106__out0;
input [0:0] inst_cellmath__121__106__in0,
	inst_cellmath__121__106__in1;
AND2XL inst_cellmath__121__106__I0 (.Y(inst_cellmath__121__106__out0[0]), .A(inst_cellmath__121__106__in0[0]), .B(inst_cellmath__121__106__in1[0]));
endmodule

`ifdef arith_fdrq_A_bdw410776230_bdw_COMPILED
`else
`define arith_fdrq_A_bdw410776230_bdw_COMPILED
module arith_fdrq_A_bdw410776230_bdw (
	r,
	d,
	clk,
	q
	); /* architecture "gate_level" */ 
input  r,
	d;
input  clk;
output  q;
wire  data;
DFFQXL arith_fdrq_A_I0 (.Q(q), .D(data), .CK(clk));
AND2XL arith_fdrq_A_I1 (.Y(data), .A(d), .B(r));
endmodule
`endif //  `ifdef arith_fdrq_A_bdw410776230_bdw_COMPILED

module cynw_cm_float_div_ieee_inst_cellmath__12__18__bdw410776230_bdw (
	inst_cellmath__12__18__out0,
	inst_cellmath__12__18__in0
	); /* architecture "gate_level" */ 
output [3:0] inst_cellmath__12__18__out0;
input [3:0] inst_cellmath__12__18__in0;
wire N44,N48;
INVXL inst_cellmath__12__18__I15 (.Y(inst_cellmath__12__18__out0[0]), .A(inst_cellmath__12__18__in0[0]));
ADDHX1 inst_cellmath__12__18__I16 (.CO(N44), .S(inst_cellmath__12__18__out0[1]), .A(inst_cellmath__12__18__in0[1]), .B(inst_cellmath__12__18__in0[0]));
ADDHX1 inst_cellmath__12__18__I17 (.CO(N48), .S(inst_cellmath__12__18__out0[2]), .A(inst_cellmath__12__18__in0[2]), .B(N44));
XOR2XL inst_cellmath__12__18__I18 (.Y(inst_cellmath__12__18__out0[3]), .A(inst_cellmath__12__18__in0[3]), .B(N48));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__12__19__bdw410776230_bdw (
	inst_cellmath__12__19__out0,
	inst_cellmath__12__19__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__12__19__out0;
input [3:0] inst_cellmath__12__19__in0;
wire N7,N8;
NAND2XL inst_cellmath__12__19__I0 (.Y(N7), .A(inst_cellmath__12__19__in0[3]), .B(inst_cellmath__12__19__in0[0]));
NAND2XL inst_cellmath__12__19__I1 (.Y(N8), .A(inst_cellmath__12__19__in0[2]), .B(inst_cellmath__12__19__in0[1]));
NOR2XL inst_cellmath__12__19__I2 (.Y(inst_cellmath__12__19__out0[0]), .A(N7), .B(N8));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__12_0_bdw410776230_bdw (
	inst_cellmath__12_0_out0,
	inst_cellmath__12_0_in0,
	inst_cellmath__12_0_in1
	); /* architecture "gate_level" */ 
output [3:0] inst_cellmath__12_0_out0;
input [0:0] inst_cellmath__12_0_in0;
input [3:0] inst_cellmath__12_0_in1;
OR2XL inst_cellmath__12_0_I9 (.Y(inst_cellmath__12_0_out0[0]), .A(inst_cellmath__12_0_in0[0]), .B(inst_cellmath__12_0_in1[0]));
OR2XL inst_cellmath__12_0_I10 (.Y(inst_cellmath__12_0_out0[1]), .A(inst_cellmath__12_0_in0[0]), .B(inst_cellmath__12_0_in1[1]));
OR2XL inst_cellmath__12_0_I11 (.Y(inst_cellmath__12_0_out0[2]), .A(inst_cellmath__12_0_in0[0]), .B(inst_cellmath__12_0_in1[2]));
OR2XL inst_cellmath__12_0_I12 (.Y(inst_cellmath__12_0_out0[3]), .A(inst_cellmath__12_0_in0[0]), .B(inst_cellmath__12_0_in1[3]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__46_0_bdw410776230_bdw (
	inst_cellmath__46_0_out0,
	inst_cellmath__46_0_in0,
	inst_cellmath__46_0_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__46_0_out0;
input [24:0] inst_cellmath__46_0_in0;
input  inst_cellmath__46_0_in1;
wire N155;
INVXL inst_cellmath__46_0_I51 (.Y(N155), .A(inst_cellmath__46_0_in1));
NAND2BXL inst_cellmath__46_0_I1 (.Y(inst_cellmath__46_0_out0[0]), .AN(inst_cellmath__46_0_in0[0]), .B(N155));
AND2XL inst_cellmath__46_0_I2 (.Y(inst_cellmath__46_0_out0[1]), .A(N155), .B(inst_cellmath__46_0_in0[1]));
AND2XL inst_cellmath__46_0_I3 (.Y(inst_cellmath__46_0_out0[2]), .A(N155), .B(inst_cellmath__46_0_in0[2]));
AND2XL inst_cellmath__46_0_I4 (.Y(inst_cellmath__46_0_out0[3]), .A(N155), .B(inst_cellmath__46_0_in0[3]));
AND2XL inst_cellmath__46_0_I5 (.Y(inst_cellmath__46_0_out0[4]), .A(N155), .B(inst_cellmath__46_0_in0[4]));
AND2XL inst_cellmath__46_0_I6 (.Y(inst_cellmath__46_0_out0[5]), .A(N155), .B(inst_cellmath__46_0_in0[5]));
AND2XL inst_cellmath__46_0_I7 (.Y(inst_cellmath__46_0_out0[6]), .A(N155), .B(inst_cellmath__46_0_in0[6]));
AND2XL inst_cellmath__46_0_I8 (.Y(inst_cellmath__46_0_out0[7]), .A(N155), .B(inst_cellmath__46_0_in0[7]));
AND2XL inst_cellmath__46_0_I9 (.Y(inst_cellmath__46_0_out0[8]), .A(N155), .B(inst_cellmath__46_0_in0[8]));
AND2XL inst_cellmath__46_0_I10 (.Y(inst_cellmath__46_0_out0[9]), .A(N155), .B(inst_cellmath__46_0_in0[9]));
AND2XL inst_cellmath__46_0_I11 (.Y(inst_cellmath__46_0_out0[10]), .A(N155), .B(inst_cellmath__46_0_in0[10]));
AND2XL inst_cellmath__46_0_I12 (.Y(inst_cellmath__46_0_out0[11]), .A(N155), .B(inst_cellmath__46_0_in0[11]));
AND2XL inst_cellmath__46_0_I13 (.Y(inst_cellmath__46_0_out0[12]), .A(N155), .B(inst_cellmath__46_0_in0[12]));
AND2XL inst_cellmath__46_0_I14 (.Y(inst_cellmath__46_0_out0[13]), .A(N155), .B(inst_cellmath__46_0_in0[13]));
AND2XL inst_cellmath__46_0_I15 (.Y(inst_cellmath__46_0_out0[14]), .A(N155), .B(inst_cellmath__46_0_in0[14]));
AND2XL inst_cellmath__46_0_I16 (.Y(inst_cellmath__46_0_out0[15]), .A(N155), .B(inst_cellmath__46_0_in0[15]));
AND2XL inst_cellmath__46_0_I17 (.Y(inst_cellmath__46_0_out0[16]), .A(N155), .B(inst_cellmath__46_0_in0[16]));
AND2XL inst_cellmath__46_0_I18 (.Y(inst_cellmath__46_0_out0[17]), .A(N155), .B(inst_cellmath__46_0_in0[17]));
AND2XL inst_cellmath__46_0_I19 (.Y(inst_cellmath__46_0_out0[18]), .A(N155), .B(inst_cellmath__46_0_in0[18]));
AND2XL inst_cellmath__46_0_I20 (.Y(inst_cellmath__46_0_out0[19]), .A(N155), .B(inst_cellmath__46_0_in0[19]));
AND2XL inst_cellmath__46_0_I21 (.Y(inst_cellmath__46_0_out0[20]), .A(N155), .B(inst_cellmath__46_0_in0[20]));
AND2XL inst_cellmath__46_0_I22 (.Y(inst_cellmath__46_0_out0[21]), .A(N155), .B(inst_cellmath__46_0_in0[21]));
AND2XL inst_cellmath__46_0_I23 (.Y(inst_cellmath__46_0_out0[22]), .A(N155), .B(inst_cellmath__46_0_in0[22]));
AND2XL inst_cellmath__46_0_I24 (.Y(inst_cellmath__46_0_out0[23]), .A(N155), .B(inst_cellmath__46_0_in0[23]));
AND2XL inst_cellmath__46_0_I25 (.Y(inst_cellmath__46_0_out0[24]), .A(N155), .B(inst_cellmath__46_0_in0[24]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__47_0_bdw410776230_bdw (
	inst_cellmath__47_0_out0,
	inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__47_0_out0;
input [24:0] inst_cellmath__47_0_in0;
input  inst_cellmath__47_0_in1;
wire N205,N212;
INVXL inst_cellmath__47_0_I51 (.Y(N205), .A(inst_cellmath__47_0_in1));
INVXL inst_cellmath__47_0_I58 (.Y(N212), .A(N205));
NOR2BX1 inst_cellmath__47_0_I241 (.Y(inst_cellmath__47_0_out0[0]), .AN(inst_cellmath__47_0_in0[0]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I242 (.Y(inst_cellmath__47_0_out0[1]), .AN(inst_cellmath__47_0_in0[1]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I243 (.Y(inst_cellmath__47_0_out0[2]), .AN(inst_cellmath__47_0_in0[2]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I244 (.Y(inst_cellmath__47_0_out0[3]), .AN(inst_cellmath__47_0_in0[3]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I245 (.Y(inst_cellmath__47_0_out0[4]), .AN(inst_cellmath__47_0_in0[4]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I246 (.Y(inst_cellmath__47_0_out0[5]), .AN(inst_cellmath__47_0_in0[5]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I247 (.Y(inst_cellmath__47_0_out0[6]), .AN(inst_cellmath__47_0_in0[6]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I248 (.Y(inst_cellmath__47_0_out0[7]), .AN(inst_cellmath__47_0_in0[7]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I249 (.Y(inst_cellmath__47_0_out0[8]), .AN(inst_cellmath__47_0_in0[8]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I250 (.Y(inst_cellmath__47_0_out0[9]), .AN(inst_cellmath__47_0_in0[9]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I251 (.Y(inst_cellmath__47_0_out0[10]), .AN(inst_cellmath__47_0_in0[10]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I252 (.Y(inst_cellmath__47_0_out0[11]), .AN(inst_cellmath__47_0_in0[11]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I253 (.Y(inst_cellmath__47_0_out0[12]), .AN(inst_cellmath__47_0_in0[12]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I254 (.Y(inst_cellmath__47_0_out0[13]), .AN(inst_cellmath__47_0_in0[13]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I255 (.Y(inst_cellmath__47_0_out0[14]), .AN(inst_cellmath__47_0_in0[14]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I256 (.Y(inst_cellmath__47_0_out0[15]), .AN(inst_cellmath__47_0_in0[15]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I257 (.Y(inst_cellmath__47_0_out0[16]), .AN(inst_cellmath__47_0_in0[16]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I258 (.Y(inst_cellmath__47_0_out0[17]), .AN(inst_cellmath__47_0_in0[17]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I259 (.Y(inst_cellmath__47_0_out0[18]), .AN(inst_cellmath__47_0_in0[18]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I260 (.Y(inst_cellmath__47_0_out0[19]), .AN(inst_cellmath__47_0_in0[19]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I261 (.Y(inst_cellmath__47_0_out0[20]), .AN(inst_cellmath__47_0_in0[20]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I262 (.Y(inst_cellmath__47_0_out0[21]), .AN(inst_cellmath__47_0_in0[21]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I263 (.Y(inst_cellmath__47_0_out0[22]), .AN(inst_cellmath__47_0_in0[22]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I264 (.Y(inst_cellmath__47_0_out0[23]), .AN(inst_cellmath__47_0_in0[23]), .B(N212));
NOR2BX1 inst_cellmath__47_0_I265 (.Y(inst_cellmath__47_0_out0[24]), .AN(inst_cellmath__47_0_in0[24]), .B(N212));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__48__47__bdw410776230_bdw (
	inst_cellmath__48__47__out0,
	inst_cellmath__48__47__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__48__47__out0;
input [1:0] inst_cellmath__48__47__in0;
NAND2XL inst_cellmath__48__47__I0 (.Y(inst_cellmath__48__47__out0[0]), .A(inst_cellmath__48__47__in0[1]), .B(inst_cellmath__48__47__in0[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__48__44__bdw410776230_bdw (
	inst_cellmath__48__44__out0,
	inst_cellmath__48__44__in0,
	inst_cellmath__48__44__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__48__44__out0;
input [2:1] inst_cellmath__48__44__in0;
input [0:0] inst_cellmath__48__44__in1;
MX2XL inst_cellmath__48__44__I2 (.Y(inst_cellmath__48__44__out0[0]), .A(inst_cellmath__48__44__in0[1]), .B(inst_cellmath__48__44__in1[0]), .S0(inst_cellmath__48__44__in0[2]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__42_0_bdw410776230_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3,
	inst_cellmath__42_0_in4
	); /* architecture "gate_level" */ 
output [26:0] inst_cellmath__42_0_out0;
input [0:0] inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1;
input [24:0] inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3;
input  inst_cellmath__42_0_in4;
wire N361;
BUFX2 inst_cellmath__42_0_I90 (.Y(N361), .A(inst_cellmath__42_0_in4));
MX2XL inst_cellmath__42_0_I56 (.Y(inst_cellmath__42_0_out0[2]), .A(inst_cellmath__42_0_in2[0]), .B(inst_cellmath__42_0_in3[0]), .S0(N361));
MX2XL inst_cellmath__42_0_I57 (.Y(inst_cellmath__42_0_out0[3]), .A(inst_cellmath__42_0_in2[1]), .B(inst_cellmath__42_0_in3[1]), .S0(N361));
MX2XL inst_cellmath__42_0_I58 (.Y(inst_cellmath__42_0_out0[4]), .A(inst_cellmath__42_0_in2[2]), .B(inst_cellmath__42_0_in3[2]), .S0(N361));
MX2XL inst_cellmath__42_0_I59 (.Y(inst_cellmath__42_0_out0[5]), .A(inst_cellmath__42_0_in2[3]), .B(inst_cellmath__42_0_in3[3]), .S0(N361));
MX2XL inst_cellmath__42_0_I60 (.Y(inst_cellmath__42_0_out0[6]), .A(inst_cellmath__42_0_in2[4]), .B(inst_cellmath__42_0_in3[4]), .S0(N361));
MX2XL inst_cellmath__42_0_I61 (.Y(inst_cellmath__42_0_out0[7]), .A(inst_cellmath__42_0_in2[5]), .B(inst_cellmath__42_0_in3[5]), .S0(N361));
MX2XL inst_cellmath__42_0_I62 (.Y(inst_cellmath__42_0_out0[8]), .A(inst_cellmath__42_0_in2[6]), .B(inst_cellmath__42_0_in3[6]), .S0(N361));
MX2XL inst_cellmath__42_0_I63 (.Y(inst_cellmath__42_0_out0[9]), .A(inst_cellmath__42_0_in2[7]), .B(inst_cellmath__42_0_in3[7]), .S0(N361));
MX2XL inst_cellmath__42_0_I64 (.Y(inst_cellmath__42_0_out0[10]), .A(inst_cellmath__42_0_in2[8]), .B(inst_cellmath__42_0_in3[8]), .S0(N361));
MX2XL inst_cellmath__42_0_I65 (.Y(inst_cellmath__42_0_out0[11]), .A(inst_cellmath__42_0_in2[9]), .B(inst_cellmath__42_0_in3[9]), .S0(N361));
MX2XL inst_cellmath__42_0_I66 (.Y(inst_cellmath__42_0_out0[12]), .A(inst_cellmath__42_0_in2[10]), .B(inst_cellmath__42_0_in3[10]), .S0(N361));
MX2XL inst_cellmath__42_0_I67 (.Y(inst_cellmath__42_0_out0[13]), .A(inst_cellmath__42_0_in2[11]), .B(inst_cellmath__42_0_in3[11]), .S0(N361));
MX2XL inst_cellmath__42_0_I68 (.Y(inst_cellmath__42_0_out0[14]), .A(inst_cellmath__42_0_in2[12]), .B(inst_cellmath__42_0_in3[12]), .S0(N361));
MX2XL inst_cellmath__42_0_I69 (.Y(inst_cellmath__42_0_out0[15]), .A(inst_cellmath__42_0_in2[13]), .B(inst_cellmath__42_0_in3[13]), .S0(N361));
MX2XL inst_cellmath__42_0_I70 (.Y(inst_cellmath__42_0_out0[16]), .A(inst_cellmath__42_0_in2[14]), .B(inst_cellmath__42_0_in3[14]), .S0(N361));
MX2XL inst_cellmath__42_0_I71 (.Y(inst_cellmath__42_0_out0[17]), .A(inst_cellmath__42_0_in2[15]), .B(inst_cellmath__42_0_in3[15]), .S0(N361));
MX2XL inst_cellmath__42_0_I72 (.Y(inst_cellmath__42_0_out0[18]), .A(inst_cellmath__42_0_in2[16]), .B(inst_cellmath__42_0_in3[16]), .S0(N361));
MX2XL inst_cellmath__42_0_I73 (.Y(inst_cellmath__42_0_out0[19]), .A(inst_cellmath__42_0_in2[17]), .B(inst_cellmath__42_0_in3[17]), .S0(N361));
MX2XL inst_cellmath__42_0_I74 (.Y(inst_cellmath__42_0_out0[20]), .A(inst_cellmath__42_0_in2[18]), .B(inst_cellmath__42_0_in3[18]), .S0(N361));
MX2XL inst_cellmath__42_0_I75 (.Y(inst_cellmath__42_0_out0[21]), .A(inst_cellmath__42_0_in2[19]), .B(inst_cellmath__42_0_in3[19]), .S0(N361));
MX2XL inst_cellmath__42_0_I76 (.Y(inst_cellmath__42_0_out0[22]), .A(inst_cellmath__42_0_in2[20]), .B(inst_cellmath__42_0_in3[20]), .S0(N361));
MX2XL inst_cellmath__42_0_I77 (.Y(inst_cellmath__42_0_out0[23]), .A(inst_cellmath__42_0_in2[21]), .B(inst_cellmath__42_0_in3[21]), .S0(N361));
MX2XL inst_cellmath__42_0_I78 (.Y(inst_cellmath__42_0_out0[24]), .A(inst_cellmath__42_0_in2[22]), .B(inst_cellmath__42_0_in3[22]), .S0(N361));
MX2XL inst_cellmath__42_0_I79 (.Y(inst_cellmath__42_0_out0[25]), .A(inst_cellmath__42_0_in2[23]), .B(inst_cellmath__42_0_in3[23]), .S0(N361));
MX2XL inst_cellmath__42_0_I80 (.Y(inst_cellmath__42_0_out0[26]), .A(inst_cellmath__42_0_in2[24]), .B(inst_cellmath__42_0_in3[24]), .S0(N361));
assign inst_cellmath__42_0_out0[0] = inst_cellmath__42_0_in0[0];
assign inst_cellmath__42_0_out0[1] = inst_cellmath__42_0_in1[0];
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__50_0_bdw410776230_bdw (
	inst_cellmath__50_0_out0,
	inst_cellmath__50_0_in0,
	inst_cellmath__50_0_in1
	); /* architecture "gate_level" */ 
output [1:0] inst_cellmath__50_0_out0;
input [0:0] inst_cellmath__50_0_in0,
	inst_cellmath__50_0_in1;
INVXL inst_cellmath__50_0_I19 (.Y(inst_cellmath__50_0_out0[0]), .A(inst_cellmath__50_0_in0[0]));
XOR2XL inst_cellmath__50_0_I17 (.Y(inst_cellmath__50_0_out0[1]), .A(inst_cellmath__50_0_in1[0]), .B(inst_cellmath__50_0_out0[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__43__56__bdw410776230_bdw (
	inst_cellmath__43__56__out0,
	inst_cellmath__43__56__in0,
	inst_cellmath__43__56__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__43__56__out0;
input [0:0] inst_cellmath__43__56__in0,
	inst_cellmath__43__56__in1;
OR2XL inst_cellmath__43__56__I0 (.Y(inst_cellmath__43__56__out0[0]), .A(inst_cellmath__43__56__in0[0]), .B(inst_cellmath__43__56__in1[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__43__55__bdw410776230_bdw (
	inst_cellmath__43__55__out0,
	inst_cellmath__43__55__in0,
	inst_cellmath__43__55__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__43__55__out0;
input [2:2] inst_cellmath__43__55__in0;
input [0:0] inst_cellmath__43__55__in1;
wire N16;
INVXL inst_cellmath__43__55__I4 (.Y(N16), .A(inst_cellmath__43__55__in0[2]));
AND2XL inst_cellmath__43__55__I1 (.Y(inst_cellmath__43__55__out0[0]), .A(N16), .B(inst_cellmath__43__55__in1[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__43_0_bdw410776230_bdw (
	inst_cellmath__43_0_out0,
	inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1,
	inst_cellmath__43_0_in2,
	inst_cellmath__43_0_in3
	); /* architecture "gate_level" */ 
output [26:0] inst_cellmath__43_0_out0;
input [1:0] inst_cellmath__43_0_in0;
input [24:0] inst_cellmath__43_0_in1,
	inst_cellmath__43_0_in2;
input [0:0] inst_cellmath__43_0_in3;
wire N361;
BUFX2 inst_cellmath__43_0_I90 (.Y(N361), .A(inst_cellmath__43_0_in3[0]));
MX2XL inst_cellmath__43_0_I56 (.Y(inst_cellmath__43_0_out0[2]), .A(inst_cellmath__43_0_in1[0]), .B(inst_cellmath__43_0_in2[0]), .S0(N361));
MX2XL inst_cellmath__43_0_I57 (.Y(inst_cellmath__43_0_out0[3]), .A(inst_cellmath__43_0_in1[1]), .B(inst_cellmath__43_0_in2[1]), .S0(N361));
MX2XL inst_cellmath__43_0_I58 (.Y(inst_cellmath__43_0_out0[4]), .A(inst_cellmath__43_0_in1[2]), .B(inst_cellmath__43_0_in2[2]), .S0(N361));
MX2XL inst_cellmath__43_0_I59 (.Y(inst_cellmath__43_0_out0[5]), .A(inst_cellmath__43_0_in1[3]), .B(inst_cellmath__43_0_in2[3]), .S0(N361));
MX2XL inst_cellmath__43_0_I60 (.Y(inst_cellmath__43_0_out0[6]), .A(inst_cellmath__43_0_in1[4]), .B(inst_cellmath__43_0_in2[4]), .S0(N361));
MX2XL inst_cellmath__43_0_I61 (.Y(inst_cellmath__43_0_out0[7]), .A(inst_cellmath__43_0_in1[5]), .B(inst_cellmath__43_0_in2[5]), .S0(N361));
MX2XL inst_cellmath__43_0_I62 (.Y(inst_cellmath__43_0_out0[8]), .A(inst_cellmath__43_0_in1[6]), .B(inst_cellmath__43_0_in2[6]), .S0(N361));
MX2XL inst_cellmath__43_0_I63 (.Y(inst_cellmath__43_0_out0[9]), .A(inst_cellmath__43_0_in1[7]), .B(inst_cellmath__43_0_in2[7]), .S0(N361));
MX2XL inst_cellmath__43_0_I64 (.Y(inst_cellmath__43_0_out0[10]), .A(inst_cellmath__43_0_in1[8]), .B(inst_cellmath__43_0_in2[8]), .S0(N361));
MX2XL inst_cellmath__43_0_I65 (.Y(inst_cellmath__43_0_out0[11]), .A(inst_cellmath__43_0_in1[9]), .B(inst_cellmath__43_0_in2[9]), .S0(N361));
MX2XL inst_cellmath__43_0_I66 (.Y(inst_cellmath__43_0_out0[12]), .A(inst_cellmath__43_0_in1[10]), .B(inst_cellmath__43_0_in2[10]), .S0(N361));
MX2XL inst_cellmath__43_0_I67 (.Y(inst_cellmath__43_0_out0[13]), .A(inst_cellmath__43_0_in1[11]), .B(inst_cellmath__43_0_in2[11]), .S0(N361));
MX2XL inst_cellmath__43_0_I68 (.Y(inst_cellmath__43_0_out0[14]), .A(inst_cellmath__43_0_in1[12]), .B(inst_cellmath__43_0_in2[12]), .S0(N361));
MX2XL inst_cellmath__43_0_I69 (.Y(inst_cellmath__43_0_out0[15]), .A(inst_cellmath__43_0_in1[13]), .B(inst_cellmath__43_0_in2[13]), .S0(N361));
MX2XL inst_cellmath__43_0_I70 (.Y(inst_cellmath__43_0_out0[16]), .A(inst_cellmath__43_0_in1[14]), .B(inst_cellmath__43_0_in2[14]), .S0(N361));
MX2XL inst_cellmath__43_0_I71 (.Y(inst_cellmath__43_0_out0[17]), .A(inst_cellmath__43_0_in1[15]), .B(inst_cellmath__43_0_in2[15]), .S0(N361));
MX2XL inst_cellmath__43_0_I72 (.Y(inst_cellmath__43_0_out0[18]), .A(inst_cellmath__43_0_in1[16]), .B(inst_cellmath__43_0_in2[16]), .S0(N361));
MX2XL inst_cellmath__43_0_I73 (.Y(inst_cellmath__43_0_out0[19]), .A(inst_cellmath__43_0_in1[17]), .B(inst_cellmath__43_0_in2[17]), .S0(N361));
MX2XL inst_cellmath__43_0_I74 (.Y(inst_cellmath__43_0_out0[20]), .A(inst_cellmath__43_0_in1[18]), .B(inst_cellmath__43_0_in2[18]), .S0(N361));
MX2XL inst_cellmath__43_0_I75 (.Y(inst_cellmath__43_0_out0[21]), .A(inst_cellmath__43_0_in1[19]), .B(inst_cellmath__43_0_in2[19]), .S0(N361));
MX2XL inst_cellmath__43_0_I76 (.Y(inst_cellmath__43_0_out0[22]), .A(inst_cellmath__43_0_in1[20]), .B(inst_cellmath__43_0_in2[20]), .S0(N361));
MX2XL inst_cellmath__43_0_I77 (.Y(inst_cellmath__43_0_out0[23]), .A(inst_cellmath__43_0_in1[21]), .B(inst_cellmath__43_0_in2[21]), .S0(N361));
MX2XL inst_cellmath__43_0_I78 (.Y(inst_cellmath__43_0_out0[24]), .A(inst_cellmath__43_0_in1[22]), .B(inst_cellmath__43_0_in2[22]), .S0(N361));
MX2XL inst_cellmath__43_0_I79 (.Y(inst_cellmath__43_0_out0[25]), .A(inst_cellmath__43_0_in1[23]), .B(inst_cellmath__43_0_in2[23]), .S0(N361));
MX2XL inst_cellmath__43_0_I80 (.Y(inst_cellmath__43_0_out0[26]), .A(inst_cellmath__43_0_in1[24]), .B(inst_cellmath__43_0_in2[24]), .S0(N361));
assign inst_cellmath__43_0_out0[0] = inst_cellmath__43_0_in0[0];
assign inst_cellmath__43_0_out0[1] = inst_cellmath__43_0_in0[1];
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__56_2mx_bdw410776230_bdw (
	inst_it2_cellmath__56_2mx_out0,
	inst_it2_cellmath__56_2mx_in0,
	inst_it2_cellmath__56_2mx_in1
	); /* architecture "gate_level" */ 
output [25:0] inst_it2_cellmath__56_2mx_out0;
input [2:2] inst_it2_cellmath__56_2mx_in0;
input [24:1] inst_it2_cellmath__56_2mx_in1;
wire N340;
INVXL inst_it2_cellmath__56_2mx_I92 (.Y(inst_it2_cellmath__56_2mx_out0[0]), .A(inst_it2_cellmath__56_2mx_in0[2]));
INVXL inst_it2_cellmath__56_2mx_I87 (.Y(N340), .A(inst_it2_cellmath__56_2mx_out0[0]));
XNOR2X1 inst_it2_cellmath__56_2mx_I29 (.Y(inst_it2_cellmath__56_2mx_out0[1]), .A(inst_it2_cellmath__56_2mx_in1[1]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I30 (.Y(inst_it2_cellmath__56_2mx_out0[2]), .A(inst_it2_cellmath__56_2mx_in1[2]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I31 (.Y(inst_it2_cellmath__56_2mx_out0[3]), .A(inst_it2_cellmath__56_2mx_in1[3]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I32 (.Y(inst_it2_cellmath__56_2mx_out0[4]), .A(inst_it2_cellmath__56_2mx_in1[4]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I33 (.Y(inst_it2_cellmath__56_2mx_out0[5]), .A(inst_it2_cellmath__56_2mx_in1[5]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I34 (.Y(inst_it2_cellmath__56_2mx_out0[6]), .A(inst_it2_cellmath__56_2mx_in1[6]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I35 (.Y(inst_it2_cellmath__56_2mx_out0[7]), .A(inst_it2_cellmath__56_2mx_in1[7]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I36 (.Y(inst_it2_cellmath__56_2mx_out0[8]), .A(inst_it2_cellmath__56_2mx_in1[8]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I37 (.Y(inst_it2_cellmath__56_2mx_out0[9]), .A(inst_it2_cellmath__56_2mx_in1[9]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I38 (.Y(inst_it2_cellmath__56_2mx_out0[10]), .A(inst_it2_cellmath__56_2mx_in1[10]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I39 (.Y(inst_it2_cellmath__56_2mx_out0[11]), .A(inst_it2_cellmath__56_2mx_in1[11]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I40 (.Y(inst_it2_cellmath__56_2mx_out0[12]), .A(inst_it2_cellmath__56_2mx_in1[12]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I41 (.Y(inst_it2_cellmath__56_2mx_out0[13]), .A(inst_it2_cellmath__56_2mx_in1[13]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I42 (.Y(inst_it2_cellmath__56_2mx_out0[14]), .A(inst_it2_cellmath__56_2mx_in1[14]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I43 (.Y(inst_it2_cellmath__56_2mx_out0[15]), .A(inst_it2_cellmath__56_2mx_in1[15]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I44 (.Y(inst_it2_cellmath__56_2mx_out0[16]), .A(inst_it2_cellmath__56_2mx_in1[16]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I45 (.Y(inst_it2_cellmath__56_2mx_out0[17]), .A(inst_it2_cellmath__56_2mx_in1[17]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I46 (.Y(inst_it2_cellmath__56_2mx_out0[18]), .A(inst_it2_cellmath__56_2mx_in1[18]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I47 (.Y(inst_it2_cellmath__56_2mx_out0[19]), .A(inst_it2_cellmath__56_2mx_in1[19]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I48 (.Y(inst_it2_cellmath__56_2mx_out0[20]), .A(inst_it2_cellmath__56_2mx_in1[20]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I49 (.Y(inst_it2_cellmath__56_2mx_out0[21]), .A(inst_it2_cellmath__56_2mx_in1[21]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I50 (.Y(inst_it2_cellmath__56_2mx_out0[22]), .A(inst_it2_cellmath__56_2mx_in1[22]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I51 (.Y(inst_it2_cellmath__56_2mx_out0[23]), .A(inst_it2_cellmath__56_2mx_in1[23]), .B(N340));
XNOR2X1 inst_it2_cellmath__56_2mx_I52 (.Y(inst_it2_cellmath__56_2mx_out0[24]), .A(inst_it2_cellmath__56_2mx_in1[24]), .B(N340));
assign inst_it2_cellmath__56_2mx_out0[25] = inst_it2_cellmath__56_2mx_out0[0];
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__57_2mx_bdw410776230_bdw (
	inst_it2_cellmath__57_2mx_out0,
	inst_it2_cellmath__57_2mx_in0,
	inst_it2_cellmath__57_2mx_in1
	); /* architecture "gate_level" */ 
output [25:0] inst_it2_cellmath__57_2mx_out0;
input [2:2] inst_it2_cellmath__57_2mx_in0;
input [25:2] inst_it2_cellmath__57_2mx_in1;
wire N271,N274;
INVXL buf1_A_I139 (.Y(N274), .A(inst_it2_cellmath__57_2mx_in0[2]));
INVXL buf1_A_I140 (.Y(N271), .A(N274));
INVXL inst_it2_cellmath__57_2mx_I111 (.Y(inst_it2_cellmath__57_2mx_out0[1]), .A(N271));
MXI2XL inst_it2_cellmath__57_2mx_I114 (.Y(inst_it2_cellmath__57_2mx_out0[2]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[2]));
MXI2XL inst_it2_cellmath__57_2mx_I115 (.Y(inst_it2_cellmath__57_2mx_out0[3]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[3]));
MXI2XL inst_it2_cellmath__57_2mx_I116 (.Y(inst_it2_cellmath__57_2mx_out0[4]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[4]));
MXI2XL inst_it2_cellmath__57_2mx_I117 (.Y(inst_it2_cellmath__57_2mx_out0[5]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[5]));
MXI2XL inst_it2_cellmath__57_2mx_I118 (.Y(inst_it2_cellmath__57_2mx_out0[6]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[6]));
MXI2XL inst_it2_cellmath__57_2mx_I119 (.Y(inst_it2_cellmath__57_2mx_out0[7]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[7]));
MXI2XL inst_it2_cellmath__57_2mx_I120 (.Y(inst_it2_cellmath__57_2mx_out0[8]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[8]));
MXI2XL inst_it2_cellmath__57_2mx_I121 (.Y(inst_it2_cellmath__57_2mx_out0[9]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[9]));
MXI2XL inst_it2_cellmath__57_2mx_I122 (.Y(inst_it2_cellmath__57_2mx_out0[10]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[10]));
MXI2XL inst_it2_cellmath__57_2mx_I123 (.Y(inst_it2_cellmath__57_2mx_out0[11]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[11]));
MXI2XL inst_it2_cellmath__57_2mx_I124 (.Y(inst_it2_cellmath__57_2mx_out0[12]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[12]));
MXI2XL inst_it2_cellmath__57_2mx_I125 (.Y(inst_it2_cellmath__57_2mx_out0[13]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[13]));
MXI2XL inst_it2_cellmath__57_2mx_I126 (.Y(inst_it2_cellmath__57_2mx_out0[14]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[14]));
MXI2XL inst_it2_cellmath__57_2mx_I127 (.Y(inst_it2_cellmath__57_2mx_out0[15]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[15]));
MXI2XL inst_it2_cellmath__57_2mx_I128 (.Y(inst_it2_cellmath__57_2mx_out0[16]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[16]));
MXI2XL inst_it2_cellmath__57_2mx_I129 (.Y(inst_it2_cellmath__57_2mx_out0[17]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[17]));
MXI2XL inst_it2_cellmath__57_2mx_I130 (.Y(inst_it2_cellmath__57_2mx_out0[18]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[18]));
MXI2XL inst_it2_cellmath__57_2mx_I131 (.Y(inst_it2_cellmath__57_2mx_out0[19]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[19]));
MXI2XL inst_it2_cellmath__57_2mx_I132 (.Y(inst_it2_cellmath__57_2mx_out0[20]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[20]));
MXI2XL inst_it2_cellmath__57_2mx_I133 (.Y(inst_it2_cellmath__57_2mx_out0[21]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[21]));
MXI2XL inst_it2_cellmath__57_2mx_I134 (.Y(inst_it2_cellmath__57_2mx_out0[22]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[22]));
MXI2XL inst_it2_cellmath__57_2mx_I135 (.Y(inst_it2_cellmath__57_2mx_out0[23]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[23]));
MXI2XL inst_it2_cellmath__57_2mx_I136 (.Y(inst_it2_cellmath__57_2mx_out0[24]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[24]));
MXI2XL inst_it2_cellmath__57_2mx_I137 (.Y(inst_it2_cellmath__57_2mx_out0[25]), .A(N271), .B(inst_it2_cellmath__57_2mx_out0[1]), .S0(inst_it2_cellmath__57_2mx_in1[25]));
assign inst_it2_cellmath__57_2mx_out0[0] = inst_it2_cellmath__57_2mx_out0[1];
endmodule

module cynw_cm_float_div_ieee_inst_fa_1820_10_bdw410776230_bdw (
	inst_fa_1820_10_out0,
	inst_fa_1820_10_out1,
	inst_fa_1820_10_in0,
	inst_fa_1820_10_in1,
	inst_fa_1820_10_in2,
	inst_fa_1820_10_in3
	); /* architecture "gate_level" */ 
output [25:0] inst_fa_1820_10_out0;
output [24:0] inst_fa_1820_10_out1;
input  inst_fa_1820_10_in0;
input [25:0] inst_fa_1820_10_in1;
input [23:0] inst_fa_1820_10_in2;
input [22:0] inst_fa_1820_10_in3;
ADDHX1 inst_fa_1820_10_I2 (.CO(inst_fa_1820_10_out1[2]), .S(inst_fa_1820_10_out0[2]), .A(inst_fa_1820_10_in2[0]), .B(inst_fa_1820_10_in1[2]));
ADDFX1 inst_fa_1820_10_I3 (.CO(inst_fa_1820_10_out1[3]), .S(inst_fa_1820_10_out0[3]), .A(inst_fa_1820_10_in2[1]), .B(inst_fa_1820_10_in3[0]), .CI(inst_fa_1820_10_in1[3]));
ADDFX1 inst_fa_1820_10_I4 (.CO(inst_fa_1820_10_out1[4]), .S(inst_fa_1820_10_out0[4]), .A(inst_fa_1820_10_in2[2]), .B(inst_fa_1820_10_in3[1]), .CI(inst_fa_1820_10_in1[4]));
ADDFX1 inst_fa_1820_10_I5 (.CO(inst_fa_1820_10_out1[5]), .S(inst_fa_1820_10_out0[5]), .A(inst_fa_1820_10_in2[3]), .B(inst_fa_1820_10_in3[2]), .CI(inst_fa_1820_10_in1[5]));
ADDFX1 inst_fa_1820_10_I6 (.CO(inst_fa_1820_10_out1[6]), .S(inst_fa_1820_10_out0[6]), .A(inst_fa_1820_10_in2[4]), .B(inst_fa_1820_10_in3[3]), .CI(inst_fa_1820_10_in1[6]));
ADDFX1 inst_fa_1820_10_I7 (.CO(inst_fa_1820_10_out1[7]), .S(inst_fa_1820_10_out0[7]), .A(inst_fa_1820_10_in2[5]), .B(inst_fa_1820_10_in3[4]), .CI(inst_fa_1820_10_in1[7]));
ADDFX1 inst_fa_1820_10_I8 (.CO(inst_fa_1820_10_out1[8]), .S(inst_fa_1820_10_out0[8]), .A(inst_fa_1820_10_in2[6]), .B(inst_fa_1820_10_in3[5]), .CI(inst_fa_1820_10_in1[8]));
ADDFX1 inst_fa_1820_10_I9 (.CO(inst_fa_1820_10_out1[9]), .S(inst_fa_1820_10_out0[9]), .A(inst_fa_1820_10_in2[7]), .B(inst_fa_1820_10_in3[6]), .CI(inst_fa_1820_10_in1[9]));
ADDFX1 inst_fa_1820_10_I10 (.CO(inst_fa_1820_10_out1[10]), .S(inst_fa_1820_10_out0[10]), .A(inst_fa_1820_10_in2[8]), .B(inst_fa_1820_10_in3[7]), .CI(inst_fa_1820_10_in1[10]));
ADDFX1 inst_fa_1820_10_I11 (.CO(inst_fa_1820_10_out1[11]), .S(inst_fa_1820_10_out0[11]), .A(inst_fa_1820_10_in2[9]), .B(inst_fa_1820_10_in3[8]), .CI(inst_fa_1820_10_in1[11]));
ADDFX1 inst_fa_1820_10_I12 (.CO(inst_fa_1820_10_out1[12]), .S(inst_fa_1820_10_out0[12]), .A(inst_fa_1820_10_in2[10]), .B(inst_fa_1820_10_in3[9]), .CI(inst_fa_1820_10_in1[12]));
ADDFX1 inst_fa_1820_10_I13 (.CO(inst_fa_1820_10_out1[13]), .S(inst_fa_1820_10_out0[13]), .A(inst_fa_1820_10_in2[11]), .B(inst_fa_1820_10_in3[10]), .CI(inst_fa_1820_10_in1[13]));
ADDFX1 inst_fa_1820_10_I14 (.CO(inst_fa_1820_10_out1[14]), .S(inst_fa_1820_10_out0[14]), .A(inst_fa_1820_10_in2[12]), .B(inst_fa_1820_10_in3[11]), .CI(inst_fa_1820_10_in1[14]));
ADDFX1 inst_fa_1820_10_I15 (.CO(inst_fa_1820_10_out1[15]), .S(inst_fa_1820_10_out0[15]), .A(inst_fa_1820_10_in2[13]), .B(inst_fa_1820_10_in3[12]), .CI(inst_fa_1820_10_in1[15]));
ADDFX1 inst_fa_1820_10_I16 (.CO(inst_fa_1820_10_out1[16]), .S(inst_fa_1820_10_out0[16]), .A(inst_fa_1820_10_in2[14]), .B(inst_fa_1820_10_in3[13]), .CI(inst_fa_1820_10_in1[16]));
ADDFX1 inst_fa_1820_10_I17 (.CO(inst_fa_1820_10_out1[17]), .S(inst_fa_1820_10_out0[17]), .A(inst_fa_1820_10_in2[15]), .B(inst_fa_1820_10_in3[14]), .CI(inst_fa_1820_10_in1[17]));
ADDFX1 inst_fa_1820_10_I18 (.CO(inst_fa_1820_10_out1[18]), .S(inst_fa_1820_10_out0[18]), .A(inst_fa_1820_10_in2[16]), .B(inst_fa_1820_10_in3[15]), .CI(inst_fa_1820_10_in1[18]));
ADDFX1 inst_fa_1820_10_I19 (.CO(inst_fa_1820_10_out1[19]), .S(inst_fa_1820_10_out0[19]), .A(inst_fa_1820_10_in2[17]), .B(inst_fa_1820_10_in3[16]), .CI(inst_fa_1820_10_in1[19]));
ADDFX1 inst_fa_1820_10_I20 (.CO(inst_fa_1820_10_out1[20]), .S(inst_fa_1820_10_out0[20]), .A(inst_fa_1820_10_in2[18]), .B(inst_fa_1820_10_in3[17]), .CI(inst_fa_1820_10_in1[20]));
ADDFX1 inst_fa_1820_10_I21 (.CO(inst_fa_1820_10_out1[21]), .S(inst_fa_1820_10_out0[21]), .A(inst_fa_1820_10_in2[19]), .B(inst_fa_1820_10_in3[18]), .CI(inst_fa_1820_10_in1[21]));
ADDFX1 inst_fa_1820_10_I22 (.CO(inst_fa_1820_10_out1[22]), .S(inst_fa_1820_10_out0[22]), .A(inst_fa_1820_10_in2[20]), .B(inst_fa_1820_10_in3[19]), .CI(inst_fa_1820_10_in1[22]));
ADDFX1 inst_fa_1820_10_I23 (.CO(inst_fa_1820_10_out1[23]), .S(inst_fa_1820_10_out0[23]), .A(inst_fa_1820_10_in2[21]), .B(inst_fa_1820_10_in3[20]), .CI(inst_fa_1820_10_in1[23]));
ADDFX1 inst_fa_1820_10_I24 (.CO(inst_fa_1820_10_out1[24]), .S(inst_fa_1820_10_out0[24]), .A(inst_fa_1820_10_in2[22]), .B(inst_fa_1820_10_in3[21]), .CI(inst_fa_1820_10_in1[24]));
XOR3XL inst_fa_1820_10_I115 (.Y(inst_fa_1820_10_out0[25]), .A(inst_fa_1820_10_in3[22]), .B(inst_fa_1820_10_in2[23]), .C(inst_fa_1820_10_in1[25]));
assign inst_fa_1820_10_out0[0] = inst_fa_1820_10_in1[0];
assign inst_fa_1820_10_out0[1] = inst_fa_1820_10_in1[1];
assign inst_fa_1820_10_out1[0] = inst_fa_1820_10_in0;
assign inst_fa_1820_10_out1[1] = 1'B0;
endmodule

module cynw_cm_float_div_ieee_inst_fa_1839_10_bdw410776230_bdw (
	inst_fa_1839_10_out0,
	inst_fa_1839_10_out1,
	inst_fa_1839_10_in0,
	inst_fa_1839_10_in1,
	inst_fa_1839_10_in2
	); /* architecture "gate_level" */ 
output [25:0] inst_fa_1839_10_out0;
output [24:0] inst_fa_1839_10_out1;
input [25:0] inst_fa_1839_10_in0;
input [24:0] inst_fa_1839_10_in1;
input [25:0] inst_fa_1839_10_in2;
wire N207;
ADDHX1 inst_fa_1839_10_I0 (.CO(inst_fa_1839_10_out1[0]), .S(inst_fa_1839_10_out0[0]), .A(inst_fa_1839_10_in0[0]), .B(inst_fa_1839_10_in2[0]));
ADDFX1 inst_fa_1839_10_I1 (.CO(inst_fa_1839_10_out1[1]), .S(inst_fa_1839_10_out0[1]), .A(inst_fa_1839_10_in1[0]), .B(inst_fa_1839_10_in0[1]), .CI(inst_fa_1839_10_in2[1]));
ADDFX1 inst_fa_1839_10_I2 (.CO(inst_fa_1839_10_out1[2]), .S(inst_fa_1839_10_out0[2]), .A(inst_fa_1839_10_in1[1]), .B(inst_fa_1839_10_in0[2]), .CI(inst_fa_1839_10_in2[2]));
ADDFX1 inst_fa_1839_10_I3 (.CO(inst_fa_1839_10_out1[3]), .S(inst_fa_1839_10_out0[3]), .A(inst_fa_1839_10_in1[2]), .B(inst_fa_1839_10_in0[3]), .CI(inst_fa_1839_10_in2[3]));
ADDFX1 inst_fa_1839_10_I4 (.CO(inst_fa_1839_10_out1[4]), .S(inst_fa_1839_10_out0[4]), .A(inst_fa_1839_10_in1[3]), .B(inst_fa_1839_10_in0[4]), .CI(inst_fa_1839_10_in2[4]));
ADDFX1 inst_fa_1839_10_I5 (.CO(inst_fa_1839_10_out1[5]), .S(inst_fa_1839_10_out0[5]), .A(inst_fa_1839_10_in1[4]), .B(inst_fa_1839_10_in0[5]), .CI(inst_fa_1839_10_in2[5]));
ADDFX1 inst_fa_1839_10_I6 (.CO(inst_fa_1839_10_out1[6]), .S(inst_fa_1839_10_out0[6]), .A(inst_fa_1839_10_in1[5]), .B(inst_fa_1839_10_in0[6]), .CI(inst_fa_1839_10_in2[6]));
ADDFX1 inst_fa_1839_10_I7 (.CO(inst_fa_1839_10_out1[7]), .S(inst_fa_1839_10_out0[7]), .A(inst_fa_1839_10_in1[6]), .B(inst_fa_1839_10_in0[7]), .CI(inst_fa_1839_10_in2[7]));
ADDFX1 inst_fa_1839_10_I8 (.CO(inst_fa_1839_10_out1[8]), .S(inst_fa_1839_10_out0[8]), .A(inst_fa_1839_10_in1[7]), .B(inst_fa_1839_10_in0[8]), .CI(inst_fa_1839_10_in2[8]));
ADDFX1 inst_fa_1839_10_I9 (.CO(inst_fa_1839_10_out1[9]), .S(inst_fa_1839_10_out0[9]), .A(inst_fa_1839_10_in1[8]), .B(inst_fa_1839_10_in0[9]), .CI(inst_fa_1839_10_in2[9]));
ADDFX1 inst_fa_1839_10_I10 (.CO(inst_fa_1839_10_out1[10]), .S(inst_fa_1839_10_out0[10]), .A(inst_fa_1839_10_in1[9]), .B(inst_fa_1839_10_in0[10]), .CI(inst_fa_1839_10_in2[10]));
ADDFX1 inst_fa_1839_10_I11 (.CO(inst_fa_1839_10_out1[11]), .S(inst_fa_1839_10_out0[11]), .A(inst_fa_1839_10_in1[10]), .B(inst_fa_1839_10_in0[11]), .CI(inst_fa_1839_10_in2[11]));
ADDFX1 inst_fa_1839_10_I12 (.CO(inst_fa_1839_10_out1[12]), .S(inst_fa_1839_10_out0[12]), .A(inst_fa_1839_10_in1[11]), .B(inst_fa_1839_10_in0[12]), .CI(inst_fa_1839_10_in2[12]));
ADDFX1 inst_fa_1839_10_I13 (.CO(inst_fa_1839_10_out1[13]), .S(inst_fa_1839_10_out0[13]), .A(inst_fa_1839_10_in1[12]), .B(inst_fa_1839_10_in0[13]), .CI(inst_fa_1839_10_in2[13]));
ADDFX1 inst_fa_1839_10_I14 (.CO(inst_fa_1839_10_out1[14]), .S(inst_fa_1839_10_out0[14]), .A(inst_fa_1839_10_in1[13]), .B(inst_fa_1839_10_in0[14]), .CI(inst_fa_1839_10_in2[14]));
ADDFX1 inst_fa_1839_10_I15 (.CO(inst_fa_1839_10_out1[15]), .S(inst_fa_1839_10_out0[15]), .A(inst_fa_1839_10_in1[14]), .B(inst_fa_1839_10_in0[15]), .CI(inst_fa_1839_10_in2[15]));
ADDFX1 inst_fa_1839_10_I16 (.CO(inst_fa_1839_10_out1[16]), .S(inst_fa_1839_10_out0[16]), .A(inst_fa_1839_10_in1[15]), .B(inst_fa_1839_10_in0[16]), .CI(inst_fa_1839_10_in2[16]));
ADDFX1 inst_fa_1839_10_I17 (.CO(inst_fa_1839_10_out1[17]), .S(inst_fa_1839_10_out0[17]), .A(inst_fa_1839_10_in1[16]), .B(inst_fa_1839_10_in0[17]), .CI(inst_fa_1839_10_in2[17]));
ADDFX1 inst_fa_1839_10_I18 (.CO(inst_fa_1839_10_out1[18]), .S(inst_fa_1839_10_out0[18]), .A(inst_fa_1839_10_in1[17]), .B(inst_fa_1839_10_in0[18]), .CI(inst_fa_1839_10_in2[18]));
ADDFX1 inst_fa_1839_10_I19 (.CO(inst_fa_1839_10_out1[19]), .S(inst_fa_1839_10_out0[19]), .A(inst_fa_1839_10_in1[18]), .B(inst_fa_1839_10_in0[19]), .CI(inst_fa_1839_10_in2[19]));
ADDFX1 inst_fa_1839_10_I20 (.CO(inst_fa_1839_10_out1[20]), .S(inst_fa_1839_10_out0[20]), .A(inst_fa_1839_10_in1[19]), .B(inst_fa_1839_10_in0[20]), .CI(inst_fa_1839_10_in2[20]));
ADDFX1 inst_fa_1839_10_I21 (.CO(inst_fa_1839_10_out1[21]), .S(inst_fa_1839_10_out0[21]), .A(inst_fa_1839_10_in1[20]), .B(inst_fa_1839_10_in0[21]), .CI(inst_fa_1839_10_in2[21]));
ADDFX1 inst_fa_1839_10_I22 (.CO(inst_fa_1839_10_out1[22]), .S(inst_fa_1839_10_out0[22]), .A(inst_fa_1839_10_in1[21]), .B(inst_fa_1839_10_in0[22]), .CI(inst_fa_1839_10_in2[22]));
ADDFX1 inst_fa_1839_10_I23 (.CO(inst_fa_1839_10_out1[23]), .S(inst_fa_1839_10_out0[23]), .A(inst_fa_1839_10_in1[22]), .B(inst_fa_1839_10_in0[23]), .CI(inst_fa_1839_10_in2[23]));
ADDFX1 inst_fa_1839_10_I24 (.CO(inst_fa_1839_10_out1[24]), .S(inst_fa_1839_10_out0[24]), .A(inst_fa_1839_10_in1[23]), .B(inst_fa_1839_10_in0[24]), .CI(inst_fa_1839_10_in2[24]));
ADDFX1 inst_fa_1839_10_I25 (.CO(N207), .S(inst_fa_1839_10_out0[25]), .A(inst_fa_1839_10_in1[24]), .B(inst_fa_1839_10_in0[25]), .CI(inst_fa_1839_10_in2[25]));
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__64__71__bdw410776230_bdw (
	inst_it2_cellmath__64__71__out0,
	inst_it2_cellmath__64__71__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_it2_cellmath__64__71__out0;
input [1:0] inst_it2_cellmath__64__71__in0;
NAND2XL inst_it2_cellmath__64__71__I0 (.Y(inst_it2_cellmath__64__71__out0[0]), .A(inst_it2_cellmath__64__71__in0[1]), .B(inst_it2_cellmath__64__71__in0[0]));
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__64__68__bdw410776230_bdw (
	inst_it2_cellmath__64__68__out0,
	inst_it2_cellmath__64__68__in0,
	inst_it2_cellmath__64__68__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_it2_cellmath__64__68__out0;
input [2:1] inst_it2_cellmath__64__68__in0;
input [0:0] inst_it2_cellmath__64__68__in1;
MX2XL inst_it2_cellmath__64__68__I2 (.Y(inst_it2_cellmath__64__68__out0[0]), .A(inst_it2_cellmath__64__68__in0[1]), .B(inst_it2_cellmath__64__68__in1[0]), .S0(inst_it2_cellmath__64__68__in0[2]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__40_0_bdw410776230_bdw (
	inst_cellmath__40_0_out0,
	inst_cellmath__40_0_in0,
	inst_cellmath__40_0_in1,
	inst_cellmath__40_0_in2,
	inst_cellmath__40_0_in3,
	inst_cellmath__40_0_in4
	); /* architecture "gate_level" */ 
output [28:0] inst_cellmath__40_0_out0;
input [0:0] inst_cellmath__40_0_in0,
	inst_cellmath__40_0_in1;
input  inst_cellmath__40_0_in2;
input [26:0] inst_cellmath__40_0_in3,
	inst_cellmath__40_0_in4;
wire N388;
BUFX2 inst_cellmath__40_0_I97 (.Y(N388), .A(inst_cellmath__40_0_in2));
MX2XL inst_cellmath__40_0_I60 (.Y(inst_cellmath__40_0_out0[2]), .A(inst_cellmath__40_0_in3[0]), .B(inst_cellmath__40_0_in4[0]), .S0(N388));
MX2XL inst_cellmath__40_0_I61 (.Y(inst_cellmath__40_0_out0[3]), .A(inst_cellmath__40_0_in3[1]), .B(inst_cellmath__40_0_in4[1]), .S0(N388));
MX2XL inst_cellmath__40_0_I62 (.Y(inst_cellmath__40_0_out0[4]), .A(inst_cellmath__40_0_in3[2]), .B(inst_cellmath__40_0_in4[2]), .S0(N388));
MX2XL inst_cellmath__40_0_I63 (.Y(inst_cellmath__40_0_out0[5]), .A(inst_cellmath__40_0_in3[3]), .B(inst_cellmath__40_0_in4[3]), .S0(N388));
MX2XL inst_cellmath__40_0_I64 (.Y(inst_cellmath__40_0_out0[6]), .A(inst_cellmath__40_0_in3[4]), .B(inst_cellmath__40_0_in4[4]), .S0(N388));
MX2XL inst_cellmath__40_0_I65 (.Y(inst_cellmath__40_0_out0[7]), .A(inst_cellmath__40_0_in3[5]), .B(inst_cellmath__40_0_in4[5]), .S0(N388));
MX2XL inst_cellmath__40_0_I66 (.Y(inst_cellmath__40_0_out0[8]), .A(inst_cellmath__40_0_in3[6]), .B(inst_cellmath__40_0_in4[6]), .S0(N388));
MX2XL inst_cellmath__40_0_I67 (.Y(inst_cellmath__40_0_out0[9]), .A(inst_cellmath__40_0_in3[7]), .B(inst_cellmath__40_0_in4[7]), .S0(N388));
MX2XL inst_cellmath__40_0_I68 (.Y(inst_cellmath__40_0_out0[10]), .A(inst_cellmath__40_0_in3[8]), .B(inst_cellmath__40_0_in4[8]), .S0(N388));
MX2XL inst_cellmath__40_0_I69 (.Y(inst_cellmath__40_0_out0[11]), .A(inst_cellmath__40_0_in3[9]), .B(inst_cellmath__40_0_in4[9]), .S0(N388));
MX2XL inst_cellmath__40_0_I70 (.Y(inst_cellmath__40_0_out0[12]), .A(inst_cellmath__40_0_in3[10]), .B(inst_cellmath__40_0_in4[10]), .S0(N388));
MX2XL inst_cellmath__40_0_I71 (.Y(inst_cellmath__40_0_out0[13]), .A(inst_cellmath__40_0_in3[11]), .B(inst_cellmath__40_0_in4[11]), .S0(N388));
MX2XL inst_cellmath__40_0_I72 (.Y(inst_cellmath__40_0_out0[14]), .A(inst_cellmath__40_0_in3[12]), .B(inst_cellmath__40_0_in4[12]), .S0(N388));
MX2XL inst_cellmath__40_0_I73 (.Y(inst_cellmath__40_0_out0[15]), .A(inst_cellmath__40_0_in3[13]), .B(inst_cellmath__40_0_in4[13]), .S0(N388));
MX2XL inst_cellmath__40_0_I74 (.Y(inst_cellmath__40_0_out0[16]), .A(inst_cellmath__40_0_in3[14]), .B(inst_cellmath__40_0_in4[14]), .S0(N388));
MX2XL inst_cellmath__40_0_I75 (.Y(inst_cellmath__40_0_out0[17]), .A(inst_cellmath__40_0_in3[15]), .B(inst_cellmath__40_0_in4[15]), .S0(N388));
MX2XL inst_cellmath__40_0_I76 (.Y(inst_cellmath__40_0_out0[18]), .A(inst_cellmath__40_0_in3[16]), .B(inst_cellmath__40_0_in4[16]), .S0(N388));
MX2XL inst_cellmath__40_0_I77 (.Y(inst_cellmath__40_0_out0[19]), .A(inst_cellmath__40_0_in3[17]), .B(inst_cellmath__40_0_in4[17]), .S0(N388));
MX2XL inst_cellmath__40_0_I78 (.Y(inst_cellmath__40_0_out0[20]), .A(inst_cellmath__40_0_in3[18]), .B(inst_cellmath__40_0_in4[18]), .S0(N388));
MX2XL inst_cellmath__40_0_I79 (.Y(inst_cellmath__40_0_out0[21]), .A(inst_cellmath__40_0_in3[19]), .B(inst_cellmath__40_0_in4[19]), .S0(N388));
MX2XL inst_cellmath__40_0_I80 (.Y(inst_cellmath__40_0_out0[22]), .A(inst_cellmath__40_0_in3[20]), .B(inst_cellmath__40_0_in4[20]), .S0(N388));
MX2XL inst_cellmath__40_0_I81 (.Y(inst_cellmath__40_0_out0[23]), .A(inst_cellmath__40_0_in3[21]), .B(inst_cellmath__40_0_in4[21]), .S0(N388));
MX2XL inst_cellmath__40_0_I82 (.Y(inst_cellmath__40_0_out0[24]), .A(inst_cellmath__40_0_in3[22]), .B(inst_cellmath__40_0_in4[22]), .S0(N388));
MX2XL inst_cellmath__40_0_I83 (.Y(inst_cellmath__40_0_out0[25]), .A(inst_cellmath__40_0_in3[23]), .B(inst_cellmath__40_0_in4[23]), .S0(N388));
MX2XL inst_cellmath__40_0_I84 (.Y(inst_cellmath__40_0_out0[26]), .A(inst_cellmath__40_0_in3[24]), .B(inst_cellmath__40_0_in4[24]), .S0(N388));
MX2XL inst_cellmath__40_0_I85 (.Y(inst_cellmath__40_0_out0[27]), .A(inst_cellmath__40_0_in3[25]), .B(inst_cellmath__40_0_in4[25]), .S0(N388));
MX2XL inst_cellmath__40_0_I86 (.Y(inst_cellmath__40_0_out0[28]), .A(inst_cellmath__40_0_in3[26]), .B(inst_cellmath__40_0_in4[26]), .S0(N388));
assign inst_cellmath__40_0_out0[0] = inst_cellmath__40_0_in0[0];
assign inst_cellmath__40_0_out0[1] = inst_cellmath__40_0_in1[0];
endmodule

module cynw_cm_float_div_ieee_inst_it2_cellmath__66_0_bdw410776230_bdw (
	inst_it2_cellmath__66_0_out0,
	inst_it2_cellmath__66_0_in0,
	inst_it2_cellmath__66_0_in1
	); /* architecture "gate_level" */ 
output [1:0] inst_it2_cellmath__66_0_out0;
input [0:0] inst_it2_cellmath__66_0_in0,
	inst_it2_cellmath__66_0_in1;
INVXL inst_it2_cellmath__66_0_I19 (.Y(inst_it2_cellmath__66_0_out0[0]), .A(inst_it2_cellmath__66_0_in0[0]));
XOR2XL inst_it2_cellmath__66_0_I17 (.Y(inst_it2_cellmath__66_0_out0[1]), .A(inst_it2_cellmath__66_0_in1[0]), .B(inst_it2_cellmath__66_0_out0[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__41__80__bdw410776230_bdw (
	inst_cellmath__41__80__out0,
	inst_cellmath__41__80__in0,
	inst_cellmath__41__80__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__41__80__out0;
input [0:0] inst_cellmath__41__80__in0,
	inst_cellmath__41__80__in1;
OR2XL inst_cellmath__41__80__I0 (.Y(inst_cellmath__41__80__out0[0]), .A(inst_cellmath__41__80__in0[0]), .B(inst_cellmath__41__80__in1[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__41__79__bdw410776230_bdw (
	inst_cellmath__41__79__out0,
	inst_cellmath__41__79__in0,
	inst_cellmath__41__79__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__41__79__out0;
input [2:2] inst_cellmath__41__79__in0;
input [0:0] inst_cellmath__41__79__in1;
wire N16;
INVXL inst_cellmath__41__79__I4 (.Y(N16), .A(inst_cellmath__41__79__in0[2]));
AND2XL inst_cellmath__41__79__I1 (.Y(inst_cellmath__41__79__out0[0]), .A(N16), .B(inst_cellmath__41__79__in1[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__41_0_bdw410776230_bdw (
	inst_cellmath__41_0_out0,
	inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3
	); /* architecture "gate_level" */ 
output [28:0] inst_cellmath__41_0_out0;
input [1:0] inst_cellmath__41_0_in0;
input [26:0] inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2;
input [0:0] inst_cellmath__41_0_in3;
wire N388;
BUFX2 inst_cellmath__41_0_I97 (.Y(N388), .A(inst_cellmath__41_0_in3[0]));
MX2XL inst_cellmath__41_0_I60 (.Y(inst_cellmath__41_0_out0[2]), .A(inst_cellmath__41_0_in1[0]), .B(inst_cellmath__41_0_in2[0]), .S0(N388));
MX2XL inst_cellmath__41_0_I61 (.Y(inst_cellmath__41_0_out0[3]), .A(inst_cellmath__41_0_in1[1]), .B(inst_cellmath__41_0_in2[1]), .S0(N388));
MX2XL inst_cellmath__41_0_I62 (.Y(inst_cellmath__41_0_out0[4]), .A(inst_cellmath__41_0_in1[2]), .B(inst_cellmath__41_0_in2[2]), .S0(N388));
MX2XL inst_cellmath__41_0_I63 (.Y(inst_cellmath__41_0_out0[5]), .A(inst_cellmath__41_0_in1[3]), .B(inst_cellmath__41_0_in2[3]), .S0(N388));
MX2XL inst_cellmath__41_0_I64 (.Y(inst_cellmath__41_0_out0[6]), .A(inst_cellmath__41_0_in1[4]), .B(inst_cellmath__41_0_in2[4]), .S0(N388));
MX2XL inst_cellmath__41_0_I65 (.Y(inst_cellmath__41_0_out0[7]), .A(inst_cellmath__41_0_in1[5]), .B(inst_cellmath__41_0_in2[5]), .S0(N388));
MX2XL inst_cellmath__41_0_I66 (.Y(inst_cellmath__41_0_out0[8]), .A(inst_cellmath__41_0_in1[6]), .B(inst_cellmath__41_0_in2[6]), .S0(N388));
MX2XL inst_cellmath__41_0_I67 (.Y(inst_cellmath__41_0_out0[9]), .A(inst_cellmath__41_0_in1[7]), .B(inst_cellmath__41_0_in2[7]), .S0(N388));
MX2XL inst_cellmath__41_0_I68 (.Y(inst_cellmath__41_0_out0[10]), .A(inst_cellmath__41_0_in1[8]), .B(inst_cellmath__41_0_in2[8]), .S0(N388));
MX2XL inst_cellmath__41_0_I69 (.Y(inst_cellmath__41_0_out0[11]), .A(inst_cellmath__41_0_in1[9]), .B(inst_cellmath__41_0_in2[9]), .S0(N388));
MX2XL inst_cellmath__41_0_I70 (.Y(inst_cellmath__41_0_out0[12]), .A(inst_cellmath__41_0_in1[10]), .B(inst_cellmath__41_0_in2[10]), .S0(N388));
MX2XL inst_cellmath__41_0_I71 (.Y(inst_cellmath__41_0_out0[13]), .A(inst_cellmath__41_0_in1[11]), .B(inst_cellmath__41_0_in2[11]), .S0(N388));
MX2XL inst_cellmath__41_0_I72 (.Y(inst_cellmath__41_0_out0[14]), .A(inst_cellmath__41_0_in1[12]), .B(inst_cellmath__41_0_in2[12]), .S0(N388));
MX2XL inst_cellmath__41_0_I73 (.Y(inst_cellmath__41_0_out0[15]), .A(inst_cellmath__41_0_in1[13]), .B(inst_cellmath__41_0_in2[13]), .S0(N388));
MX2XL inst_cellmath__41_0_I74 (.Y(inst_cellmath__41_0_out0[16]), .A(inst_cellmath__41_0_in1[14]), .B(inst_cellmath__41_0_in2[14]), .S0(N388));
MX2XL inst_cellmath__41_0_I75 (.Y(inst_cellmath__41_0_out0[17]), .A(inst_cellmath__41_0_in1[15]), .B(inst_cellmath__41_0_in2[15]), .S0(N388));
MX2XL inst_cellmath__41_0_I76 (.Y(inst_cellmath__41_0_out0[18]), .A(inst_cellmath__41_0_in1[16]), .B(inst_cellmath__41_0_in2[16]), .S0(N388));
MX2XL inst_cellmath__41_0_I77 (.Y(inst_cellmath__41_0_out0[19]), .A(inst_cellmath__41_0_in1[17]), .B(inst_cellmath__41_0_in2[17]), .S0(N388));
MX2XL inst_cellmath__41_0_I78 (.Y(inst_cellmath__41_0_out0[20]), .A(inst_cellmath__41_0_in1[18]), .B(inst_cellmath__41_0_in2[18]), .S0(N388));
MX2XL inst_cellmath__41_0_I79 (.Y(inst_cellmath__41_0_out0[21]), .A(inst_cellmath__41_0_in1[19]), .B(inst_cellmath__41_0_in2[19]), .S0(N388));
MX2XL inst_cellmath__41_0_I80 (.Y(inst_cellmath__41_0_out0[22]), .A(inst_cellmath__41_0_in1[20]), .B(inst_cellmath__41_0_in2[20]), .S0(N388));
MX2XL inst_cellmath__41_0_I81 (.Y(inst_cellmath__41_0_out0[23]), .A(inst_cellmath__41_0_in1[21]), .B(inst_cellmath__41_0_in2[21]), .S0(N388));
MX2XL inst_cellmath__41_0_I82 (.Y(inst_cellmath__41_0_out0[24]), .A(inst_cellmath__41_0_in1[22]), .B(inst_cellmath__41_0_in2[22]), .S0(N388));
MX2XL inst_cellmath__41_0_I83 (.Y(inst_cellmath__41_0_out0[25]), .A(inst_cellmath__41_0_in1[23]), .B(inst_cellmath__41_0_in2[23]), .S0(N388));
MX2XL inst_cellmath__41_0_I84 (.Y(inst_cellmath__41_0_out0[26]), .A(inst_cellmath__41_0_in1[24]), .B(inst_cellmath__41_0_in2[24]), .S0(N388));
MX2XL inst_cellmath__41_0_I85 (.Y(inst_cellmath__41_0_out0[27]), .A(inst_cellmath__41_0_in1[25]), .B(inst_cellmath__41_0_in2[25]), .S0(N388));
MX2XL inst_cellmath__41_0_I86 (.Y(inst_cellmath__41_0_out0[28]), .A(inst_cellmath__41_0_in1[26]), .B(inst_cellmath__41_0_in2[26]), .S0(N388));
assign inst_cellmath__41_0_out0[0] = inst_cellmath__41_0_in0[0];
assign inst_cellmath__41_0_out0[1] = inst_cellmath__41_0_in0[1];
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__67_0_bdw410776230_bdw (
	inst_cellmath__67_0_out0,
	inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__67_0_out0;
input [30:23] inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1;
wire N64,N66,N68,N70,N72,N74,N76 
	,N95,N99,N100,N103,N104,N107,N108,N111 
	,N112,N115,N116,N119,N122,N126,N128,N130 
	,N132,N134,N136,N138;
INVXL inst_cellmath__67_0_I18 (.Y(N64), .A(inst_cellmath__67_0_in0[23]));
INVXL inst_cellmath__67_0_I19 (.Y(N66), .A(inst_cellmath__67_0_in0[24]));
INVXL inst_cellmath__67_0_I20 (.Y(N68), .A(inst_cellmath__67_0_in0[25]));
INVXL inst_cellmath__67_0_I21 (.Y(N70), .A(inst_cellmath__67_0_in0[26]));
INVXL inst_cellmath__67_0_I22 (.Y(N72), .A(inst_cellmath__67_0_in0[27]));
INVXL inst_cellmath__67_0_I23 (.Y(N74), .A(inst_cellmath__67_0_in0[28]));
INVXL inst_cellmath__67_0_I24 (.Y(N76), .A(inst_cellmath__67_0_in0[29]));
INVXL inst_cellmath__67_0_I39 (.Y(N95), .A(inst_cellmath__67_0_in1[24]));
XNOR2X1 hap1_A_I54 (.Y(N99), .A(inst_cellmath__67_0_in1[24]), .B(N68));
OR2XL hap1_A_I55 (.Y(N100), .A(inst_cellmath__67_0_in1[24]), .B(N68));
XNOR2X1 hap1_A_I56 (.Y(N103), .A(inst_cellmath__67_0_in1[26]), .B(N70));
OR2XL hap1_A_I57 (.Y(N104), .A(inst_cellmath__67_0_in1[26]), .B(N70));
XNOR2X1 hap1_A_I58 (.Y(N107), .A(inst_cellmath__67_0_in1[27]), .B(N72));
OR2XL hap1_A_I59 (.Y(N108), .A(inst_cellmath__67_0_in1[27]), .B(N72));
XNOR2X1 hap1_A_I60 (.Y(N111), .A(inst_cellmath__67_0_in1[28]), .B(N74));
OR2XL hap1_A_I61 (.Y(N112), .A(inst_cellmath__67_0_in1[28]), .B(N74));
XNOR2X1 hap1_A_I62 (.Y(N115), .A(inst_cellmath__67_0_in1[29]), .B(N76));
OR2XL hap1_A_I63 (.Y(N116), .A(inst_cellmath__67_0_in1[29]), .B(N76));
XNOR2X1 inst_cellmath__67_0_I45 (.Y(N119), .A(inst_cellmath__67_0_in1[30]), .B(inst_cellmath__67_0_in0[30]));
XNOR2X1 hap1_A_I64 (.Y(inst_cellmath__67_0_out0[0]), .A(N64), .B(inst_cellmath__67_0_in1[23]));
OR2XL hap1_A_I65 (.Y(N122), .A(N64), .B(inst_cellmath__67_0_in1[23]));
ADDFX1 inst_cellmath__67_0_I47 (.CO(N126), .S(inst_cellmath__67_0_out0[1]), .A(N95), .B(N66), .CI(N122));
ADDFX1 inst_cellmath__67_0_I48 (.CO(N128), .S(inst_cellmath__67_0_out0[2]), .A(N99), .B(inst_cellmath__67_0_in1[25]), .CI(N126));
ADDFX1 inst_cellmath__67_0_I49 (.CO(N130), .S(inst_cellmath__67_0_out0[3]), .A(N103), .B(N100), .CI(N128));
ADDFX1 inst_cellmath__67_0_I50 (.CO(N132), .S(inst_cellmath__67_0_out0[4]), .A(N107), .B(N104), .CI(N130));
ADDFX1 inst_cellmath__67_0_I51 (.CO(N134), .S(inst_cellmath__67_0_out0[5]), .A(N111), .B(N108), .CI(N132));
ADDFX1 inst_cellmath__67_0_I52 (.CO(N136), .S(inst_cellmath__67_0_out0[6]), .A(N115), .B(N112), .CI(N134));
ADDFX1 inst_cellmath__67_0_I53 (.CO(N138), .S(inst_cellmath__67_0_out0[7]), .A(N119), .B(N116), .CI(N136));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__68_0_bdw410776230_bdw (
	inst_cellmath__68_0_out0,
	inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__68_0_out0;
input [30:23] inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1;
wire N66,N68,N70,N72,N74,N76,N78 
	,N80,N98,N103,N107,N109,N111,N113,N115 
	,N117,N119;
INVXL inst_cellmath__68_0_I18 (.Y(N66), .A(inst_cellmath__68_0_in0[23]));
INVXL inst_cellmath__68_0_I19 (.Y(N68), .A(inst_cellmath__68_0_in0[24]));
INVXL inst_cellmath__68_0_I20 (.Y(N70), .A(inst_cellmath__68_0_in0[25]));
INVXL inst_cellmath__68_0_I21 (.Y(N72), .A(inst_cellmath__68_0_in0[26]));
INVXL inst_cellmath__68_0_I22 (.Y(N74), .A(inst_cellmath__68_0_in0[27]));
INVXL inst_cellmath__68_0_I23 (.Y(N76), .A(inst_cellmath__68_0_in0[28]));
INVXL inst_cellmath__68_0_I24 (.Y(N78), .A(inst_cellmath__68_0_in0[29]));
INVXL inst_cellmath__68_0_I25 (.Y(N80), .A(inst_cellmath__68_0_in0[30]));
INVXL inst_cellmath__68_0_I40 (.Y(N98), .A(inst_cellmath__68_0_in1[30]));
ADDHX1 inst_cellmath__68_0_I41 (.CO(N103), .S(inst_cellmath__68_0_out0[0]), .A(inst_cellmath__68_0_in1[23]), .B(N66));
ADDFX1 inst_cellmath__68_0_I42 (.CO(N107), .S(inst_cellmath__68_0_out0[1]), .A(N68), .B(inst_cellmath__68_0_in1[24]), .CI(N103));
ADDFX1 inst_cellmath__68_0_I43 (.CO(N109), .S(inst_cellmath__68_0_out0[2]), .A(N70), .B(inst_cellmath__68_0_in1[25]), .CI(N107));
ADDFX1 inst_cellmath__68_0_I44 (.CO(N111), .S(inst_cellmath__68_0_out0[3]), .A(N72), .B(inst_cellmath__68_0_in1[26]), .CI(N109));
ADDFX1 inst_cellmath__68_0_I45 (.CO(N113), .S(inst_cellmath__68_0_out0[4]), .A(N74), .B(inst_cellmath__68_0_in1[27]), .CI(N111));
ADDFX1 inst_cellmath__68_0_I46 (.CO(N115), .S(inst_cellmath__68_0_out0[5]), .A(N76), .B(inst_cellmath__68_0_in1[28]), .CI(N113));
ADDFX1 inst_cellmath__68_0_I47 (.CO(N117), .S(inst_cellmath__68_0_out0[6]), .A(N78), .B(inst_cellmath__68_0_in1[29]), .CI(N115));
ADDFX1 inst_cellmath__68_0_I48 (.CO(N119), .S(inst_cellmath__68_0_out0[7]), .A(N80), .B(N98), .CI(N117));
XNOR2X1 hap1_A_I52 (.Y(inst_cellmath__68_0_out0[8]), .A(inst_cellmath__68_0_in1[30]), .B(N119));
NOR2XL hap1_A_I53 (.Y(inst_cellmath__68_0_out0[9]), .A(inst_cellmath__68_0_in1[30]), .B(N119));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__69__82__bdw410776230_bdw (
	inst_cellmath__69__82__out0,
	inst_cellmath__69__82__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__69__82__out0;
input [7:0] inst_cellmath__69__82__in0;
wire N11,N17,N19;
AND2XL inst_cellmath__69__82__I0 (.Y(N11), .A(inst_cellmath__69__82__in0[0]), .B(inst_cellmath__69__82__in0[1]));
NAND3XL inst_cellmath__69__82__I15 (.Y(N17), .A(inst_cellmath__69__82__in0[3]), .B(inst_cellmath__69__82__in0[4]), .C(inst_cellmath__69__82__in0[7]));
NAND4X1 inst_cellmath__69__82__I16 (.Y(N19), .A(inst_cellmath__69__82__in0[2]), .B(N11), .C(inst_cellmath__69__82__in0[6]), .D(inst_cellmath__69__82__in0[5]));
NOR2X6 inst_cellmath__69__82__I9 (.Y(inst_cellmath__69__82__out0[0]), .A(N17), .B(N19));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__69__81__bdw410776230_bdw (
	inst_cellmath__69__81__out0,
	inst_cellmath__69__81__in0,
	inst_cellmath__69__81__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__69__81__out0;
input [0:0] inst_cellmath__69__81__in0;
input [8:8] inst_cellmath__69__81__in1;
OR2XL inst_cellmath__69__81__I0 (.Y(inst_cellmath__69__81__out0[0]), .A(inst_cellmath__69__81__in1[8]), .B(inst_cellmath__69__81__in0[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__69_0_bdw410776230_bdw (
	inst_cellmath__69_0_out0,
	inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__69_0_out0;
input [0:0] inst_cellmath__69_0_in0;
input [9:9] inst_cellmath__69_0_in1;
NOR2BX1 inst_cellmath__69_0_I3 (.Y(inst_cellmath__69_0_out0), .AN(inst_cellmath__69_0_in0[0]), .B(inst_cellmath__69_0_in1[9]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__70__83__bdw410776230_bdw (
	inst_cellmath__70__83__out0,
	inst_cellmath__70__83__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__70__83__out0;
input [8:0] inst_cellmath__70__83__in0;
wire N12,N13,N16,N20,N53,N54,N55 
	;
NOR2XL inst_cellmath__70__83__I0 (.Y(N12), .A(inst_cellmath__70__83__in0[0]), .B(inst_cellmath__70__83__in0[1]));
NOR2XL inst_cellmath__70__83__I1 (.Y(N13), .A(inst_cellmath__70__83__in0[2]), .B(inst_cellmath__70__83__in0[3]));
NOR2XL inst_cellmath__70__83__I4 (.Y(N16), .A(inst_cellmath__70__83__in0[6]), .B(inst_cellmath__70__83__in0[7]));
INVXL inst_cellmath__70__83__I20 (.Y(N53), .A(inst_cellmath__70__83__in0[8]));
INVXL inst_cellmath__70__83__I21 (.Y(N54), .A(inst_cellmath__70__83__in0[4]));
INVXL inst_cellmath__70__83__I22 (.Y(N55), .A(inst_cellmath__70__83__in0[5]));
AND4XL inst_cellmath__70__83__I31 (.Y(N20), .A(N53), .B(N54), .C(N55), .D(N12));
NAND3XL inst_cellmath__70__83__I29 (.Y(inst_cellmath__70__83__out0[0]), .A(N13), .B(N16), .C(N20));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__70_0_bdw410776230_bdw (
	inst_cellmath__70_0_out0,
	inst_cellmath__70_0_in0,
	inst_cellmath__70_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__70_0_out0;
input [0:0] inst_cellmath__70_0_in0;
input [9:9] inst_cellmath__70_0_in1;
NAND2BXL inst_cellmath__70_0_I2 (.Y(inst_cellmath__70_0_out0), .AN(inst_cellmath__70_0_in1[9]), .B(inst_cellmath__70_0_in0[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__71_0_bdw410776230_bdw (
	inst_cellmath__71_0_out0,
	inst_cellmath__71_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__71_0_out0;
input [9:0] inst_cellmath__71_0_in0;
wire N15,N16,N17,N22,N23;
NAND3BXL inst_cellmath__71_0_I64 (.Y(N15), .AN(inst_cellmath__71_0_in0[9]), .B(inst_cellmath__71_0_in0[0]), .C(inst_cellmath__71_0_in0[1]));
NAND2XL inst_cellmath__71_0_I3 (.Y(N16), .A(inst_cellmath__71_0_in0[2]), .B(inst_cellmath__71_0_in0[3]));
NAND2XL inst_cellmath__71_0_I4 (.Y(N17), .A(inst_cellmath__71_0_in0[4]), .B(inst_cellmath__71_0_in0[6]));
NOR2XL inst_cellmath__71_0_I9 (.Y(N22), .A(N16), .B(N17));
NAND3BXL inst_cellmath__71_0_I66 (.Y(N23), .AN(inst_cellmath__71_0_in0[8]), .B(inst_cellmath__71_0_in0[7]), .C(N22));
NOR3BXL inst_cellmath__71_0_I67 (.Y(inst_cellmath__71_0_out0), .AN(inst_cellmath__71_0_in0[5]), .B(N15), .C(N23));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__72_0_bdw410776230_bdw (
	inst_cellmath__72_0_out0,
	inst_cellmath__72_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__72_0_out0;
input [8:0] inst_cellmath__72_0_in0;
wire N14,N15,N21,N64,N65;
NOR2XL inst_cellmath__72_0_I2 (.Y(N14), .A(inst_cellmath__72_0_in0[2]), .B(inst_cellmath__72_0_in0[3]));
NOR2XL inst_cellmath__72_0_I3 (.Y(N15), .A(inst_cellmath__72_0_in0[4]), .B(inst_cellmath__72_0_in0[6]));
INVXL inst_cellmath__72_0_I22 (.Y(N64), .A(inst_cellmath__72_0_in0[7]));
INVXL inst_cellmath__72_0_I23 (.Y(N65), .A(inst_cellmath__72_0_in0[8]));
NAND4XL inst_cellmath__72_0_I33 (.Y(N21), .A(N64), .B(N65), .C(N14), .D(N15));
NOR4BX1 inst_cellmath__72_0_I67 (.Y(inst_cellmath__72_0_out0), .AN(inst_cellmath__72_0_in0[0]), .B(inst_cellmath__72_0_in0[1]), .C(inst_cellmath__72_0_in0[5]), .D(N21));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__73_0_bdw410776230_bdw (
	inst_cellmath__73_0_out0,
	inst_cellmath__73_0_in0,
	inst_cellmath__73_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__73_0_out0;
input  inst_cellmath__73_0_in0,
	inst_cellmath__73_0_in1;
NOR2BX1 inst_cellmath__73_0_I3 (.Y(inst_cellmath__73_0_out0), .AN(inst_cellmath__73_0_in1), .B(inst_cellmath__73_0_in0));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__74_0_bdw410776230_bdw (
	inst_cellmath__74_0_out0,
	inst_cellmath__74_0_in0,
	inst_cellmath__74_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__74_0_out0;
input  inst_cellmath__74_0_in0,
	inst_cellmath__74_0_in1;
OR2XL inst_cellmath__74_0_I0 (.Y(inst_cellmath__74_0_out0), .A(inst_cellmath__74_0_in0), .B(inst_cellmath__74_0_in1));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__75_0_bdw410776230_bdw (
	inst_cellmath__75_0_out0,
	inst_cellmath__75_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__75_0_out0;
input [30:23] inst_cellmath__75_0_in0;
wire N11,N12,N13,N14;
NAND2XL inst_cellmath__75_0_I0 (.Y(N11), .A(inst_cellmath__75_0_in0[30]), .B(inst_cellmath__75_0_in0[24]));
NAND2XL inst_cellmath__75_0_I1 (.Y(N12), .A(inst_cellmath__75_0_in0[29]), .B(inst_cellmath__75_0_in0[25]));
NAND2XL inst_cellmath__75_0_I2 (.Y(N13), .A(inst_cellmath__75_0_in0[27]), .B(inst_cellmath__75_0_in0[28]));
NAND2XL inst_cellmath__75_0_I3 (.Y(N14), .A(inst_cellmath__75_0_in0[26]), .B(inst_cellmath__75_0_in0[23]));
NOR4X1 inst_cellmath__75_0_I25 (.Y(inst_cellmath__75_0_out0), .A(N12), .B(N11), .C(N13), .D(N14));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__76_0_bdw410776230_bdw (
	inst_cellmath__76_0_out0,
	inst_cellmath__76_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__76_0_out0;
input [30:23] inst_cellmath__76_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__76_0_I0 (.Y(N11), .A(inst_cellmath__76_0_in0[25]), .B(inst_cellmath__76_0_in0[27]));
NAND2XL inst_cellmath__76_0_I1 (.Y(N12), .A(inst_cellmath__76_0_in0[28]), .B(inst_cellmath__76_0_in0[23]));
NAND2XL inst_cellmath__76_0_I2 (.Y(N13), .A(inst_cellmath__76_0_in0[29]), .B(inst_cellmath__76_0_in0[24]));
NAND2XL inst_cellmath__76_0_I3 (.Y(N14), .A(inst_cellmath__76_0_in0[30]), .B(inst_cellmath__76_0_in0[26]));
NOR2XL inst_cellmath__76_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__76_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__76_0_I6 (.Y(inst_cellmath__76_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__77_0_bdw410776230_bdw (
	inst_cellmath__77_0_out0,
	inst_cellmath__77_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__77_0_out0;
input [22:0] inst_cellmath__77_0_in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N40,N45,N47,N48 
	,N73,N167;
NOR2XL inst_cellmath__77_0_I0 (.Y(N26), .A(inst_cellmath__77_0_in0[1]), .B(inst_cellmath__77_0_in0[2]));
NOR2XL inst_cellmath__77_0_I1 (.Y(N27), .A(inst_cellmath__77_0_in0[18]), .B(inst_cellmath__77_0_in0[16]));
NOR2XL inst_cellmath__77_0_I2 (.Y(N28), .A(inst_cellmath__77_0_in0[14]), .B(inst_cellmath__77_0_in0[12]));
NOR2XL inst_cellmath__77_0_I3 (.Y(N29), .A(inst_cellmath__77_0_in0[10]), .B(inst_cellmath__77_0_in0[8]));
NOR2XL inst_cellmath__77_0_I4 (.Y(N30), .A(inst_cellmath__77_0_in0[6]), .B(inst_cellmath__77_0_in0[4]));
NOR2XL inst_cellmath__77_0_I5 (.Y(N31), .A(inst_cellmath__77_0_in0[19]), .B(inst_cellmath__77_0_in0[17]));
NOR2XL inst_cellmath__77_0_I6 (.Y(N32), .A(inst_cellmath__77_0_in0[15]), .B(inst_cellmath__77_0_in0[13]));
NOR2XL inst_cellmath__77_0_I7 (.Y(N33), .A(inst_cellmath__77_0_in0[11]), .B(inst_cellmath__77_0_in0[9]));
NOR2XL inst_cellmath__77_0_I8 (.Y(N34), .A(inst_cellmath__77_0_in0[7]), .B(inst_cellmath__77_0_in0[5]));
NOR2XL inst_cellmath__77_0_I9 (.Y(N35), .A(inst_cellmath__77_0_in0[3]), .B(inst_cellmath__77_0_in0[0]));
NOR2XL inst_cellmath__77_0_I10 (.Y(N36), .A(inst_cellmath__77_0_in0[22]), .B(inst_cellmath__77_0_in0[21]));
NAND2XL inst_cellmath__77_0_I14 (.Y(N40), .A(N29), .B(N30));
AND4XL inst_cellmath__77_0_I35 (.Y(N45), .A(N32), .B(N34), .C(N33), .D(N31));
NAND3XL hyperpropagate_4_1_A_I78 (.Y(N167), .A(N26), .B(N35), .C(N36));
NOR2XL hyperpropagate_4_1_A_I79 (.Y(N48), .A(inst_cellmath__77_0_in0[20]), .B(N167));
NAND3XL hyperpropagate_4_1_A_I39 (.Y(N73), .A(N27), .B(N28), .C(N45));
NOR2XL hyperpropagate_4_1_A_I40 (.Y(N47), .A(N40), .B(N73));
NAND2XL inst_cellmath__77_0_I23 (.Y(inst_cellmath__77_0_out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__78_0_bdw410776230_bdw (
	inst_cellmath__78_0_out0,
	inst_cellmath__78_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__78_0_out0;
input [22:0] inst_cellmath__78_0_in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N40,N45,N47,N48 
	,N113,N207;
NOR2XL inst_cellmath__78_0_I0 (.Y(N26), .A(inst_cellmath__78_0_in0[1]), .B(inst_cellmath__78_0_in0[2]));
NOR2XL inst_cellmath__78_0_I1 (.Y(N27), .A(inst_cellmath__78_0_in0[18]), .B(inst_cellmath__78_0_in0[16]));
NOR2XL inst_cellmath__78_0_I2 (.Y(N28), .A(inst_cellmath__78_0_in0[14]), .B(inst_cellmath__78_0_in0[12]));
NOR2XL inst_cellmath__78_0_I3 (.Y(N29), .A(inst_cellmath__78_0_in0[10]), .B(inst_cellmath__78_0_in0[8]));
NOR2XL inst_cellmath__78_0_I4 (.Y(N30), .A(inst_cellmath__78_0_in0[6]), .B(inst_cellmath__78_0_in0[4]));
NOR2XL inst_cellmath__78_0_I5 (.Y(N31), .A(inst_cellmath__78_0_in0[19]), .B(inst_cellmath__78_0_in0[17]));
NOR2XL inst_cellmath__78_0_I6 (.Y(N32), .A(inst_cellmath__78_0_in0[15]), .B(inst_cellmath__78_0_in0[13]));
NOR2XL inst_cellmath__78_0_I7 (.Y(N33), .A(inst_cellmath__78_0_in0[11]), .B(inst_cellmath__78_0_in0[9]));
NOR2XL inst_cellmath__78_0_I8 (.Y(N34), .A(inst_cellmath__78_0_in0[7]), .B(inst_cellmath__78_0_in0[5]));
NOR2XL inst_cellmath__78_0_I9 (.Y(N35), .A(inst_cellmath__78_0_in0[3]), .B(inst_cellmath__78_0_in0[0]));
NOR2XL inst_cellmath__78_0_I10 (.Y(N36), .A(inst_cellmath__78_0_in0[20]), .B(inst_cellmath__78_0_in0[22]));
NAND2XL inst_cellmath__78_0_I14 (.Y(N40), .A(N29), .B(N30));
AND4XL inst_cellmath__78_0_I56 (.Y(N45), .A(N32), .B(N34), .C(N33), .D(N31));
NAND3XL hyperpropagate_4_1_A_I99 (.Y(N207), .A(N35), .B(N26), .C(N36));
NOR2XL hyperpropagate_4_1_A_I100 (.Y(N48), .A(inst_cellmath__78_0_in0[21]), .B(N207));
NAND3XL hyperpropagate_4_1_A_I60 (.Y(N113), .A(N27), .B(N28), .C(N45));
NOR2XL hyperpropagate_4_1_A_I61 (.Y(N47), .A(N40), .B(N113));
NAND2XL inst_cellmath__78_0_I23 (.Y(inst_cellmath__78_0_out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__79_1_bdw410776230_bdw (
	inst_cellmath__79_1_out0,
	inst_cellmath__79_1_in0,
	inst_cellmath__79_1_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__79_1_out0;
input  inst_cellmath__79_1_in0,
	inst_cellmath__79_1_in1;
AND2XL inst_cellmath__79_1_I0 (.Y(inst_cellmath__79_1_out0), .A(inst_cellmath__79_1_in1), .B(inst_cellmath__79_1_in0));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__80_0_bdw410776230_bdw (
	inst_cellmath__80_0_out0,
	inst_cellmath__80_0_in0,
	inst_cellmath__80_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__80_0_out0;
input  inst_cellmath__80_0_in0,
	inst_cellmath__80_0_in1;
AND2XL inst_cellmath__80_0_I0 (.Y(inst_cellmath__80_0_out0), .A(inst_cellmath__80_0_in1), .B(inst_cellmath__80_0_in0));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__83_0_bdw410776230_bdw (
	inst_cellmath__83_0_out0,
	inst_cellmath__83_0_in0,
	inst_cellmath__83_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__83_0_out0;
input  inst_cellmath__83_0_in0,
	inst_cellmath__83_0_in1;
NOR2BX1 inst_cellmath__83_0_I2 (.Y(inst_cellmath__83_0_out0), .AN(inst_cellmath__83_0_in1), .B(inst_cellmath__83_0_in0));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__84_0_bdw410776230_bdw (
	inst_cellmath__84_0_out0,
	inst_cellmath__84_0_in0,
	inst_cellmath__84_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__84_0_out0;
input  inst_cellmath__84_0_in0,
	inst_cellmath__84_0_in1;
NOR2BX1 inst_cellmath__84_0_I2 (.Y(inst_cellmath__84_0_out0), .AN(inst_cellmath__84_0_in1), .B(inst_cellmath__84_0_in0));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__85__85__bdw410776230_bdw (
	inst_cellmath__85__85__out0,
	inst_cellmath__85__85__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__85__85__out0;
input [30:23] inst_cellmath__85__85__in0;
wire N11,N12,N13,N14;
NOR2XL inst_cellmath__85__85__I0 (.Y(N11), .A(inst_cellmath__85__85__in0[30]), .B(inst_cellmath__85__85__in0[24]));
NOR2XL inst_cellmath__85__85__I1 (.Y(N12), .A(inst_cellmath__85__85__in0[29]), .B(inst_cellmath__85__85__in0[25]));
NOR2XL inst_cellmath__85__85__I2 (.Y(N13), .A(inst_cellmath__85__85__in0[27]), .B(inst_cellmath__85__85__in0[28]));
NOR2XL inst_cellmath__85__85__I3 (.Y(N14), .A(inst_cellmath__85__85__in0[26]), .B(inst_cellmath__85__85__in0[23]));
AND4XL inst_cellmath__85__85__I16 (.Y(inst_cellmath__85__85__out0), .A(N11), .B(N12), .C(N13), .D(N14));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__86__86__bdw410776230_bdw (
	inst_cellmath__86__86__out0,
	inst_cellmath__86__86__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__86__86__out0;
input [30:23] inst_cellmath__86__86__in0;
wire N11,N12,N13,N14;
NOR2XL inst_cellmath__86__86__I0 (.Y(N11), .A(inst_cellmath__86__86__in0[25]), .B(inst_cellmath__86__86__in0[27]));
NOR2XL inst_cellmath__86__86__I1 (.Y(N12), .A(inst_cellmath__86__86__in0[28]), .B(inst_cellmath__86__86__in0[23]));
NOR2XL inst_cellmath__86__86__I2 (.Y(N13), .A(inst_cellmath__86__86__in0[29]), .B(inst_cellmath__86__86__in0[24]));
NOR2XL inst_cellmath__86__86__I3 (.Y(N14), .A(inst_cellmath__86__86__in0[30]), .B(inst_cellmath__86__86__in0[26]));
AND4XL inst_cellmath__86__86__I16 (.Y(inst_cellmath__86__86__out0), .A(N11), .B(N13), .C(N12), .D(N14));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__87__87__bdw410776230_bdw (
	inst_cellmath__87__87__out0,
	inst_cellmath__87__87__in0,
	inst_cellmath__87__87__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__87__87__out0;
input  inst_cellmath__87__87__in0,
	inst_cellmath__87__87__in1;
AND2XL inst_cellmath__87__87__I0 (.Y(inst_cellmath__87__87__out0[0]), .A(inst_cellmath__87__87__in1), .B(inst_cellmath__87__87__in0));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__87__88__bdw410776230_bdw (
	inst_cellmath__87__88__out0,
	inst_cellmath__87__88__in0,
	inst_cellmath__87__88__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__87__88__out0;
input  inst_cellmath__87__88__in0,
	inst_cellmath__87__88__in1;
AND2XL inst_cellmath__87__88__I0 (.Y(inst_cellmath__87__88__out0[0]), .A(inst_cellmath__87__88__in0), .B(inst_cellmath__87__88__in1));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__87_0_bdw410776230_bdw (
	inst_cellmath__87_0_out0,
	inst_cellmath__87_0_in0,
	inst_cellmath__87_0_in1,
	inst_cellmath__87_0_in2,
	inst_cellmath__87_0_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__87_0_out0;
input [0:0] inst_cellmath__87_0_in0,
	inst_cellmath__87_0_in1;
input  inst_cellmath__87_0_in2,
	inst_cellmath__87_0_in3;
OR4X1 inst_cellmath__87_0_I6 (.Y(inst_cellmath__87_0_out0), .A(inst_cellmath__87_0_in0[0]), .B(inst_cellmath__87_0_in3), .C(inst_cellmath__87_0_in2), .D(inst_cellmath__87_0_in1[0]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__88_0_bdw410776230_bdw (
	inst_cellmath__88_0_out0,
	inst_cellmath__88_0_in0,
	inst_cellmath__88_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__88_0_out0;
input  inst_cellmath__88_0_in0,
	inst_cellmath__88_0_in1;
OR2XL inst_cellmath__88_0_I0 (.Y(inst_cellmath__88_0_out0), .A(inst_cellmath__88_0_in0), .B(inst_cellmath__88_0_in1));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__89_0_bdw410776230_bdw (
	inst_cellmath__89_0_out0,
	inst_cellmath__89_0_in0,
	inst_cellmath__89_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__89_0_out0;
input  inst_cellmath__89_0_in0,
	inst_cellmath__89_0_in1;
OR2XL inst_cellmath__89_0_I0 (.Y(inst_cellmath__89_0_out0), .A(inst_cellmath__89_0_in0), .B(inst_cellmath__89_0_in1));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__91_0_bdw410776230_bdw (
	inst_cellmath__91_0_out0,
	inst_cellmath__91_0_in0,
	inst_cellmath__91_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__91_0_out0;
input [31:31] inst_cellmath__91_0_in0,
	inst_cellmath__91_0_in1;
XOR2XL inst_cellmath__91_0_I0 (.Y(inst_cellmath__91_0_out0), .A(inst_cellmath__91_0_in0[31]), .B(inst_cellmath__91_0_in1[31]));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__92__95__bdw410776230_bdw (
	inst_cellmath__92__95__out0,
	inst_cellmath__92__95__in0,
	inst_cellmath__92__95__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__92__95__out0;
input  inst_cellmath__92__95__in0,
	inst_cellmath__92__95__in1;
OR2XL inst_cellmath__92__95__I0 (.Y(inst_cellmath__92__95__out0[0]), .A(inst_cellmath__92__95__in0), .B(inst_cellmath__92__95__in1));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__90_2WWMM_bdw410776230_bdw (
	inst_cellmath__90_2WWMM_out0,
	inst_cellmath__90_2WWMM_in0,
	inst_cellmath__90_2WWMM_in1,
	inst_cellmath__90_2WWMM_in2,
	inst_cellmath__90_2WWMM_in3,
	inst_cellmath__90_2WWMM_in4,
	inst_cellmath__90_2WWMM_in5,
	inst_cellmath__90_2WWMM_in6
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__90_2WWMM_out0;
input [31:31] inst_cellmath__90_2WWMM_in0;
input [21:0] inst_cellmath__90_2WWMM_in1;
input [0:0] inst_cellmath__90_2WWMM_in2;
input [31:31] inst_cellmath__90_2WWMM_in3;
input [21:0] inst_cellmath__90_2WWMM_in4;
input  inst_cellmath__90_2WWMM_in5,
	inst_cellmath__90_2WWMM_in6;
wire N124,N128,N246;
NOR2BX1 inst_cellmath__90_2WWMM_I132 (.Y(N246), .AN(inst_cellmath__90_2WWMM_in5), .B(inst_cellmath__90_2WWMM_in6));
NOR2XL inst_cellmath__90_2WWMM_I2 (.Y(N124), .A(inst_cellmath__90_2WWMM_in5), .B(inst_cellmath__90_2WWMM_in6));
AOI22XL inst_cellmath__90_2WWMM_I6 (.Y(N128), .A0(inst_cellmath__90_2WWMM_in3[31]), .A1(inst_cellmath__90_2WWMM_in6), .B0(N246), .B1(inst_cellmath__90_2WWMM_in0[31]));
AO22XL inst_cellmath__90_2WWMM_I7 (.Y(inst_cellmath__90_2WWMM_out0[1]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[0]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[0]));
AO22XL inst_cellmath__90_2WWMM_I8 (.Y(inst_cellmath__90_2WWMM_out0[2]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[1]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[1]));
AO22XL inst_cellmath__90_2WWMM_I9 (.Y(inst_cellmath__90_2WWMM_out0[3]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[2]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[2]));
AO22XL inst_cellmath__90_2WWMM_I10 (.Y(inst_cellmath__90_2WWMM_out0[4]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[3]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[3]));
AO22XL inst_cellmath__90_2WWMM_I11 (.Y(inst_cellmath__90_2WWMM_out0[5]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[4]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[4]));
AO22XL inst_cellmath__90_2WWMM_I12 (.Y(inst_cellmath__90_2WWMM_out0[6]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[5]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[5]));
AO22XL inst_cellmath__90_2WWMM_I13 (.Y(inst_cellmath__90_2WWMM_out0[7]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[6]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[6]));
AO22XL inst_cellmath__90_2WWMM_I14 (.Y(inst_cellmath__90_2WWMM_out0[8]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[7]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[7]));
AO22XL inst_cellmath__90_2WWMM_I15 (.Y(inst_cellmath__90_2WWMM_out0[9]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[8]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[8]));
AO22XL inst_cellmath__90_2WWMM_I16 (.Y(inst_cellmath__90_2WWMM_out0[10]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[9]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[9]));
AO22XL inst_cellmath__90_2WWMM_I17 (.Y(inst_cellmath__90_2WWMM_out0[11]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[10]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[10]));
AO22XL inst_cellmath__90_2WWMM_I18 (.Y(inst_cellmath__90_2WWMM_out0[12]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[11]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[11]));
AO22XL inst_cellmath__90_2WWMM_I19 (.Y(inst_cellmath__90_2WWMM_out0[13]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[12]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[12]));
AO22XL inst_cellmath__90_2WWMM_I20 (.Y(inst_cellmath__90_2WWMM_out0[14]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[13]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[13]));
AO22XL inst_cellmath__90_2WWMM_I21 (.Y(inst_cellmath__90_2WWMM_out0[15]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[14]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[14]));
AO22XL inst_cellmath__90_2WWMM_I22 (.Y(inst_cellmath__90_2WWMM_out0[16]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[15]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[15]));
AO22XL inst_cellmath__90_2WWMM_I23 (.Y(inst_cellmath__90_2WWMM_out0[17]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[16]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[16]));
AO22XL inst_cellmath__90_2WWMM_I24 (.Y(inst_cellmath__90_2WWMM_out0[18]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[17]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[17]));
AO22XL inst_cellmath__90_2WWMM_I25 (.Y(inst_cellmath__90_2WWMM_out0[19]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[18]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[18]));
AO22XL inst_cellmath__90_2WWMM_I26 (.Y(inst_cellmath__90_2WWMM_out0[20]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[19]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[19]));
AO22XL inst_cellmath__90_2WWMM_I27 (.Y(inst_cellmath__90_2WWMM_out0[21]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[20]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[20]));
AO22XL inst_cellmath__90_2WWMM_I28 (.Y(inst_cellmath__90_2WWMM_out0[22]), .A0(inst_cellmath__90_2WWMM_in6), .A1(inst_cellmath__90_2WWMM_in4[21]), .B0(N246), .B1(inst_cellmath__90_2WWMM_in1[21]));
OAI2BB1X1 inst_cellmath__90_2WWMM_I133 (.Y(inst_cellmath__90_2WWMM_out0[0]), .A0N(N124), .A1N(inst_cellmath__90_2WWMM_in2[0]), .B0(N128));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__96_0_bdw410776230_bdw (
	inst_cellmath__96_0_out0,
	inst_cellmath__96_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__96_0_out0;
input [3:0] inst_cellmath__96_0_in0;
wire N43,N45;
INVXL inst_cellmath__96_0_I22 (.Y(N43), .A(inst_cellmath__96_0_in0[3]));
NAND4XL inst_cellmath__96_0_I23 (.Y(N45), .A(inst_cellmath__96_0_in0[0]), .B(inst_cellmath__96_0_in0[1]), .C(inst_cellmath__96_0_in0[2]), .D(N43));
INVXL inst_cellmath__96_0_I24 (.Y(inst_cellmath__96_0_out0), .A(N45));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__133__109__bdw410776230_bdw (
	inst_cellmath__133__109__out0,
	inst_cellmath__133__109__in0,
	inst_cellmath__133__109__in1,
	inst_cellmath__133__109__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__133__109__out0;
input  inst_cellmath__133__109__in0,
	inst_cellmath__133__109__in1,
	inst_cellmath__133__109__in2;
OR3XL inst_cellmath__133__109__I3 (.Y(inst_cellmath__133__109__out0[0]), .A(inst_cellmath__133__109__in0), .B(inst_cellmath__133__109__in1), .C(inst_cellmath__133__109__in2));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__135_0_bdw410776230_bdw (
	inst_cellmath__135_0_out0,
	inst_cellmath__135_0_in0,
	inst_cellmath__135_0_in1,
	inst_cellmath__135_0_in2,
	inst_cellmath__135_0_in3,
	inst_cellmath__135_0_in4
	); /* architecture "gate_level" */ 
output  inst_cellmath__135_0_out0;
input  inst_cellmath__135_0_in0,
	inst_cellmath__135_0_in1,
	inst_cellmath__135_0_in2,
	inst_cellmath__135_0_in3,
	inst_cellmath__135_0_in4;
wire N11,N12,N33;
NOR2XL inst_cellmath__135_0_I1 (.Y(N12), .A(inst_cellmath__135_0_in1), .B(inst_cellmath__135_0_in3));
INVXL inst_cellmath__135_0_I10 (.Y(N33), .A(inst_cellmath__135_0_in4));
NOR3BXL inst_cellmath__135_0_I12 (.Y(N11), .AN(N33), .B(inst_cellmath__135_0_in0), .C(inst_cellmath__135_0_in2));
NAND2X6 inst_cellmath__135_0_I5 (.Y(inst_cellmath__135_0_out0), .A(N12), .B(N11));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__136_0_bdw410776230_bdw (
	inst_cellmath__136_0_out0,
	inst_cellmath__136_0_in0,
	inst_cellmath__136_0_in1,
	inst_cellmath__136_0_in2,
	inst_cellmath__136_0_in3,
	inst_cellmath__136_0_in4
	); /* architecture "gate_level" */ 
output  inst_cellmath__136_0_out0;
input  inst_cellmath__136_0_in0,
	inst_cellmath__136_0_in1,
	inst_cellmath__136_0_in2,
	inst_cellmath__136_0_in3,
	inst_cellmath__136_0_in4;
wire N8,N11,N12,N33,N34,N35;
NOR2XL inst_cellmath__136_0_I0 (.Y(N8), .A(inst_cellmath__136_0_in1), .B(inst_cellmath__136_0_in0));
INVXL inst_cellmath__136_0_I10 (.Y(N33), .A(inst_cellmath__136_0_in2));
INVXL inst_cellmath__136_0_I11 (.Y(N34), .A(inst_cellmath__136_0_in3));
NAND2XL inst_cellmath__136_0_I1 (.Y(N12), .A(N33), .B(N34));
INVXL inst_cellmath__136_0_I12 (.Y(N35), .A(inst_cellmath__136_0_in4));
NAND2XL inst_cellmath__136_0_I3 (.Y(N11), .A(N35), .B(N8));
OR2XL inst_cellmath__136_0_I5 (.Y(inst_cellmath__136_0_out0), .A(N12), .B(N11));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__137_2_bdw410776230_bdw (
	inst_cellmath__137_2_out0,
	inst_cellmath__137_2_in0,
	inst_cellmath__137_2_in1,
	inst_cellmath__137_2_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__137_2_out0;
input  inst_cellmath__137_2_in0,
	inst_cellmath__137_2_in1,
	inst_cellmath__137_2_in2;
MX2XL inst_cellmath__137_2_I2 (.Y(inst_cellmath__137_2_out0), .A(inst_cellmath__137_2_in1), .B(inst_cellmath__137_2_in0), .S0(inst_cellmath__137_2_in2));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__113__113__bdw410776230_bdw (
	inst_cellmath__113__113__out0,
	inst_cellmath__113__113__in0,
	inst_cellmath__113__113__in1,
	inst_cellmath__113__113__in2,
	inst_cellmath__113__113__in3,
	inst_cellmath__113__113__in4
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__113__113__out0;
input  inst_cellmath__113__113__in0;
input [0:0] inst_cellmath__113__113__in1;
input  inst_cellmath__113__113__in2;
input [7:0] inst_cellmath__113__113__in3,
	inst_cellmath__113__113__in4;
wire N37,N39,N41,N43,N45,N47,N49 
	,N51,N80,N82,N92;
NOR2XL inst_cellmath__113__113__I0 (.Y(N80), .A(inst_cellmath__113__113__in2), .B(inst_cellmath__113__113__in0));
NOR2BX1 inst_cellmath__113__113__I43 (.Y(N82), .AN(inst_cellmath__113__113__in2), .B(inst_cellmath__113__113__in0));
AOI22XL inst_cellmath__113__113__I6 (.Y(N37), .A0(inst_cellmath__113__113__in4[0]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[0]));
AOI22XL inst_cellmath__113__113__I7 (.Y(N39), .A0(inst_cellmath__113__113__in4[1]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[1]));
AOI22XL inst_cellmath__113__113__I8 (.Y(N41), .A0(inst_cellmath__113__113__in4[2]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[2]));
AOI22XL inst_cellmath__113__113__I9 (.Y(N43), .A0(inst_cellmath__113__113__in4[3]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[3]));
AOI22XL inst_cellmath__113__113__I10 (.Y(N45), .A0(inst_cellmath__113__113__in4[4]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[4]));
AOI22XL inst_cellmath__113__113__I11 (.Y(N47), .A0(inst_cellmath__113__113__in4[5]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[5]));
AOI22XL inst_cellmath__113__113__I12 (.Y(N49), .A0(inst_cellmath__113__113__in4[6]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[6]));
AOI22XL inst_cellmath__113__113__I13 (.Y(N51), .A0(inst_cellmath__113__113__in4[7]), .A1(N82), .B0(N80), .B1(inst_cellmath__113__113__in3[7]));
NAND2XL inst_cellmath__113__113__I47 (.Y(N92), .A(inst_cellmath__113__113__in0), .B(inst_cellmath__113__113__in1[0]));
NAND2XL inst_cellmath__113__113__I25 (.Y(inst_cellmath__113__113__out0[0]), .A(N92), .B(N37));
NAND2XL inst_cellmath__113__113__I26 (.Y(inst_cellmath__113__113__out0[1]), .A(N92), .B(N39));
NAND2XL inst_cellmath__113__113__I27 (.Y(inst_cellmath__113__113__out0[2]), .A(N92), .B(N41));
NAND2XL inst_cellmath__113__113__I28 (.Y(inst_cellmath__113__113__out0[3]), .A(N92), .B(N43));
NAND2XL inst_cellmath__113__113__I29 (.Y(inst_cellmath__113__113__out0[4]), .A(N92), .B(N45));
NAND2XL inst_cellmath__113__113__I30 (.Y(inst_cellmath__113__113__out0[5]), .A(N92), .B(N47));
NAND2XL inst_cellmath__113__113__I31 (.Y(inst_cellmath__113__113__out0[6]), .A(N92), .B(N49));
NAND2XL inst_cellmath__113__113__I32 (.Y(inst_cellmath__113__113__out0[7]), .A(N92), .B(N51));
endmodule

module cynw_cm_float_div_ieee_inst_cellmath__113__115__U_2WWMM_bdw410776230_bdw (
	inst_cellmath__113__115__U_2WWMM_out0,
	inst_cellmath__113__115__U_2WWMM_in0,
	inst_cellmath__113__115__U_2WWMM_in1,
	inst_cellmath__113__115__U_2WWMM_in2,
	inst_cellmath__113__115__U_2WWMM_in3,
	inst_cellmath__113__115__U_2WWMM_in4
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__113__115__U_2WWMM_out0;
input  inst_cellmath__113__115__U_2WWMM_in0;
input [22:1] inst_cellmath__113__115__U_2WWMM_in1;
input [0:0] inst_cellmath__113__115__U_2WWMM_in2;
input [21:0] inst_cellmath__113__115__U_2WWMM_in3;
input  inst_cellmath__113__115__U_2WWMM_in4;
wire N298,N299;
AND2XL inst_cellmath__113__115__U_2WWMM_I119 (.Y(N298), .A(inst_cellmath__113__115__U_2WWMM_in4), .B(inst_cellmath__113__115__U_2WWMM_in0));
INVXL inst_cellmath__113__115__U_2WWMM_I57 (.Y(N299), .A(inst_cellmath__113__115__U_2WWMM_in0));
AO22XL inst_cellmath__113__115__U_2WWMM_I7 (.Y(inst_cellmath__113__115__U_2WWMM_out0[0]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[0]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in2[0]));
AO22XL inst_cellmath__113__115__U_2WWMM_I8 (.Y(inst_cellmath__113__115__U_2WWMM_out0[1]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[1]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[1]));
AO22XL inst_cellmath__113__115__U_2WWMM_I9 (.Y(inst_cellmath__113__115__U_2WWMM_out0[2]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[2]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[2]));
AO22XL inst_cellmath__113__115__U_2WWMM_I10 (.Y(inst_cellmath__113__115__U_2WWMM_out0[3]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[3]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[3]));
AO22XL inst_cellmath__113__115__U_2WWMM_I11 (.Y(inst_cellmath__113__115__U_2WWMM_out0[4]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[4]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[4]));
AO22XL inst_cellmath__113__115__U_2WWMM_I12 (.Y(inst_cellmath__113__115__U_2WWMM_out0[5]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[5]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[5]));
AO22XL inst_cellmath__113__115__U_2WWMM_I13 (.Y(inst_cellmath__113__115__U_2WWMM_out0[6]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[6]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[6]));
AO22XL inst_cellmath__113__115__U_2WWMM_I14 (.Y(inst_cellmath__113__115__U_2WWMM_out0[7]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[7]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[7]));
AO22XL inst_cellmath__113__115__U_2WWMM_I15 (.Y(inst_cellmath__113__115__U_2WWMM_out0[8]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[8]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[8]));
AO22XL inst_cellmath__113__115__U_2WWMM_I16 (.Y(inst_cellmath__113__115__U_2WWMM_out0[9]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[9]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[9]));
AO22XL inst_cellmath__113__115__U_2WWMM_I17 (.Y(inst_cellmath__113__115__U_2WWMM_out0[10]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[10]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[10]));
AO22XL inst_cellmath__113__115__U_2WWMM_I18 (.Y(inst_cellmath__113__115__U_2WWMM_out0[11]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[11]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[11]));
AO22XL inst_cellmath__113__115__U_2WWMM_I19 (.Y(inst_cellmath__113__115__U_2WWMM_out0[12]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[12]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[12]));
AO22XL inst_cellmath__113__115__U_2WWMM_I20 (.Y(inst_cellmath__113__115__U_2WWMM_out0[13]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[13]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[13]));
AO22XL inst_cellmath__113__115__U_2WWMM_I21 (.Y(inst_cellmath__113__115__U_2WWMM_out0[14]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[14]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[14]));
AO22XL inst_cellmath__113__115__U_2WWMM_I22 (.Y(inst_cellmath__113__115__U_2WWMM_out0[15]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[15]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[15]));
AO22XL inst_cellmath__113__115__U_2WWMM_I23 (.Y(inst_cellmath__113__115__U_2WWMM_out0[16]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[16]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[16]));
AO22XL inst_cellmath__113__115__U_2WWMM_I24 (.Y(inst_cellmath__113__115__U_2WWMM_out0[17]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[17]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[17]));
AO22XL inst_cellmath__113__115__U_2WWMM_I25 (.Y(inst_cellmath__113__115__U_2WWMM_out0[18]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[18]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[18]));
AO22XL inst_cellmath__113__115__U_2WWMM_I26 (.Y(inst_cellmath__113__115__U_2WWMM_out0[19]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[19]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[19]));
AO22XL inst_cellmath__113__115__U_2WWMM_I27 (.Y(inst_cellmath__113__115__U_2WWMM_out0[20]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[20]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[20]));
AO22XL inst_cellmath__113__115__U_2WWMM_I28 (.Y(inst_cellmath__113__115__U_2WWMM_out0[21]), .A0(N298), .A1(inst_cellmath__113__115__U_2WWMM_in3[21]), .B0(N299), .B1(inst_cellmath__113__115__U_2WWMM_in1[21]));
AO21XL inst_cellmath__113__115__U_2WWMM_I61 (.Y(inst_cellmath__113__115__U_2WWMM_out0[22]), .A0(N299), .A1(inst_cellmath__113__115__U_2WWMM_in1[22]), .B0(N298));
endmodule

/* CADENCE  uLLyQwzZqxw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




