/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:30 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_mul_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x;
wire  DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__33;
wire [9:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34;
wire  DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__41,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__42;
wire [47:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43;
wire [7:0] DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54;
wire  DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__60,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__61,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N267,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N268,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N269,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N270,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N272,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N273,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N274,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N276,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1314,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1318,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1338,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1340,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1361,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1369,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1372,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1374,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1378,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1380,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1383,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1389,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1393,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1425,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1429,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1451,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1483,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1485,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1489,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1491,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1494,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1500,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1504,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1551,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1552,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1553,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1554,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1555,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1556,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1557,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1558,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1559,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1561,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1563,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1564,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1566,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1567,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1569,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1570,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1571,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1572,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1574,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1576,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1577,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1578,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1579,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1580,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1581,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1582,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1583,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1584,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1585,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1586,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1587,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1588,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1589,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1590,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1591,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1592,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1593,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1594,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1595,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1596,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1597,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1600,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1601,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1602,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1603,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1604,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1605,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1606,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1607,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1608,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1609,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1610,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1611,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1612,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1613,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1614,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1616,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1617,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1618,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1619,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1620,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1622,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1624,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1625,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1626,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1627,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1628,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1631,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1632,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1633,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1634,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1636,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1637,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1638,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1639,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1640,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1641,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1642,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1643,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1644,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1645,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1646,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1647,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1648,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1650,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1651,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1652,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1654,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1655,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1656,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1657,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1659,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1660,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1661,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1662,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1664,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1665,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1666,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1667,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1668,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1669,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1670,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1671,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1673,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1674,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1675,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1676,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1677,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1678,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1679,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1680,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1681,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1683,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1684,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1685,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1686,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1687,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1690,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1691,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1692,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1693,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1694,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1696,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1698,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1699,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1700,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1701,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1703,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1704,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1705,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1707,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1708,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1709,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1710,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1711,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1712,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1713,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1714,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1715,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1716,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1717,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1718,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1719,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1720,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1721,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1722,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1723,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1725,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1727,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1728,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1729,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1730,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1731,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1733,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1734,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1735,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1736,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1737,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1738,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1739,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1740,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1741,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1742,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1743,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1744,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1745,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1746,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1747,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1748,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1750,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1751,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1752,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1753,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1754,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1755,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1757,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1759,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1760,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1761,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1762,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1763,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1764,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1766,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1767,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1769,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1771,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1773,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1774,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1775,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1776,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1779,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1780,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1781,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1782,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1783,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1784,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1785,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1786,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1787,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1788,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1791,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1792,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1793,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1796,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1799,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1800,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1801,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1802,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1804,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1805,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1806,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1807,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1808,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1809,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1810,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1811,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1812,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1813,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1815,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1816,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1817,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1818,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1819,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1821,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1822,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1824,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1825,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1826,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1827,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1828,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1830,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1832,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1834,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1835,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1837,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1838,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1839,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1840,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1841,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1842,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1843,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1844,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1845,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1847,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1848,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1849,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1852,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1853,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1855,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1856,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1858,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1859,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1860,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1861,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1862,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1863,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1864,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1865,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1866,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1867,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1869,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1870,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1872,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1873,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1874,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1875,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1876,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1877,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1878,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1879,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1880,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1881,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1882,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1883,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1884,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1885,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1886,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1887,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1888,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1889,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1890,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1891,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1892,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1893,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1894,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1896,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1897,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1899,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1900,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1903,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1905,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1906,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1907,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1908,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1909,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1910,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1911,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1912,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1913,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1914,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1915,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1916,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1918,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1919,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1920,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1921,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1922,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1924,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1925,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1926,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1927,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1929,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1930,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1932,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1934,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1935,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1936,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1938,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1939,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1940,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1942,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1944,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1946,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1947,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1949,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1950,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1951,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1952,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1953,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1954,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1956,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1957,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1958,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1959,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1960,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1961,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1962,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1963,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1964,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1965,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1966,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1967,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1968,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1969,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1972,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1973,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1974,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1975,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1976,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1977,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1978,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1979,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1980,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1981,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1982,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1983,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1984,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1985,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1986,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1987,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1988,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1990,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1991,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1993,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1994,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1995,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1996,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1997,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1998,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1999,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2000,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2001,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2003,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2004,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2005,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2007,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2008,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2009,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2010,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2011,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2012,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2013,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2014,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2015,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2016,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2017,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2018,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2019,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2020,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2022,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2023,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2024,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2026,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2027,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2028,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2029,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2030,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2031,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2032,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2034,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2035,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2036,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2037,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2038,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2039,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2040,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2041,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2042,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2043,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2044,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2046,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2047,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2048,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2051,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2052,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2053,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2055,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2056,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2057,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2058,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2060,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2061,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2062,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2064,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2065,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2066,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2067,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2069,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2070,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2071,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2073,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2074,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2075,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2076,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2077,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2079,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2080,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2082,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2083,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2084,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2085,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2086,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2087,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2089,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2090,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2091,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2092,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2093,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2094,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2095,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2096,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2097,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2098,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2101,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2102,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2103,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2104,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2105,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2106,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2108,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2109,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2110,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2111,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2112,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2113,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2114,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2116,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2117,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2118,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2119,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2121,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2123,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2124,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2125,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2126,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2127,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2128,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2129,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2130,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2131,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2132,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2133,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2134,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2136,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2137,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2138,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2140,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2141,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2143,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2144,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2145,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2148,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2149,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2151,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2153,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2154,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2156,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2157,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2158,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2160,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2161,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2162,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2163,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2164,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2165,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2166,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2167,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2168,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2170,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2171,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2172,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2173,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2174,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2175,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2176,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2177,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2179,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2180,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2181,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2183,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2184,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2185,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2186,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2187,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2188,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2190,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2193,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2194,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2195,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2197,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2198,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2199,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2200,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2203,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2204,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2205,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2207,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2208,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2209,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2210,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2211,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2212,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2213,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2214,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2215,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2216,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2217,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2219,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2220,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2221,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2223,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2224,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2225,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2226,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2227,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2228,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2229,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2231,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2233,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2234,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2235,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2236,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2238,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2239,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2240,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2242,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2243,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2244,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2246,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2247,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2248,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2249,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2250,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2251,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2253,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2254,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2255,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2256,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2257,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2258,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2259,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2260,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2262,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2263,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2264,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2265,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2266,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2267,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2269,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2270,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2271,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2272,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2273,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2274,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2276,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2277,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2278,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2279,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2280,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2282,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2283,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2284,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2286,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2287,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2288,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2290,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2291,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2292,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2293,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2295,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2296,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2298,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2299,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2300,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2302,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2303,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2304,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2305,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2306,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2308,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2309,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2310,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2311,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2313,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2314,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2315,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2317,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2318,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2319,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2320,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2321,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2322,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2324,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2325,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2326,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2328,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2329,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2332,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2333,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2334,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2336,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2337,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2338,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2339,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2340,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2341,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2342,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2343,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2344,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2345,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2346,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2347,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2348,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2350,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2352,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2353,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2355,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2356,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2357,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2358,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2360,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2361,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2362,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2363,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2364,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2365,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2366,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2367,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2368,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2369,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2370,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2371,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2373,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2374,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2376,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2377,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2378,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2379,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2380,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2382,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2383,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2384,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2385,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2386,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2387,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2388,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2389,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2390,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2391,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2392,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2393,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2395,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2396,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2397,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2398,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2401,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2402,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2404,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2405,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2406,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2407,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2409,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2410,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2411,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2412,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2413,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2414,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2415,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2416,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2417,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2419,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2420,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2421,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2422,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2424,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2425,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2426,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2427,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2428,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2429,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2430,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2431,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2432,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2434,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2435,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2436,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2437,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2438,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2439,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2441,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2442,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2443,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2444,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2445,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2446,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2448,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2451,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2452,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2454,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2455,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2456,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2457,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2459,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2460,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2461,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2463,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2464,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2465,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2466,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2467,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2468,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2469,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2471,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2473,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2474,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2475,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2476,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2477,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2478,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2479,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2481,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2482,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2483,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2484,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2485,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2486,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2487,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2488,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2490,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2491,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2492,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2493,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2494,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2495,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2497,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2498,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2499,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2500,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2501,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2502,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2503,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2505,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2506,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2507,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2508,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2509,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2511,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2512,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2514,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2515,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2516,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2517,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2518,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2519,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2521,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2522,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2523,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2524,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2525,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2526,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2527,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2529,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2531,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2532,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2533,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2534,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2535,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2536,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2537,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2538,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2540,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2542,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2543,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2545,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2546,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2547,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2548,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2550,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2551,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2553,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2554,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2555,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2557,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2558,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2559,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2560,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2561,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2562,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2563,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2564,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2565,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2566,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2567,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2568,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2569,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2571,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2572,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2574,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2575,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2576,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2577,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2579,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2580,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2581,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2582,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2585,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2586,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2588,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2589,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2590,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2591,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2592,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2593,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2594,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2595,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2596,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2597,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2600,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2601,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2602,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2603,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2604,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2605,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2606,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2608,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2610,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2611,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2612,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2613,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2614,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2615,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2616,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2617,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2618,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2619,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2620,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2624,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2625,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2626,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2627,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2628,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2629,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2631,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2632,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2633,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2634,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2635,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2637,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2638,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2640,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2641,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2642,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2643,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2644,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2645,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2646,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2648,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2650,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2651,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2652,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2653,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2654,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2655,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2657,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2658,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2659,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2661,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2662,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2663,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2664,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2665,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2666,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2667,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2668,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2669,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2672,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2673,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2674,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2675,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2676,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2678,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2679,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2680,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2681,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2683,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2684,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2685,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2686,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2687,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2689,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2690,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2691,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2692,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2693,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2695,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2696,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2698,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2699,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2700,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2701,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2702,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2703,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2704,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2707,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2708,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2709,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2710,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2711,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2713,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2714,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2717,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2719,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2721,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2722,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2723,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2724,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2725,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2727,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2728,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2730,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2731,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2732,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2733,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2734,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2735,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2736,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2737,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2738,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2739,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2740,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2742,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2743,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2744,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2745,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2748,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2749,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2750,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2751,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2752,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2754,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2755,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2756,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2757,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2758,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2760,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2761,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2763,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2764,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2765,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2766,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2767,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2768,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2769,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2770,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2771,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2772,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2773,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2774,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2775,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2776,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2778,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2779,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2780,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2781,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2782,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2783,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2784,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2785,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2786,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2788,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2789,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2790,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2792,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2793,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2794,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2795,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2796,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2797,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2798,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2799,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2800,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2803,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2804,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2805,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2807,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2808,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2809,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2810,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2811,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2813,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2814,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2815,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2816,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2817,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2818,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2819,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2820,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2821,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2823,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2824,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2825,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2827,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2828,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2829,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2830,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2833,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2834,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2836,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2837,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2838,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2839,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2840,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2841,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2842,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2843,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2844,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2845,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2846,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2847,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2849,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2850,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2851,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2852,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2853,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2854,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2855,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2856,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2857,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2859,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2860,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2861,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2862,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2863,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2864,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2865,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2867,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2868,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2869,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2872,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2873,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2874,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2875,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2876,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2878,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2879,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2880,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2882,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2883,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2884,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2885,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2886,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2887,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2888,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2889,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2890,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2892,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2893,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2894,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2895,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2896,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2897,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2898,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2899,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2900,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2901,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2903,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2904,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2906,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2907,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2908,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2909,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2910,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2913,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2914,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2915,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2916,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2917,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2918,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2919,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2920,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2922,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2923,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2924,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2925,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2926,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2927,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2928,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2931,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2932,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2933,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2934,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2935,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2936,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2937,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2939,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2940,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2941,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2942,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2944,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2945,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2946,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2947,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2948,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2949,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2950,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2951,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2952,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2953,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2955,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2956,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2957,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2958,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2959,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2962,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2963,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2964,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2965,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2966,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2968,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2969,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2970,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2971,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2972,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2973,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2974,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2975,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2976,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2979,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2980,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2981,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2982,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2983,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2985,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2986,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2987,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2988,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2989,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2990,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2991,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2993,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2994,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2995,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2996,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2997,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2998,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2999,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3000,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3001,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3003,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3004,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3005,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3007,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3008,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3009,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3010,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3012,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3013,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3014,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3015,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3016,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3017,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3018,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3019,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3020,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3021,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3022,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3023,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3025,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3026,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3027,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3028,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3030,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3031,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3034,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3035,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3036,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3037,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3039,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3040,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3041,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3042,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3043,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3044,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3046,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3047,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3048,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3049,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3051,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3052,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3053,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3054,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3055,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3057,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3058,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3059,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3061,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3063,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3064,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3065,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3067,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3069,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3070,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3071,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3073,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3075,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3076,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3078,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3079,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3080,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3081,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3082,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3083,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3086,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3087,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3088,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3089,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3090,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3092,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3093,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3094,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3096,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3097,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3098,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3100,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3101,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3102,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3103,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3104,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3105,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3107,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3108,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3109,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3110,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3111,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3112,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3113,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3115,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3116,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3117,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3118,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3119,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3120,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3121,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3122,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3124,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3125,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3126,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3127,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3128,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3130,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3131,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3133,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3134,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3135,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3136,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3137,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3138,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3139,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3140,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3141,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3142,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3143,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3144,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3147,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3149,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3150,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3151,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3152,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3153,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3155,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3156,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3158,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3159,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3160,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3161,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3162,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3163,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3164,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3165,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3166,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3167,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3168,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3169,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3170,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3171,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3173,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3174,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3175,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3176,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3177,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3178,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3179,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3181,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3182,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3183,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3185,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3186,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3187,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3188,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3189,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3191,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3192,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3193,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3194,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3195,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3196,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3197,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3198,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3199,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3200,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3201,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3203,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3205,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3206,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3208,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3209,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3210,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3211,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3212,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3213,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3215,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3216,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3217,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3219,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3220,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3221,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3222,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3223,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3224,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3225,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3226,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3227,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3229,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3230,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3231,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3232,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3233,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3234,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3235,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3238,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3239,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3240,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3241,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3242,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3243,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3244,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3245,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3246,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3247,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3248,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3249,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3250,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3252,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3253,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3255,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3256,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3257,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3258,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3259,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3261,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3262,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3264,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3265,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3266,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3267,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3268,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3269,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3270,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3271,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3272,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3273,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3274,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3275,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3276,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3277,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3279,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3280,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3282,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3283,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3284,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3285,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3286,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3288,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3289,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3290,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3292,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3293,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3295,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3296,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3297,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3298,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3300,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3301,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3302,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3304,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3305,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3307,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3308,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3309,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3310,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3313,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3314,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3315,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3316,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3317,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3318,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3319,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3320,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3321,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3323,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3324,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3325,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3327,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3328,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3329,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3330,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3331,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3333,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3334,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3336,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3337,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3338,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3339,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3340,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3341,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3342,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3343,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3344,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3345,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3346,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3348,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3349,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3350,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3351,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3353,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3354,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3355,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3356,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3357,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3358,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3360,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3361,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3364,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3366,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3368,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3369,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3371,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3372,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3373,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3374,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3375,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3376,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3377,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3378,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3379,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3380,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3381,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3384,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3385,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3387,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3389,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3390,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3391,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3392,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3393,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3395,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3396,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3397,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3399,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3400,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3401,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3402,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3403,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3404,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3405,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3406,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3407,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3410,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3411,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3413,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3414,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3415,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3416,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3417,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3418,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3419,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3420,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3421,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3422,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3423,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3424,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3425,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3426,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3427,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3429,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3430,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3431,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3433,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3434,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3435,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3436,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3437,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3438,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3439,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3442,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3443,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3444,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3446,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3447,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3448,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3450,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3451,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3452,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3453,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3454,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3455,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3456,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3457,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3458,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3459,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3461,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3462,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3465,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3466,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3468,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3470,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3471,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3473,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3474,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3475,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3476,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3478,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3479,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3481,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3482,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3483,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3485,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3486,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3487,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3488,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3489,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3491,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3492,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3493,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3495,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3496,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3497,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3498,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3500,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3501,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3502,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3504,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3505,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3506,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3507,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3508,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3510,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3511,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3512,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5430,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5437,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5449,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5452,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5456,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5457,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5462,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5468,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5477,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5480,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5501,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5505,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5507,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5529,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5530,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5534,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5538,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5564,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5566,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5575,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5580,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5618,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5625,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5627,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5669,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5672,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5677,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5680,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5684,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5687,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5692,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5694,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5697,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5700,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5705,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5707,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5711,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5714,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5719,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5722,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5727,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5729,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5732,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5735,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5741,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5743,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5747,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5750,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5755,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5759,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5762,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5766,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5770,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5776,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5778,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8064,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8072,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8078,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8085,
	DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N16704;
assign bdw_enable = !astall;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1425 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1429 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1425 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1429);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1449 = !(b_exp[0] & b_exp[1]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1451 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8072 = !((b_exp[7] & b_exp[6]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1451);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1449 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8072);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1485 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1489 = !(((b_man[0] | b_man[1]) | b_man[2]) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1485);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1472 = !(b_man[10] | b_man[9]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1491 = !(b_man[6] | b_man[5]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1480 = !(b_man[8] | b_man[7]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1500 = !(b_man[4] | b_man[3]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1483 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1472 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1491) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1480) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1500);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1494 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1504 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20 = !((((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1489) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1483) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1494) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1504);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20 | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__18 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__20;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N269 = !(((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1314 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1318 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1314 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1318);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1338 = !(a_exp[0] & a_exp[1]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1340 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8064 = !((a_exp[7] & a_exp[6]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1340);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1338 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8064);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1374 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1378 = !(((a_man[0] | a_man[1]) | a_man[2]) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1374);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1361 = !(a_man[10] | a_man[9]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1380 = !(a_man[6] | a_man[5]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1369 = !(a_man[8] | a_man[7]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1389 = !(a_man[4] | a_man[3]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1372 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1361 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1380) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1369) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1389);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1383 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1393 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19 = !((((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1378) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1372) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1383) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1393);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19 | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__17 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__19;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N270 = !(((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N269 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N270;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N268 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N267 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29 = ((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N268) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N267;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5452 = !a_exp[7];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5456 = b_exp[0] | a_exp[0];
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5449, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]} = {1'B0, a_exp[1]} + {1'B0, b_exp[1]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5456};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5468, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]} = {1'B0, a_exp[2]} + {1'B0, b_exp[2]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5449};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5480, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]} = {1'B0, a_exp[3]} + {1'B0, b_exp[3]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5468};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5462, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]} = {1'B0, a_exp[4]} + {1'B0, b_exp[4]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5480};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5477, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]} = {1'B0, a_exp[5]} + {1'B0, b_exp[5]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5462};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5457, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]} = {1'B0, a_exp[6]} + {1'B0, b_exp[6]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5477};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]} = {1'B0, b_exp[7]} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5452} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5457};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9] = !(a_exp[7] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5564 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5529 = (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5538 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0] = (!b_exp[0]) ^ a_exp[0];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5530 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8] = (!a_exp[7]) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5472;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5534 = !((((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5530) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8]) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N273 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5534 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5538) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5529));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5566 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5564 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N273);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5430 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__26 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__22);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5437 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__25 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__21);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N272 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5437 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__24);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30 = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N272) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5430 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__23);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5507 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5505 = ((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5501 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5505);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N276 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5507 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5501);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8078 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N276);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__41 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8078 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__41;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__60 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5566 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5580 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5575 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N274 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5580 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5575);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8085 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[8] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N274);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__42 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N8085 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__30 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__42;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__61 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__32 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[9]) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 = !a_man[22];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1991 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905 = !b_man[22];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3087 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3094 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480 = !b_man[21];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2231 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 = !a_man[21];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2250 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688;
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2066, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1641} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2231} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3094} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2250};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3087} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1991} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2066};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3357 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049 = !b_man[20];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3341 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2240 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3426, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2994} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3341} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3357} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2240};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 = !a_man[20];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1657 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623 = !b_man[19];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2486 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2502 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1962, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3495} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2486} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1657} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2502};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2512 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261;
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2319, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1887} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2512} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1962} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2994};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3426} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1641} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2319};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3349 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 = !a_man[19];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2769 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1911 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157 = !b_man[18];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1628 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2761 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1610, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3141} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1628} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1911} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2761};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2820, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2390} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2769} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3349} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1610};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1647 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 = !a_man[18];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3026 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2494 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2466, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2030} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3026} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1647} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2494};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1716, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3245} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2466} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3495} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2390};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2820} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1887} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1716};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 = !a_man[17];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2436 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301 = !b_man[16];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1878 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3277 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2253, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1824} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1878} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2436} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3277};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1638 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2163 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 = !a_man[16];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1587 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3010 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3107, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2683} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1587} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2163} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3010};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2108, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1684} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1638} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2253} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3107};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1903 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3286 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2751 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3215, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2788} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3286} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1903} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2751};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2170 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729 = !b_man[17];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2736 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3018 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2362, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1929} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2736} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2170} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3018};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2743 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1893 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2690 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871 = !b_man[15];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2983 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1574 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3255, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2829} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2983} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2690} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1574};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2003, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1576} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1893} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2743} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3255};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2964, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2540} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1929} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2788} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2003};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2212, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1781} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2030} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2108} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2964};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3319, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2890} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2362} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3215} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3141};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3319} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2212} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3245};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2999 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2154 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1885 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3003, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2579} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2154} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2999} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1885};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2426 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 = !a_man[15];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1843 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3270 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2149, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1725} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1843} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2426} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3270};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2859, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2434} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2149} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3003} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1824};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2681 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 = !a_man[14];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2102 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1564 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2293, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1866} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2102} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2681} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1564};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2949 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412 = !b_man[14];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2128 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1835 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3404, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2972} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2128} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2949} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1835};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3262 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2416 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2145 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3150, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2722} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2416} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3262} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2145};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1896, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3435} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3404} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2293} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3150};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1750, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3288} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2683} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1896} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1576};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1858, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3395} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2859} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1684} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1750};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2890} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1858} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1781};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2756, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2328} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2829} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1725} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2579};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1556 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2672 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2407 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2444, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2010} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2672} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1556} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2407};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2898, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2475} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2444} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2972} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1866};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3209 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978 = !b_man[13];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3235 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2092 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2691, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2263} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3235} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3209} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2092};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2991 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2941 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 = !a_man[13];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2365 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1826 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1585, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3117} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2365} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2941} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1826};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2039, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1619} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2991} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2691} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1585};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1650, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3181} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2039} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2898} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3435};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2610, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2179} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2756} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2434} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1650};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2540} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2610} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3395};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2137 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3253 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3466 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556 = !b_man[12];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2380 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2357 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3083, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2659} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2380} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3466} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2357};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3296, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2868} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3253} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2137} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3083};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1816 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2928 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2664 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2839, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2411} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2928} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1816} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2664};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3199 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 = !a_man[12];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2620 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2083 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1979, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1553} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2620} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3199} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2083};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2397 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3511 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3244 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1734, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3264} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3511} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2397} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3244};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2188, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1760} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1979} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2839} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1734};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1791, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3327} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2722} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3296} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2188};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3043, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2618} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2263} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3117} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2010};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2650, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2221} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3043} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1619} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2475};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2505, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2075} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1791} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2328} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2650};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3288} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2505} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2179};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3457 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 = !a_man[11];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2880 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2345 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3479, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3054} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2880} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3457} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2345};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1762 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122 = !b_man[11];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3483 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2613 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2626, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2197} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3483} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1762} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2613};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2074 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3192 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2920 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2379, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1950} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3192} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2074} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2920};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2588, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2160} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2626} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3479} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2379};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2658 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1809 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3502 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3232, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2807} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1809} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2658} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3502};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3443, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3013} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3232} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2659} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1553};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1939, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3472} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2588} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2868} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3443};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2018 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702 = !b_man[10];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2629 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2873 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3273, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2846} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2629} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2018} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2873};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2388 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1755 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 = !a_man[10];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3139 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2604 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2166, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1739} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3139} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1755} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2604};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2124, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1704} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2388} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3273} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2166};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2336, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1905} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2411} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3264} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2124};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2797, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2370} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1760} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2336} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2618};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3505, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3075} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1939} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3327} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2797};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3181} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3505} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2075};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033;
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1875, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3413} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3054} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1950} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2807};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2914 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2065 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1801 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1914, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3450} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2065} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2914} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1801};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2338 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3449 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3183 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3020, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2597} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3449} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2338} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3183};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2982, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2559} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3020} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1914} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2197};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3193, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2765} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2982} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1875} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2160};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2595 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1747 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3442 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2814, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2387} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1747} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2595} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3442};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2012 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 = !a_man[9];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3401 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2861 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1958, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3487} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3401} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2012} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2861};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3174 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2326 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2057 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1712, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3241} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2326} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3174} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2057};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1667, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3200} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1958} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2814} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1712};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3492 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2648 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2283 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228 = !b_man[9];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1769 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3128 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3063, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2635} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1769} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2283} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3128};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2772, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2343} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2648} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3492} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3063};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1787 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2904 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2638 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2566, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2131} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2904} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1787} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2638};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2525, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2094} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2566} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2846} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1739};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2731, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2304} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2772} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1667} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2525};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2084, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1660} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3013} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2731} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1905};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1694, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3223} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3193} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3472} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2084};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2221} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1694} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3075};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2274 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 = !a_man[8];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1701 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3119 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2854, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2428} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1701} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2274} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3119};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2547 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806 = !b_man[8];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2879 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3391 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1998, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1569} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2879} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2547} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3391};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2853 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2005 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1741 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1745, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3282} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2005} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2853} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1741};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3420, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2990} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1998} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2854} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1745};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3377, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2947} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2597} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3450} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3420};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1627, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3161} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1704} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3377} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2559};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2048 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3167 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2896 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3459, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3028} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3167} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2048} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2896};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3434 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2590 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2318 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2605, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2174} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2590} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3434} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2318};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2314, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1880} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2605} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3459} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2635};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3168, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2738} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3487} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2387} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3241};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2270, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1844} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2343} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2314} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3168};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2483, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2051} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3413} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2270} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2304};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2939, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2517} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1627} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2765} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2483};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2370} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2939} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3223};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2803 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375 = !b_man[7];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2020 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1692 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2034, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1611} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2020} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2803} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1692};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1779 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2537 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 = !a_man[7];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1954 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3379 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2894, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2469} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1954} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2537} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3379};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2355, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1924} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1779} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2034} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2894};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1733 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2844 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2581 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2642, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2215} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2844} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1733} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2581};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3111 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2265 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1997 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1785, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3323} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2265} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3111} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1997};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2309 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3425 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3159 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3500, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3069} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3425} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2309} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3159};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3211, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2782} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1785} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2642} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3500};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2060, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1636} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2131} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2355} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3211};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3126, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2699} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3200} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2094} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2060};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2103, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1676} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1569} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2428} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3282};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2888 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2038 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3059 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948 = !b_man[6];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3127 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1947 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3185, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2760} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3127} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3059} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1947};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2395, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1965} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2038} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2888} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3185};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2957, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2535} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2174} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3028} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2395};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2916, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2490} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2103} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2990} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2957};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2016, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1593} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2947} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2916} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1844};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3336, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2909} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3126} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3161} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2016};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1660} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3336} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2517};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3147 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2300 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2029 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1580, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3109} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2300} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3147} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2029};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2572 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1723 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3419 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2686, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2257} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1723} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2572} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3419};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2143, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1719} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2686} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1580} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1611};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3372 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2527 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2255 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2934, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2507} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2527} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3372} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2255};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2794 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 = !a_man[6];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2211 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1681 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2079, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1654} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2211} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2794} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1681};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1987 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3101 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2838 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1828, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3366} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3101} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1987} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2838};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3248, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2823} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2079} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2934} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1828};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2997, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2574} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2469} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3323} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2215};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1853, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3389} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3248} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2143} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2997};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1810, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3346} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1880} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2738} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1853};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3049 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 = !a_man[5];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2474 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1936 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2373, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1944} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2474} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3049} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1936};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3318 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477 = !b_man[5];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2273 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2205 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3474, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3046} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2273} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3318} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2205};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1671 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2784 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2519 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3226, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2800} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2784} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1671} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2519};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2438, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2007} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3474} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2373} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3226};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2828 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1981 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1715 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2975, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2553} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1981} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2828} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1715};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2246 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3364 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3092 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2118, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1698} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3364} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2246} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3092};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3411 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2565 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2291 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1869, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3407} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2565} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3411} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2291};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3292, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2863} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2118} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2975} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1869};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1889, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3429} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3069} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2438} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3292};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2708, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2279} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1924} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2782} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1889};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2667, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2238} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1636} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2708} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2490};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2876, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2451} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1810} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2699} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2667};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2051} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2876} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2909};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370;
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2183, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1753} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2760} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1654} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2507};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2750, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2322} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1965} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2183} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2823};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1603, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3137} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1676} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2535} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2750};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3036, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2615} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3366} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2257} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3109};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1644, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3175} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3036} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1719} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2574};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2461, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2026} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3389} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1644} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2279};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1559, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3090} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1603} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3346} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2461};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1593} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1559} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2451};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3330, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2903} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2800} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1698} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2553};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2792, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2363} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3330} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2007} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2863};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2509 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1662 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3354 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1555, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3086} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1662} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2509} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3354};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1926 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3041 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2774 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2661, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2233} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3041} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1926} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2774};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3082 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2236 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1973 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2414, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1983} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2236} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3082} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1973};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1622, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3155} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2661} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1555} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2414};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1618 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050 = !b_man[4];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3381 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2465 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2913, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2485} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3381} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1618} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2465};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3138 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3310 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 = !a_man[4];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2730 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2193 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1807, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3340} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2730} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3310} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2193};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2725, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2298} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3138} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2913} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1807};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1708 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2819 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2555 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3267, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2840} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2819} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1708} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2555};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2478, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2042} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3267} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3046} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1944};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1934, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3468} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2725} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1622} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2478};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2498, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2069} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1934} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2792} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3429};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2282 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3403 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1874 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623 = !b_man[3];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2526 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2721 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3453, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3022} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2526} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1874} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2721};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2162, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1736} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3403} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2282} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3453};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2185 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3302 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3031 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3203, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2775} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3302} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2185} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3031};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1609 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 = !a_man[3];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2989 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2457 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2348, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1918} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2989} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1609} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2457};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2767 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1916 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1652 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2097, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1669} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1916} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2767} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1652};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3016, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2591} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2348} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3203} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2097};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2224, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1796} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3407} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2162} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3016};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1686, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3219} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2224} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1753} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2615};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3356, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2924} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2322} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1686} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3175};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3315, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2885} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2498} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3137} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3356};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2238} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3315} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3090};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306;
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1664, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3195} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3086} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1983} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2840};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1974, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3510} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1664} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3155} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2042};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2768, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2340} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2485} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3340} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2233};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1964 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3073 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2813 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1847, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3380} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3073} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1964} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2813};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3345 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2500 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2229 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2952, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2529} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2500} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3345} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2229};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2546 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1700 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3393 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2702, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2272} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1700} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2546} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3393};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1908, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3446} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2952} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1847} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2702};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3078, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2653} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1908} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2768} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2298};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2545, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2111} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3078} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1974} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2363};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1643 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2758 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2492 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2637, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2208} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2758} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1643} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2492};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3023 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2176 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1909 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1780, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3317} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2176} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3023} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1909};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2220 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3338 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3065 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3491, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3064} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3338} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2220} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3065};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2454, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2019} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1780} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2637} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3491};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1865 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 = !a_man[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3247 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2711 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2028, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1606} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3247} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1865} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2711};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2134 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196 = !b_man[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1670 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2981 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3140, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2710} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1670} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2134} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2981};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2449 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1602 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3293 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2887, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2463} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1602} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2449} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3293};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1597, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3130} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3140} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2028} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2887};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2518, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2087} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1597} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2454} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1736};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2833, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2404} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2903} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2518} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1796};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3399, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2965} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3468} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2833} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3219};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2247, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1818} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2545} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2069} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3399};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2026} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2247} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2885};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765 = !b_man[1];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2776 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2393 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1969, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3501} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2776} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2393};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2536 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3239 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 = !a_man[1];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3508 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2123 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2824, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2398} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3508} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3239} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2123};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3243, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2816} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2536} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1969} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2824};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3057, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2628} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3380} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2272} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3243};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2200, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1771} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2775} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1669} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2529};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2267, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1838} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2200} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3057} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2340};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2805 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1957 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1691 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2389, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1960} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1957} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2805} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1691};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3309, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2878} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2389} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3022} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1918};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3374, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2944} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3309} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2591} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3446};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1728, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3257} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3374} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2267} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2653};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2210 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3329 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3058 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3178, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2752} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3329} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2210} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3058};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1634 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2748 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2482 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2325, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1892} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2748} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1634} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2482};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2796 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1946 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1680 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2071, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1646} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1946} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2796} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1680};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2993, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2569} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2325} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3178} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2071};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2442 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1591 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3283 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2576, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2144} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1591} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2442} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3283};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1856 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2971 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2704 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1722, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3252} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2971} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1856} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2704};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3015 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2168 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1900 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3430, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3000} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2168} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3015} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1900};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2136, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1714} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1722} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2576} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3430};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1884, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3422} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2710} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1606} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2463};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1953, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3482} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2136} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2993} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1884};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2742, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2317} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3317} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2208} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3064};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2811, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2382} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2742} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3130} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2019};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3118, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2695} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3195} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1953} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2811};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2582, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2153} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3118} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3510} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2404};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2286, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1862} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1728} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2111} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2582};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2924} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2286} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1818};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303 = !b_man[0];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1915 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2652 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2763, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2334} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1915} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2652};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3498 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 = !a_man[0];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1806 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2386 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1656, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3188} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1806} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3498} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2386};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2927, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2501} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2763} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3501} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1656};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2696 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1849 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1582 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3368, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2937} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1849} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2696} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1582};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2114 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3231 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2963 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2511, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2082} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3231} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2114} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2963};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3275 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2431 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2161 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2260, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1830} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2431} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3275} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2161};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1821, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3358} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2511} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3368} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2260};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1639, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3171} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1960} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2927} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1821};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1707, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3234} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1639} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2878} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1771};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2014, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1590} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2087} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2944} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1707};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2473 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1626 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3321 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2008, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1583} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1626} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2473} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3321};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1891 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3005 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2740 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3113, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2689} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3005} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1891} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2740};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3048 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2204 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1935 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2865, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2441} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2204} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3048} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1935};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2679, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2249} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3113} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2008} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2865};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1572, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3103} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2398} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3252} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2144};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2493, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2061} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2679} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2816} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1572};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2430, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1999} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3000} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1892} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2752};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3348, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2919} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2430} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1714} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2569};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2563, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2127} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2628} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2493} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3348};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2872, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2445} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2563} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1838} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2695};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3438, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3007} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2014} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3257} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2872};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2965} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3438} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1862};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2905);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1592 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2786 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1757, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3295} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2786} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1592} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2334};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2106 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3222 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2953 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2194, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1764} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3222} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2106} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2953};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3486 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2641 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2378 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3304, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2874} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2641} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3486} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2378};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2687 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1841 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1571 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3047, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2624} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1841} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2687} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1571};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2616, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2186} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3304} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2194} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3047};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3284, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2856} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1646} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1757} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2616};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2242, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1813} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3284} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3422} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2317};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3416, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2985} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3482} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2382} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2242};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1882 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2996 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2733 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2804, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2374} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2996} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1882} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2733};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3268 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2421 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2151 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1949, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3476} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2421} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3268} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2151};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2464 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1617 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3314 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1699, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3229} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1617} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2464} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3314};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3470, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3039} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1949} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2804} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1699};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3040 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2195 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1925 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3114 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2557, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2121} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2195} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3040} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1925};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2367, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1938} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2557} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3188} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2082};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2177, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1748} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3470} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2501} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2367};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3220, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2795} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2937} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1830} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2689};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3030, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2606} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3220} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3358} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2249};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3093, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2668} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2177} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3171} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3030};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2308, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1877} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3093} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3234} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2127};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1761, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3300} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3416} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1590} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2308};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2153} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1761} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3007};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3121 = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2911) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1794;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2053 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2480);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2901 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2129, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1709} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2053} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2901};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2634 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1784 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3478 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2986, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2564} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1784} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2634} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3478};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3410, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2976} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2129} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3121} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2986};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2113, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1690} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1583} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2441} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3410};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1927, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3461} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2113} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3103} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1999};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1990, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1563} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2061} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2919} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1927};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1832 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2945 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2678 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2737, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2310} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2945} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1832} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2678};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3213 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2369 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2098 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1879, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3418} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2369} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3213} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2098};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2413 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1561 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3259 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1633, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3166} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1561} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2413} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3259};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2299, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1872} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1879} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2737} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1633};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1608 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2724 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2456 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3342, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2915} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2724} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1608} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2456};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2988 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2141 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1873 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2488, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2056} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2141} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2988} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1873};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2187 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2688 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3301 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3164 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2049);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2041 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1566, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3098} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3164} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2041};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2235, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1808} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3301} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2187} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1566};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3158, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2728} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2488} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3342} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2235};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2968, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2548} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2299} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3295} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3158};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2047, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1624} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2874} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1764} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2624};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1863, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3402} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2047} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2186} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3039};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2785, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2358} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2968} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2856} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1863};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2849, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2422} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2785} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1813} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2668};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3165, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2735} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1990} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2985} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2849};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2445} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3165} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3300};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2906, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2481} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3476} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2374} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3229};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2719, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2290} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2906} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1938} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2795};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1679, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3212} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1748} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2606} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2719};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1776 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2893 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2625 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2425, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1993} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2893} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1776} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2625};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2361 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3471 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3206 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3276, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2852} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3471} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2361} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3206};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3089, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2663} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1709} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2425} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3276};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1554 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2669 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2402 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3025, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2600} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2669} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1554} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2402};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2936 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2089 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1822 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2172, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1744} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2089} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2936} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1822};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2133 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3250 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2980 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1919, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3456} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3250} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2133} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2980};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1984, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1557} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2172} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3025} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1919};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1800, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3333} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2121} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3089} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1984};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2714 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1864 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1601 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2779, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2353} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1864} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2714} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1601};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2843, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2415} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2779} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2564} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3418};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2657, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2227} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2976} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2843} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1872};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1614, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3149} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1800} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1690} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2657};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2306 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3153 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1859, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3396} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2306} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3153};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2448 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2261 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1674, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3205} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2448} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1859} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3098};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2592, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2164} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2915} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1674} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1808};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1738, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3269} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2310} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3166} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2056};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3512, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3081} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1738} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2592} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2728};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2472, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2037} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2548} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3512} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3402};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2538, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2105} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1614} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3461} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2472};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1742, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3274} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1679} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1563} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2538};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1877} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1742} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2735};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3238 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2392 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2126 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2209, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1782} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2392} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3238} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2126};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2662 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1812 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3507 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3320, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2889} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1812} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2662} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3507};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1855 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2970 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2703 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1833 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3067, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2640} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2970} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1855} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2703};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3385, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2956} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3320} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2209} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3067};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3462 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2617 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2350 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1607, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3142} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2617} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3462} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2350};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2884 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2032 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1767 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2713, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2284} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2032} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2884} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1767};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2080 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3197 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2926 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2467, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2031} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3197} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2080} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2926};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2531, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2101} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2713} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1607} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2467};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2277, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1848} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1993} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2852} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1744};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3448, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3017} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2531} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3385} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2277};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2406, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1977} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1624} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2481} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3448};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3325, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2895} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2406} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2290} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3149};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3392, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2959} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2358} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3212} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3325};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2422} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3392} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3274};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3131, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2707} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2600} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3456} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2353};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2342, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1910} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3131} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2663} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1557};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3261, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2836} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2342} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3333} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2227};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3189 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2341 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2070 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1651, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3182} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2341} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3189} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2070};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2608 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1759 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3454 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2754, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2329} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1759} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2608} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3454};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1805 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2918 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2655 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2506, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2073} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2918} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1805} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2655};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2818, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2391} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2754} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1651} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2506};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3415 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3157);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2296 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3004, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2580} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3415} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2296};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2024 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3144 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2875 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1897, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3433} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3144} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2024} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2875};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1963, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3493} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3004} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3396} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1897};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2023, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1600} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1963} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2818} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3205};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3196, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2770} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2415} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3269} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2023};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2156, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1731} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3196} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3081} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1977};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2216, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1788} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3261} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2037} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2156};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2105} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2216} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2959};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2962 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3367 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2117 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2562 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3406 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3042, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2619} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2562} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3406};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2254, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1825} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2117} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2962} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3042};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2385 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3497 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3230 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3360, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2931} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3497} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2385} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3230};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1717, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3246} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3360} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2254} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2284};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2883, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2455} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1717} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2101} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2956};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2091, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1665} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2164} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2883} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3017};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3135 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2288 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2015 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1940, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3473} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2288} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3135} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2015};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1752 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2867 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2601 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2798, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2368} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2867} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1752} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2601};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3108, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2680} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2580} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1940} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2798};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3424, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2995} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1782} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2640} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3108};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2571, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2138} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3142} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2031} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2889};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1773, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3313} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2571} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3424} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1848};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2910 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2062 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1793 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2550, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2116} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2062} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2910} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1793};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2333 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3447 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3179 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1693, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3224} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3447} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2333} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3179};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3489 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2644 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2377 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3405, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2969} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2644} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3489} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2377};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2000, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1577} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1693} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2550} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3405};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2860, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2435} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3433} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2329} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3182};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2320, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1888} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2000} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3493} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2860};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2632, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2203} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2707} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2320} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1600};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2946, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2521} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1773} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1910} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2632};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3009, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2585} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2091} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2836} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2946};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2895} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3009} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1788};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2749 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1705 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2301);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2551 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1980, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1551} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1705} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2551};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3221 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2938 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2292, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1867} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3221} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1980} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2619};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1751, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3285} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2073} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2931} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2292};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3173, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2744} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2391} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1751} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3246};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2857 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2009 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1743 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1735, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3265} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2009} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2857} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1743};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2278 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3397 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3124 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2837, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2412} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3397} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2278} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3124};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3439 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2593 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2324 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2589, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2157} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2593} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3439} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2324};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3151, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2723} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2837} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1735} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2589};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2633 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1783 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3481 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2513 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2337, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1906} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1783} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2633} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3481};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2055 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3170 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2900 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3444, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3014} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3170} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2055} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2900};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2040, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1616} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3444} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2337} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3473};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2611, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2180} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1825} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3151} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2040};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2064, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1642} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2138} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2611} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2995};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3485, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3061} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3173} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2455} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2064};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1840, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3375} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2770} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3485} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1665};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1731} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1840} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2585};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647;
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2897, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2476} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2368} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3224} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2116};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3465, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3034} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2897} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2680} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1577};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2810 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1871);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1696 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1766, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3307} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2810} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1696};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3387 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2543 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2269 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2627, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2198} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2543} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3387} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2269};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3191, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2766} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1766} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1551} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2627};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2586 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1737 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3431 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2376, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1951} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1737} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2586} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3431};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2001 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3116 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2850 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3480, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3052} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3116} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2001} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2850};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3163 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2315 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2044 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3233, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2808} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2315} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3163} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2044};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2085, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1661} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3480} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2376} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3233};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1792, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3328} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2969} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3191} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2085};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2360, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1930} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1792} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2435} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3285};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2922, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2497} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3465} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1888} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2360};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2383, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1956} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3313} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2922} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2203};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2521} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2383} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3375};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1775 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2081 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2892 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1952 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3412);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2799 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2419, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1986} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1952} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2799};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2125, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1703} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2892} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1775} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2419};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2940, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2515} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2125} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2412} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3265};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2651, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2219} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1867} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2940} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2723};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1834, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3371} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2157} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3014} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1906};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3504, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3076} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1834} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1616} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2476};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3216, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2789} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2651} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2180} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3504};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1815, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3350} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2744} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1642} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3216};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3061} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1815} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1956};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2305 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3423 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3152 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1912, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3451} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3423} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2305} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3152};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1730 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2841 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2577 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3021, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2594} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2841} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1730} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2577};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1876, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3414} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3021} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1912} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2198};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2534 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1685 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3376 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3271, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2847} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1685} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2534} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3376};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3105 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2262 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1994 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2167, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1740} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2262} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3105} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1994};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2979, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2560} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3307} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3271} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2167};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2732, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2302} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3052} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1951} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2808};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2692, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2264} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2979} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1876} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2732};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3055 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2978);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1942 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1959, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3488} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3055} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1942};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2036 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1658 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2773, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2344} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2036} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1959} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1986};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2251 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3369 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3096 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1710, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3242} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3369} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2251} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3096};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1675 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2790 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2523 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2815, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2384} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2790} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1675} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2523};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2834 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1985 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1721 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2567, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2132} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1985} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2834} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1721};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1668, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3198} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2815} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1710} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2567};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1625, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3162} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2773} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1703} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1668};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1586, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3115} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2766} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1661} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1625};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2401, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1972} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2692} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3328} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1586};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2109, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1683} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3034} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1930} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2401};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2497} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2109} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3350};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1589 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1589);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2645 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3417 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2568 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2295 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3190 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3421, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2987} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2568} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3417} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2295};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2522, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2095} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3421} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2847} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1740};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2199 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2556);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3044 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2356, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1921} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2199} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3044};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2780 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1932 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1666 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3208, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2783} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1932} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2780} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1666};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2311, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1881} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2356} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3488} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3208};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3378, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2948} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2594} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3451} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2311};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2484, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2052} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2522} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2560} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3378};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2443, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2011} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2515} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3371} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2484};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3256, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2827} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2219} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3076} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2443};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2789} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3256} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1683};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1978 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3088 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2825 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2958, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2533} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3088} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1978} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2825};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3361 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2516 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2243 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2104, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1677} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2516} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3361} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2243};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2561 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2762 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1713 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3308 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2122);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2190 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1645, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3176} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3308} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2190};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1852, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3390} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1713} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2561} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1645};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3169, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2739} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2104} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2958} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1852};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2058, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1637} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2384} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3242} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2132};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2271, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1842} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2344} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3169} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2058};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3337, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2907} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3414} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2302} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2271};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3297, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2869} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2264} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3337} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3115};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1972} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3297} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2827};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1839 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1579 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1839);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3122, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2700} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3198} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2095} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2948};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2228, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1804} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3162} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2052} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3122};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2011} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2228} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2869};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N16704 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2452 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1702);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3298 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1786, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3324} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2452} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3298};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2817 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3100, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2674} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2817} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1786} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3176};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2460, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2027} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2533} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3100} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3390};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3080 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2234 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1968 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2248, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1819} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2234} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3080} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1968};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1604, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3134} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2248} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2783} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1677};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1811, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3344} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1604} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2460} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2739};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1922 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3035 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2771 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2499, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2067} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3035} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1922} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2771};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2503 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1659 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3351 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3353, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2925} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1659} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2503} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3351};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2709, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2280} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1921} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2499} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3353};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2917, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2491} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2987} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2709} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1881};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2017, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1594} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2917} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1811} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1842};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2907} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2017} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1804};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2855, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2429} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2067} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2925} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1819};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1648 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2764 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2495 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3496, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3070} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2764} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1648} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2495};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3027 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2181 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1913 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2643, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2213} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2181} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3027} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1913};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2225 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3343 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3071 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1904 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2396, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1966} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3343} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2225} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3071};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1996, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1570} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2643} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3496} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2396};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3316, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2886} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1996} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2855} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2280};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2665, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2239} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1637} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3316} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2491};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2700} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2665} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1594};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2459 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3280 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2437 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2165 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1581, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3110} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2437} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3280} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2165};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1596 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3228);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2446 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2793, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2364} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1596} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2446};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1894 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3012 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2745 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2439, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2004} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3012} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1894} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2745};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2287, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1860} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2364} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1581} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2439};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2998, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2575} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3070} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1966} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2287};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2603, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2175} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1570} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2998} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2429};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2173 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3290 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3019 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1687, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3217} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3290} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2173} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3019};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3249, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2821} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2793} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3324} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1687};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3334 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3440 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2487 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2701 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2806);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1588 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2684, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2258} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2701} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1588};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3400, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2966} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2487} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3334} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2684};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2755 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1907 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1640 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2542, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2112} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1907} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2755} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1640};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2140, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1720} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2542} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3400} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2213};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1746, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3279} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3249} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2674} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2140};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2207, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1774} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3134} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1746} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2027};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2603} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2886} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1774};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3344} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2207} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2239};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2646 = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1845 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2375);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2693 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3436, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3008} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1845} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2693};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1631 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3011 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3289, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2864} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1631} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3436} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2258};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3143, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2717} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3217} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2112} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3289};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1890, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3427} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2821} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3143} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1720};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3279} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1890} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2175};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3001 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2158 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1886 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2587 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3186, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2757} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2158} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3001} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1886};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2427 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1578 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3272 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2332, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1899} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1578} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2427} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3272};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2184, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1754} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2332} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3186} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3110};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2035, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1612} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2966} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2184} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1860};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2575} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2035} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3427};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2955 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2148 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2155 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3266 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2096 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2942 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1620, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3156} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2096} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2942};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2830, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2405} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3266} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2148} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1620};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2935, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2508} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2830} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1899} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2757};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2951 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1948);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1837 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3477);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3079, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2654} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2951} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1837};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1567 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2685 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2417 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1975, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3506} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2685} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1567} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2417};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2076, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1655} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3079} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3008} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1975};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3037, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2612} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2004} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2076} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2864};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2935} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1754} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2612};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2717} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3037} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1612};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2226 = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2675 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1827 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1558 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2479, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2043} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1827} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2675} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1558};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1729, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3258} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2654} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2479} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3506};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1729} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1655} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2508};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2352 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3201 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3050);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2086 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2973, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2554} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3201} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2086};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2409 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1732 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3331, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2899} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2409} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2973} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3156};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3331} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2405} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3258};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3455 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1817 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2932 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2666 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3263 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1870, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2932} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1817} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2666};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1870} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2043} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2899};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2602 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2347 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2623);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3194 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3227, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2347} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3194};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2077 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2923 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2835 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3452 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2196);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2339 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765);
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2371, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3452} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2339};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2119, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2923} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2077} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2371};
assign {DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294} = {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3227} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2554} + {1'B0, DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2119};
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1584 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2851 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1995 = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3097 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2244 = ((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3303 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1798) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3335) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1765;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2673 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3184 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1945);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2631 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2244 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3097) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2673);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2130 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1995) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2631)) | ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2801) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1695));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2424 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3408 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2294);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1632 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2130 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2851) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2424);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2842 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1584) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1632)) | ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2726) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1797));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2171 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2222 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2150);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2090 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2842 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2602) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2171);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3051 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3455) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2090)) | ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2583) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3363));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1920 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1829 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3469);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2046 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3051 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2352) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1920);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2778 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1931 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2470);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1673 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2891 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2323);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1799 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2778 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2100) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1673);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2514 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2046) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2226)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1799);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2532 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2747 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3029);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3384 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3460 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2636);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2259 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2532 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3384);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3104 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2259;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2471 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1851 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2955) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2514) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3104);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2276 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3062 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3091);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3133 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1560 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2450);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2217 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2276 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1599) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3133);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2432 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2471) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2646)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2217);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2022 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2877 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2660);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2882 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3084 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1758);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1961 = (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2022 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2882;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1883 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3312 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2459) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2432) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1961);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2256 = (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N16704 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1883) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2189 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1726);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3373 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2147 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2541);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2266 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2961 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2245);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3112 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3373 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2694) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2266);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2256) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1579)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3112);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3120 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2671 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2812);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2013 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3237 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2268);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3120 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2447) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2013);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2697 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3441);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1763 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1902 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2647);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2862 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1763);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2214 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3291)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2862);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2645) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2214);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3072 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1854);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3475 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2281 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2169);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3475);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2598 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1630);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3225 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2054 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2192);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2614 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3225);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3038)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2614);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2622 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1898);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2974 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2331 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2716);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2974);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3146 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2677);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2727 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3099 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1778);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2366 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2727);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1967 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2791)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2366);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2321 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2394) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1967);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2749)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2321);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2206 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1989);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2477 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2418 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3306);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2477);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1768 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1803);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2223 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2230 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3370);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2110 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2223);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2544)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2110);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1836 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2115);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1976 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2549 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1971);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1976);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2400 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2930);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1727 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3362 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3033);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1861 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1727);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1718 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2289)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1861);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3177 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1718);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3355 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3177;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2142 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3355);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3464 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2285);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3437 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2712 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2639);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3437);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3066 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2139);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3187 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2746 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2570);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1613 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3187);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3458 = !(((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1613));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2033) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3458);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2496 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3172);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2933 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3352 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2921);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2468 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2933);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2313 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2468;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741 = !(((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2313);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__61) | ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47]) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__60));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[46] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2741) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2159;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56 | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[47] | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1552 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1923;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1982 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2078;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2410 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1552)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1982);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[45] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2410) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3365;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5705 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[46]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[45]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[22] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5705);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[44] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2848 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2510;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5766 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[45]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[44]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[21] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5766);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2908 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3240 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3145;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1820;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1711 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2715;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3240) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1711);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3339 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2330;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1802 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2908)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3339);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[43] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1802) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1653;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5719 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[44]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[43]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[20] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5719);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[42] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2135 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2759;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5669 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[43]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[42]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[19] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5669);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2303 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2241;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2734 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2584;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3160 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2303)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2734);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[41] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3160) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1901;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5732 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[42]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[41]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[18] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5732);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[40] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2423 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3006;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5684 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[41]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[40]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[17] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5684);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3251) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2822);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3398)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2967);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2558 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2832);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[39] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2558 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2152;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5747 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[40]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[39]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[16] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5747);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[38] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3490) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3260;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5697 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[39]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[38]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[15] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5697);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3281;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2809 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3077);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[37] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2809 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2403;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5759 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[38]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[37]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[14] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5759);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[36] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1992) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3509;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5711 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[37]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[36]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[13] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5711);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2068;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1689)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3218);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3053 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3332);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[35] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3053 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2656;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5776 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[36]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[35]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[12] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5776);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[34] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1777) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1795;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5727 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[35]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[34]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[11] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5727);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1814;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3305 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1621);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[33] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3305 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2902;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5677 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[34]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[33]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[10] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5677);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[32] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1562) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2045;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5741 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[33]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[32]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[9] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5741);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2698 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3136 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1933;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2676 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3499;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3102 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3068;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2676)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3102);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1605 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3467;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3136) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1605);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3125 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1868;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1595 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2698)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3125);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[31] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1595) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3154;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5692 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[32]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[31]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[8] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5692);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[30] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2025 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2297;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5755 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[31]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[30]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[7] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5755);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2093 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1568;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2524 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2120;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2950 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2093)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2524);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[29] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2950) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3409;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5707 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[30]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[29]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[6] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5707);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[28] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3095 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2552;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5770 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[29]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[28]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[5] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5770);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2182)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1756);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2346 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2372);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[27] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2346 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1697;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5722 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[28]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[27]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[4] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5722);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[26] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3388) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2802;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5672 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[27]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[26]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[3] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5672);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3428;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2596 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2621);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[25] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2596 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1943;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5735 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[26]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[25]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[2] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5735);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[24] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2670) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3045;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5687 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[25]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[24]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[1] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5687);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1988 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3299;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2781 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2440;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3210 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2006;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1678 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3322 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2781) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N3210);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2420 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2871;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2845 = ((!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1678) & (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N1988)) | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2420);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[23] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2845) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N2191;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5750 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[24]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[23]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[0] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5673 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5750);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[7] = (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__37) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__38;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633 = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0] = !DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0] | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633) | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5625 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620) & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[7] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5625) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5700 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[7]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[7]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[30] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5700) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[7]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__56 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[7]);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5627 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5] & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[6] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5627) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5762 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[6]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[6]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[29] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5762);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[5] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5620 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5714 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[5]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[5]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[28] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5714);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5618 = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633 | DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[4] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5622) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5618;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5778 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[4]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[4]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[27] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5778);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[3] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5631 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5633;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5729 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[3]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[3]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[26] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5729);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[2] = DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5641 ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5680 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[2]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[2]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[25] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5680);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[1] = (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0]) ^ DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1];
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5743 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[1]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[1]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[24] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5743);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5694 = !((DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5682 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__50[0]) | (DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5767 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__34[0]));
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[23] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5701 & DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_N5694);
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__33 = a_sign ^ b_sign;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[31] = !(DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__29 | (!DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__33));
reg x_reg_0__I1518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__I1518_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[0];
	end
assign x[0] = x_reg_0__I1518_QOUT;
reg x_reg_1__I1519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__I1519_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[1];
	end
assign x[1] = x_reg_1__I1519_QOUT;
reg x_reg_2__I1520_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__I1520_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[2];
	end
assign x[2] = x_reg_2__I1520_QOUT;
reg x_reg_3__I1521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__I1521_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[3];
	end
assign x[3] = x_reg_3__I1521_QOUT;
reg x_reg_4__I1522_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__I1522_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[4];
	end
assign x[4] = x_reg_4__I1522_QOUT;
reg x_reg_5__I1523_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__I1523_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[5];
	end
assign x[5] = x_reg_5__I1523_QOUT;
reg x_reg_6__I1524_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__I1524_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[6];
	end
assign x[6] = x_reg_6__I1524_QOUT;
reg x_reg_7__I1525_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__I1525_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[7];
	end
assign x[7] = x_reg_7__I1525_QOUT;
reg x_reg_8__I1526_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__I1526_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[8];
	end
assign x[8] = x_reg_8__I1526_QOUT;
reg x_reg_9__I1527_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__I1527_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[9];
	end
assign x[9] = x_reg_9__I1527_QOUT;
reg x_reg_10__I1528_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__I1528_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[10];
	end
assign x[10] = x_reg_10__I1528_QOUT;
reg x_reg_11__I1529_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__I1529_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[11];
	end
assign x[11] = x_reg_11__I1529_QOUT;
reg x_reg_12__I1530_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__I1530_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[12];
	end
assign x[12] = x_reg_12__I1530_QOUT;
reg x_reg_13__I1531_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__I1531_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[13];
	end
assign x[13] = x_reg_13__I1531_QOUT;
reg x_reg_14__I1532_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__I1532_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[14];
	end
assign x[14] = x_reg_14__I1532_QOUT;
reg x_reg_15__I1533_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__I1533_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[15];
	end
assign x[15] = x_reg_15__I1533_QOUT;
reg x_reg_16__I1534_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__I1534_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[16];
	end
assign x[16] = x_reg_16__I1534_QOUT;
reg x_reg_17__I1535_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__I1535_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[17];
	end
assign x[17] = x_reg_17__I1535_QOUT;
reg x_reg_18__I1536_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__I1536_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[18];
	end
assign x[18] = x_reg_18__I1536_QOUT;
reg x_reg_19__I1537_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__I1537_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[19];
	end
assign x[19] = x_reg_19__I1537_QOUT;
reg x_reg_20__I1538_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__I1538_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[20];
	end
assign x[20] = x_reg_20__I1538_QOUT;
reg x_reg_21__I1539_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__I1539_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[21];
	end
assign x[21] = x_reg_21__I1539_QOUT;
reg x_reg_22__I1540_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__I1540_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[22];
	end
assign x[22] = x_reg_22__I1540_QOUT;
reg x_reg_23__I1541_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__I1541_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[23];
	end
assign x[23] = x_reg_23__I1541_QOUT;
reg x_reg_24__I1542_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__I1542_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[24];
	end
assign x[24] = x_reg_24__I1542_QOUT;
reg x_reg_25__I1543_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__I1543_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[25];
	end
assign x[25] = x_reg_25__I1543_QOUT;
reg x_reg_26__I1544_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__I1544_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[26];
	end
assign x[26] = x_reg_26__I1544_QOUT;
reg x_reg_27__I1545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__I1545_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[27];
	end
assign x[27] = x_reg_27__I1545_QOUT;
reg x_reg_28__I1546_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I1546_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[28];
	end
assign x[28] = x_reg_28__I1546_QOUT;
reg x_reg_29__I1547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__I1547_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[29];
	end
assign x[29] = x_reg_29__I1547_QOUT;
reg x_reg_30__I1548_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I1548_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[30];
	end
assign x[30] = x_reg_30__I1548_QOUT;
reg x_reg_31__I1549_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I1549_QOUT <= DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_x[31];
	end
assign x[31] = x_reg_31__I1549_QOUT;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[0] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[1] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[2] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[3] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[4] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[5] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[6] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[7] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[8] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[9] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[10] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[11] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[12] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[13] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[14] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[15] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[16] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[17] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[18] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[19] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[20] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[21] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__43[22] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[0] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[1] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[2] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[3] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[4] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[5] = 1'B0;
assign DFT_compute_cynw_cm_float_mul_E8_M23_1_inst_inst_cellmath__54[6] = 1'B0;
endmodule

/* CADENCE  vrH5SgvcrR8= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



