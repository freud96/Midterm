/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:23:54 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42;
wire [22:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68;
wire [0:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195;
wire [20:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197;
wire [32:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N623,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5570,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5577,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5578,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5600,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5607,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5614,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5616,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5623,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5629,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5641,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5657,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5664,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5754,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5866,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5869,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6087,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6179,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6189,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6197,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6224,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6256,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6257,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6258,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6292,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6299,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6310,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6347,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6356,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6359,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6381,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6396,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7360,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7365,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7438,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7450,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7555,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7570,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7929,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8158,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8179,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8197,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8221,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8222,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8252,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8292,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8294,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8360,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8361,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8364,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8382,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8384,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8405,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8425,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8429,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8436,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8442,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8445,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8452,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8459,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8465,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8471,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8474,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8485,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8502,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8537,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8539,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8555,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8579,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8586,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8607,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8612,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8614,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8616,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8632,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8657,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8735,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8860,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8868,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8900,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9059,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9087,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9093,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10425,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10430,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10436,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10438,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10442,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10443,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10445,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10449,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10450,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10452,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10459,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10465,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10470,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10475,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10476,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10500,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10558,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10593,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10600,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10613,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10617,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10629,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10650,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10661,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10674,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10765,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10797,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10807,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10860,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10861,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10889,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11701,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11735,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11738,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11753,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11760,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11765,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11791,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11806,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11807,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11813,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11826,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11830,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11839,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11851,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11863,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11866,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11869,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11872,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11890,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11904,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11911,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11931,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11937,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12021,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12030,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12047,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12059,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12087,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12093,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12118,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12129,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12145,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12165,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12189,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12193,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12194,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12221,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12224,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12229,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12240,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12256,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12269,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12271,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12347,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12351,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12356,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12361,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12364,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12365,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12367,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12381,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12384,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12392,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12396,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12406,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12423,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12429,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12431,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12432,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12438,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12447,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12470,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12472,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12474,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12475,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12476,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12478,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12490,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12491,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12501,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12502,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12520,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12527,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12532,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12537,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12567,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12578,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12579,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12582,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12593,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12599,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12602,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12603,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12605,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12606,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12607,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12610,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12613,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12614,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12617,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12619,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12622,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12625,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12626,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12628,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12629,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12630,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12632,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12633,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12635,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12637,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12639,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12640,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12642,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12644,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12645,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12647,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12648,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12649,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12651,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12652,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12653,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12654,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12656,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12658,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12659,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12661,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12664,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12665,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12670,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12683,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12688,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12696,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12702,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12706,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12707,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12712,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12714,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12716,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12723,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12732,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12736,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12738,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12740,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12745,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12747,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12751,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12758,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12765,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12766,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12772,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12773,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12778,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12779,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12784,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12785,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12791,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12793,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12797,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12803,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12804,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12818,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12819,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12821,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12825,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12826,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12827,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12828,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12830,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12832,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12833,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12834,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12836,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12837,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12840,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12842,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12843,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12844,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12848,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12849,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12850,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12853,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12854,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12856,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12857,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12859,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12860,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12861,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12862,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12863,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12864,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12867,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12868,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12870,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12871,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12873,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12874,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12875,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12876,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12877,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12879,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12880,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12882,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12884,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12886,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12888,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12889,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12891,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12892,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12894,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12896,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12897,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12900,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12901,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12902,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12903,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12906,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12907,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12908,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12909,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12910,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12913,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12916,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12917,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12918,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12919,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12920,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12922,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12923,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12924,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12925,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12926,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12927,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12930,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12933,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12934,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12935,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12939,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12941,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12943,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12952,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12953,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12958,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12959,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12969,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12971,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12977,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12983,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12993,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13004,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13010,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13018,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13022,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13047,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13058,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13060,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13066,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13077,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13080,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13083,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13092,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13093,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13095,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13098,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13109,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13116,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13126,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13129,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13131,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13138,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13142,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13149,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13157,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13158,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13165,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13168,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13169,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13177,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13180,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13186,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13189,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13197,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13204,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13214,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13222,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13224,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13228,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13229,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13233,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13243,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13252,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13253,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13258,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13264,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13266,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13291,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13299,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13305,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13310,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13329,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13333,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13337,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14940,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14944,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14950,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14956,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14960,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14963,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14966,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14970,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14985,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14988,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14992,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14994,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15001,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15008,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15011,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15026,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15028,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15035,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15038,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15044,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15054,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15078,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15081,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15084,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15086,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15097,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15100,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15105,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15107,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15110,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15113,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15123,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15127,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15129,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15135,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15137,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15143,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15144,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15147,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15161,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15166,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15170,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15175,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15177,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15184,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15187,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15192,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15199,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15201,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15210,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15215,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15241,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15257,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15265,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15311,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15325,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15327,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15338,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15348,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15352,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15354,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15366,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15369,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15372,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15379,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15412,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15416,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15419,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15420,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15424,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15428,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15429,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15435,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15441,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15448,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15453,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15457,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15463,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15466,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15483,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15485,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15487,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15490,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15510,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15524,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15539,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15543,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15559,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15560,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15573,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15580,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15589,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15590,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15594,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16294,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16298,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16332,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16334,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16343,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16357,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16362,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16376,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16390,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16393,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16401,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16403,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16409,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16411,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16417,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16486,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16488,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16489,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16492,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16493,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16497,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16500,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16506,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16508,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16509,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16514,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16515,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16516,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16519,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16522,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16534,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16535,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16537,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16541,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16542,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16545,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16546,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16548,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16551,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16553,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16554,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16556,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16557,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16561,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16562,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16564,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16566,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16643,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16646,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16662,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16663,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16667,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16685,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16691,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16693,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16703,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16704,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16719,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16727,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16741,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16742,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16746,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16754,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16762,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16775,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16776,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16783,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16789,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16790,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16794,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16795,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16809,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16810,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16814,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17141,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17198,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17202,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17205,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17207,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17211,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17213,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17217,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17220,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17223,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17227,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17230,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17234,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17237,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17244,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17247,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17251,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17256,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17263,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23226,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23240,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23255,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23303,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23307,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23314,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23324,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23367,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23375,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23399,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23407,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23415,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23421,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23433,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44729,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44981,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44986,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45000,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45015,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45016,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45019,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45020,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45023,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45031,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45033,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45036,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45040,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45043,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45045,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45050,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45052,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45055,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45064,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45065,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45068,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45070,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45072,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45115,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45117,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45118,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45119,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45132,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45146,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45148,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45150,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45152,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45155,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45200,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45206,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45208,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45238,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45239,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45242,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45245,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45246,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45249,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45252,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45254,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45259,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45262,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45267,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45270,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45273,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45276,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45279,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45282,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45283,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45286,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45290,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45293,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45296,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45297,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45300,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45341,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45342,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45345,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45350,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45353,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45355,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45358,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45368,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45371,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45377,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45380,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45383,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45386,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45389,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45391,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45394,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45397,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45400,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45439,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45446,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45451,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45454,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45460,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45464,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45473,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45494,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45504,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45525,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45526,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45530,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45547,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45549,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45552,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45569,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45572,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45575,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45576,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45581,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45583,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45584,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45587,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45592,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45595,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45598,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45601,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45604,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45608,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45611,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45612,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45615,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45618,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45620,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45621,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45624,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45631,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45668,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45677,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45679,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45684,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45687,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45692,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45695,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45698,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45700,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45705,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45708,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45711,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45713,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45718,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45720,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45721,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45724,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45756,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45763,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45771,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45774,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45780,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45786,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45792,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45799,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45805,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45811,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45817,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45823,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45829,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45835,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45841,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45847,
	DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45854;
wire N20585,N20596,N20746,N20748,N21279,N21282,N21470 
	,N21688,N22491,N22530,N22533,N22538,N22540,N22545,N22547 
	,N22552,N22554,N22559,N22561,N22566,N22575,N22580,N22583 
	,N22585,N22594,N22597,N22599,N22606,N22611,N22616,N22621 
	,N22624,N22626,N22636,N22641,N22648,N22651,N22672,N22682 
	,N22708,N22728,N22764,N22772,N22791,N22793,N22798,N22800 
	,N22812,N22814,N22816,N22826,N22828,N22830,N22833,N22835 
	,N22837,N22841,N22843,N22845,N22848,N22850,N22852,N22858 
	,N22860,N22864,N22866,N22868,N22871,N22873,N22875,N22881 
	,N22883,N22889,N22891,N22895,N22897,N22899,N22903,N22905 
	,N22907,N22910,N22919,N22973,N22978,N22985,N22992,N23039 
	,N23041,N23043,N23049,N23051,N23099,N23101,N23103,N23137 
	,N23601,N23606,N23608,N23613,N23615,N23620,N23628,N23630 
	,N23638,N23640,N23646,N23917,N23918,N23919,N23920,N23921 
	,N23922,N23923,N23924,N23925,N23926,N23927,N23928,N23929 
	;
EDFFHQX2 x_reg_20__retimed_I14257 (.Q(N23646), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15184), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I14255 (.Q(N23640), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I14254 (.Q(N23638), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15399), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14251 (.Q(N23630), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14250 (.Q(N23628), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14247 (.Q(N23620), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15019), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14245 (.Q(N23615), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14244 (.Q(N23613), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15487), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14242 (.Q(N23608), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14241 (.Q(N23606), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15113), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14239 (.Q(N23601), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15386), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14063 (.Q(N23137), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15008), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14046 (.Q(N23103), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15490), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14045 (.Q(N23101), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14044 (.Q(N23099), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14026 (.Q(N23051), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15428), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14025 (.Q(N23049), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15283), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14023 (.Q(N23043), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14022 (.Q(N23041), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14021 (.Q(N23039), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14003 (.Q(N22992), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I14000 (.Q(N22985), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15105), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13997 (.Q(N22978), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13995 (.Q(N22973), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15071), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13973 (.Q(N22919), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15448), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13969 (.Q(N22910), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15473), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13968 (.Q(N22907), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378), .E(bdw_enable), .CK(aclk));
fdeQ_A_bdw839185604_bdw x_reg_20__retimed_I13967 (.Q(N22905), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15524), .EN(bdw_enable), .CLK(aclk));
EDFFHQX1 x_reg_20__retimed_I13966 (.Q(N22903), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15376), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13965 (.Q(N22899), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15352), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13964 (.Q(N22897), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15550), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13963 (.Q(N22895), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15207), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13962 (.Q(N22891), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13961 (.Q(N22889), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15064), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13959 (.Q(N22883), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15152), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13958 (.Q(N22881), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13956 (.Q(N22875), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15044), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13955 (.Q(N22873), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13954 (.Q(N22871), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13953 (.Q(N22868), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15463), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13952 (.Q(N22866), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15265), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13951 (.Q(N22864), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15127), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13950 (.Q(N22860), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15175), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13949 (.Q(N22858), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14981), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13947 (.Q(N22852), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15539), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13946 (.Q(N22850), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15338), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13945 (.Q(N22848), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15195), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13944 (.Q(N22845), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15435), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13943 (.Q(N22843), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13942 (.Q(N22841), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15290), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13941 (.Q(N22837), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15241), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13940 (.Q(N22835), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15054), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13939 (.Q(N22833), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15573), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13938 (.Q(N22830), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15499), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13937 (.Q(N22828), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13936 (.Q(N22826), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15161), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13932 (.Q(N22816), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14956), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13931 (.Q(N22814), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15420), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13930 (.Q(N22812), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15278), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13925 (.Q(N22800), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15135), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13924 (.Q(N22798), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14992), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13922 (.Q(N22793), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15565), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13921 (.Q(N22791), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15409), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13914 (.Q(N22772), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15297), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13911 (.Q(N22764), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15589), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13906 (.Q(N22728), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15123), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13898 (.Q(N22708), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15441), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13887 (.Q(N22682), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15518), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13883 (.Q(N22672), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15226), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13874 (.Q(N22651), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15372), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13873 (.Q(N22648), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14966), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13870 (.Q(N22641), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15559), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13868 (.Q(N22636), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15100), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13864 (.Q(N22626), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13863 (.Q(N22624), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45835), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13862 (.Q(N22621), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15397), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13860 (.Q(N22616), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14991), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13858 (.Q(N22611), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14944), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13856 (.Q(N22606), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15170), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13853 (.Q(N22599), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13852 (.Q(N22597), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45811), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13851 (.Q(N22594), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15534), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13847 (.Q(N22585), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13846 (.Q(N22583), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45829), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13845 (.Q(N22580), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15192), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13843 (.Q(N22575), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15147), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13839 (.Q(N22566), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15325), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13837 (.Q(N22561), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13836 (.Q(N22559), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45847), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13834 (.Q(N22554), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13833 (.Q(N22552), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45841), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13831 (.Q(N22547), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13830 (.Q(N22545), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45817), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13828 (.Q(N22540), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13827 (.Q(N22538), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45823), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13825 (.Q(N22533), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15583), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13824 (.Q(N22530), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15348), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I13812 (.Q(N22491), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15419), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I13554 (.Q(N21688), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15081), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I13476 (.Q(N21470), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15143), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I13410 (.Q(N21282), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I13409 (.Q(N21279), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_27__retimed_I13216 (.Q(N20748), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_27__retimed_I13215 (.Q(N20746), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I13151 (.Q(N20596), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I14386 (.Y(N23917), .A(N20596));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14391 (.Y(N23922), .A(N23917));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14390 (.Y(N23921), .A(N23917));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14389 (.Y(N23920), .A(N23917));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14388 (.Y(N23919), .A(N23917));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14387 (.Y(N23918), .A(N23917));
EDFFHQX1 x_reg_22__retimed_I13146 (.Q(N20585), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163), .E(bdw_enable), .CK(aclk));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I14392 (.Y(N23923), .A(N20585));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14393 (.Y(N23924), .A(N23923));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I0 (.Y(bdw_enable), .A(astall));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45150), .A(a_exp[6]), .B(a_exp[5]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16362), .A(a_exp[4]), .B(a_exp[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328), .A(a_exp[2]), .B(a_exp[1]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16357), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I5 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45152), .A(a_exp[7]), .B(a_exp[0]), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16357));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I6 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45150), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45152));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I7 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I8 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16464), .A(a_sign), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19));
CLKINVX6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I9 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122), .A(a_man[2]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I10 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16403), .A(a_man[0]), .B(a_man[1]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I11 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16417), .A(a_man[12]), .B(a_man[11]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I12 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16386), .A(a_man[18]), .B(a_man[17]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I13 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16397), .A(a_man[16]), .B(a_man[15]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I14 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16407), .A(a_man[14]), .B(a_man[13]));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I15 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16409), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16417), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16386), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16397), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16407));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I16 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16403), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16409));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I17 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213), .A(a_man[22]), .B(a_man[21]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I18 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16411), .A(a_man[4]), .B(a_man[3]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I19 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16380), .A(a_man[10]), .B(a_man[9]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I20 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16390), .A(a_man[8]), .B(a_man[7]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I21 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16401), .A(a_man[6]), .B(a_man[5]));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I22 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16393), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16411), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16380), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16390), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16401));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I23 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16376), .A(a_man[20]), .B(a_man[19]));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I24 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16393), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16376));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I25 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I26 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19), .B(a_sign), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__24));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I27 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I28 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I29 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268), .A(a_exp[6]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I30 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289), .A(a_exp[5]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I31 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264), .A(a_exp[4]));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I32 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I33 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287), .A(a_exp[2]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I34 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280), .A(a_exp[1]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I35 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293), .A(a_exp[3]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I36 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I37 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I38 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267), .A(a_exp[7]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I39 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I40 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7267), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7291));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I41 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7270), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I42 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7271), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7270));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I43 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7271), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7268));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I44 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[6]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I45 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I46 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16334), .A(a_exp[3]), .B(a_exp[4]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I47 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16332), .A(a_exp[5]), .B(a_exp[6]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I48 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16324), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16328), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16334), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16332));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I49 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16294), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I50 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16298), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
OA22X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I51 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139), .A0(a_exp[7]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16324), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16294), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16298));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I52 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I53 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45122), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45159));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I54 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45118), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17163), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45119));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I55 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45146), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45132), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45118));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I56 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I57 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N594), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17178));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I58 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974), .A(a_exp[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284));
CLKXOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I59 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I60 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I61 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7293), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45763));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I62 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406), .A(a_man[22]), .B(a_man[21]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I63 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I64 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .A(a_man[21]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I65 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341), .A(a_man[20]), .B(a_man[22]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I66 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I67 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965), .A(a_man[19]), .B(a_man[21]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I68 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I69 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I70 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6156), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6341));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I71 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5663));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I72 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I73 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I74 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6172));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I75 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6283), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I76 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6212), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6017), .A(a_man[19]), .B(a_man[17]), .CI(a_man[22]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I77 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594), .A(a_man[20]), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6212));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I78 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I79 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201), .A(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I80 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5833), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5644), .A(a_man[21]), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I81 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5833), .B(a_man[16]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6017));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I82 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I83 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I84 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6154), .A(a_man[15]), .B(a_man[17]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I85 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870), .A(a_man[22]));
BUFX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I86 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I87 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6261), .A(a_man[14]), .B(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I88 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6317), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6131), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010), .B(a_man[20]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6261));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I89 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5644), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6154), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6317));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I90 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I91 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6377), .A(a_man[13]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I92 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5940), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .B(a_man[19]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6377));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I93 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5962), .A(a_man[15]), .B(a_man[17]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I94 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5962), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6131));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I95 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I96 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I97 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I98 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981), .A(a_man[20]));
BUFX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I99 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5621), .A(a_man[12]), .B(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I101 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5572), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6241), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637), .B(a_man[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5621));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6077), .A(a_man[14]), .B(a_man[16]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I103 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6077), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5749));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I105 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6108), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5915), .A(a_man[13]), .B(a_man[11]), .CI(a_man[16]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605), .A(a_man[19]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I107 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6051), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5866), .A(a_man[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6108), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I108 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6190), .A(a_man[13]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I109 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6051), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6190), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6241));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I110 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I111 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I112 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .A(a_man[18]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I113 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6218), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6025), .A(a_man[12]), .B(a_man[10]), .CI(a_man[15]));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .A(a_man[17]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I115 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5721), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I116 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5671), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6218), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5721));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6292), .A(a_man[12]), .B(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I118 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5671), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6292), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5866));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I120 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6326), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6141), .A(a_man[11]), .B(a_man[9]), .CI(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I121 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6166), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6025), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6326), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6413));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I122 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6348), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5915), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6166));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6115), .A(a_man[22]), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I128 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5840), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5651), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6115), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821), .A(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I130 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5581), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6248), .A(a_man[13]), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I131 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5732), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6421), .A(a_man[7]), .B(a_man[21]), .CI(a_man[9]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5922), .A(a_man[22]), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I133 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5949), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5759), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5732), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5922));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I134 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5787), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5600), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6141), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5581), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5949));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I135 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5840), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5787));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I136 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I137 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308), .A(a_man[14]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I138 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5680), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6357), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I139 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5849), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5656), .A(a_man[6]), .B(a_man[20]), .CI(a_man[8]));
CLKINVX6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929), .A(a_man[13]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I141 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6223), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929), .B(a_man[11]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I142 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6060), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5849), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6223), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6421));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I143 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6274), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6085), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6248), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5680), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6060));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I144 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5651), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5600));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I146 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565), .A(a_man[12]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I148 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6336), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6148), .A(a_man[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I149 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5793), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6336));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I150 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5956), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5769), .A(a_man[5]), .B(a_man[19]), .CI(a_man[7]));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I151 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6174), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5956), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5656));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I152 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5895), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5793), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6357), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6174));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I153 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5895), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5759), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6085));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041), .A(a_man[11]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I156 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5589), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6255), .A(a_man[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I157 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5903), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5589));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I158 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6070), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5883), .A(a_man[4]), .B(a_man[18]), .CI(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I159 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6281), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6092), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6070), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6148), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5769));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I160 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6388), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6197), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5903), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5609), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6281));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I161 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6388), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5876), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5700));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I165 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902));
CLKINVX6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662), .A(a_man[10]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I167 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5686), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6370), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I168 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6009), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5824), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5686), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I169 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6289), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6101), .A(a_man[2]), .B(a_man[16]), .CI(a_man[4]));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I170 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6123), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6289));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155), .A(a_man[9]));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I172 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5803), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5616), .A(a_man[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I173 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6182), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5988), .A(a_man[3]), .B(a_man[17]), .CI(a_man[5]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I174 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5635), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6310), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5803), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6370), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5988));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I175 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5627), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5824), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6123), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5635));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I176 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6396), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6182), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6255), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5883));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I177 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6004), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6009), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6396));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I178 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5627), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6092), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5817));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I179 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6004), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5983), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6197));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I183 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6133), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I184 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6243), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6054), .A(a_man[14]), .B(a_man[21]), .CI(a_man[0]));
CLKINVX6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263), .A(a_man[7]));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I186 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5752), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5574), .A(a_man[5]), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I187 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6343), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6133), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6243), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5752));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I188 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5646), .A(a_man[22]), .B(a_man[15]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I189 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6407), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6214), .A(a_man[3]), .B(a_man[1]), .CI(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I190 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6233), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6407));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6318), .A(a_man[22]), .B(a_man[15]));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778), .A(a_man[8]));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I193 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5910), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I194 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5857), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5664), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6318), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6214), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5717));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I195 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5734), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6343), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6045), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5857));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I196 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5742), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5910), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6101), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5616));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I197 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6117), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5933), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6233), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5742));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I198 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6310), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5734), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5923));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I199 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6117), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6204), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6303));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I200 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5601), .A(a_man[20]), .B(a_man[13]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I205 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5867), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5674), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821));
CLKINVX8 DFT_compute_cynw_cm_float_cos_E8_M23_1_I206 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927), .A(a_man[6]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I207 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6351), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6167), .A(a_man[4]), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I208 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5595), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5601), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5867), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6351));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I209 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5966), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6054), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5942), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5574));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I210 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6224), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6036), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6157), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5966));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I211 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6224), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5566), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5560));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I213 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6087), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5896), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5819), .A(a_man[19]), .B(a_man[12]));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378), .A(a_man[5]));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I216 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5702), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6391), .A(a_man[3]), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I217 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5695), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6087), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5819), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5702));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I218 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6276), .A(a_man[20]), .B(a_man[13]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I219 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6079), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6276), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5674), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6167));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I220 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5852), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5659), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6267), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5695), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6079));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I221 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5852), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5664), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6036));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611));
NAND2X6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I224 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5925), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5736), .A(a_man[11]), .B(a_man[18]), .CI(a_man[2]));
CLKINVX6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I225 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995), .A(a_man[4]));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I226 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6305), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I227 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5810), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5623), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5925), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6305));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6152), .A(a_man[17]), .B(a_man[10]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I229 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5562), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6225), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5981));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I230 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5918), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6152), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5562));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716), .A(a_man[3]));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I232 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6038), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I233 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6297), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6110), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6038), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6120), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5736));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I234 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5958), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5623), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5918), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6297));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5629), .A(a_man[19]), .B(a_man[12]));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I236 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6192), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5629), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6391));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I237 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6337), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6192), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6381));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I238 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5958), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5891), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6150));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I239 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6337), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5780), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5659));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260));
NOR2X6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6389), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071));
CLKINVX8 DFT_compute_cynw_cm_float_cos_E8_M23_1_I246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723), .A(a_man[1]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I247 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5894), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723), .B(a_man[6]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I248 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5786), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5598), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I249 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5754), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5575), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5894), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5598), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I250 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5669), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6347), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I251 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6272), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6084), .A(a_man[0]), .B(a_man[7]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I252 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6163), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5971), .A(a_man[1]), .B(a_man[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I253 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6134), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6272), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5786), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5971));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I254 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5754), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6347), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5945));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5980), .A(a_man[9]), .B(a_man[2]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I256 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5570), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6237), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5980));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I257 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740), .A(a_man[0]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I258 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6050), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5862), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I259 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5648), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6320), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5669), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6163), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5862));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I260 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6237), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6134), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6320));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I261 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6171), .A(a_man[9]), .B(a_man[2]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I262 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6056), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5872), .A(a_man[3]), .B(a_man[10]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I263 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6314), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6171), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5872));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I264 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5937), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5748), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I265 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6021), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5837), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5748), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6050), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5570));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I266 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6127), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5837), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5648));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5848), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I269 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5578), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6246), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122), .B(a_man[11]), .CI(a_man[4]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I270 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6207), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6013), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6246));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I271 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5828), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I272 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6409), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5640), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5937), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6314));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I273 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6021), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6013), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6215));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I274 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5947), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5755), .A(a_man[5]), .B(a_man[12]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I275 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6096), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5906), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5578), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5821), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5755));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I276 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5713), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I277 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5911), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5718), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6399), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6207));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I278 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5906), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6409), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5718));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5577));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5848), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I283 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5869), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5675), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6308), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6002), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I285 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6244), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I286 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5699), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5869), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6055));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I287 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6244), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6084), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5575));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6181), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5815), .A(a_man[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I291 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6352), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6169), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5929), .B(a_man[4]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I292 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5815), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6352), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5675));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I293 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6279), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I294 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5976), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5789), .A(a_man[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5565), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I295 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5604), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6278), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041), .B(a_man[2]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I296 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5604), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I297 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6169), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5976), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I300 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5703), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155), .B(a_man[0]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I301 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6088), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662), .B(a_man[1]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I302 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5899), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I303 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6278), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6088), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I304 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I305 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6315), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I306 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6200), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I307 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6200), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6392), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I309 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5820), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5631), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I310 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5820), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6007));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I311 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6173), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I312 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I313 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5563), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I318 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I320 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6339), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5634), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6188), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6309));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I321 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6288));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I322 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6203), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5615), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5802));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I323 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6227), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6395), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5823), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6203));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I324 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5898), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5563), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6339), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6227));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I325 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I326 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5739), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5716));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5901), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5987), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6180));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5944), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5898), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5901), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5706));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I330 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5631));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6020), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I333 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6091), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6369), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5685));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I334 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5607), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5882), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6069));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5835), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6091), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5792), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5607));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5771), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5944), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6020), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5835));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5982), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6254), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5588));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6356), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5767), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5954));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I339 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5856), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5982), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6356));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6239), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5677), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6173), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5771), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5856));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I341 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6147), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6335));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6247), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5847));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6130), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5580), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5875), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6247));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5758), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6033), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6222));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6419), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5730));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6015), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6325), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5758), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6138));
OA21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6137), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6130), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6015));
OAI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5704), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6211), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6315), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6239), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6137));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6090), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6114));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I350 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6100), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6279), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5704), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6090));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I351 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6301), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5626));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I352 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5979), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5813), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6001));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I353 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5989), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6170), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5606), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5979));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6181), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6100), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5989));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6194), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6385));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5871), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5698), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5893));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5658), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6058), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6355), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5871));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6082), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6270));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I359 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5597), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5785));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6420), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6245), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5946), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5757));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5731), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5658), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6420));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I363 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5776), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6041));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I364 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6374), .A(a_man[16]), .B(a_man[9]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I365 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6259), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45245), .A(a_man[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6122), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6263));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I366 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6030), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5843), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5776), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6374), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6259));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I367 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5960), .A(a_man[17]), .B(a_man[10]));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I368 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6416), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5960), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6225), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5854));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I369 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5591), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6256), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5727), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6030), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6416));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I370 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5998), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5591), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5774));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6105), .A(a_man[15]), .B(a_man[8]));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I373 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45282), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5723), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5662));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I374 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6144), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6105), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45282));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I375 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45296), .A(a_man[16]), .B(a_man[9]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I376 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5653), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45296), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45273), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45245));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I377 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6072), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5885), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5843), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6144), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5653));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I378 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6072), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6110), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6256));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I379 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I381 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5839), .A(a_man[14]), .B(a_man[7]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I382 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45300), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6089), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6354), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5839));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I383 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45242), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5705), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5637), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6155));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I384 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6322), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6136), .A(a_man[6]), .B(a_man[13]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5995));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I385 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5650), .A(a_man[14]), .B(a_man[7]));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I386 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45238), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5740));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I387 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45270), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6322), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5650), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45290));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I388 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45246), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45286), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45242), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45270));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I389 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45254), .A(a_man[15]), .B(a_man[8]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I390 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45262), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45249), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45254), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45238), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45267));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I391 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5687), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45259), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45300), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45276), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45262));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I392 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45246), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45239), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45259));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I393 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5687), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6220), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5885));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I398 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45252), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6285), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5778), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5605), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6010));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I399 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45279), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6201), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6136));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I400 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45283), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45293), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45252), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45279));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I401 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45283), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45249), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45297));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I403 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6290), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6285), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5713), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6096));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I404 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5683), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6290), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5618));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I406 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I407 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5799), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6103));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346));
OAI2BB1X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6135), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5969), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6162));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5649), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6346), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5668));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I414 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6135), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5838), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5649));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5861), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6049));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6236));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5970), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6164), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5970));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5745), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5935));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I420 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6126), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6313));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I421 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I422 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5827));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6012), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6206));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6401), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5712), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6401));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I428 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6398), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5710));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I429 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6095));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6284), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5611));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5798), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5984));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5952), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I434 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6143), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5952));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6363));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5682), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5878));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I437 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I438 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6250));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5582), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5763));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6380), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5694), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6380));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I442 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5950), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6142));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6330), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5652));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I445 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I446 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5842), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6029));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6414), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6219));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5932), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6124), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5932));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I450 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5916));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6296));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5808));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6191));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6359), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5679), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6359));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6379), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5693));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5889), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6078));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5594), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6266));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5965), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5779));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5914), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5691), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6107), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5914));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5641), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5887), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5691));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5773), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5829), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5641));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6196), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5959), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5773));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6389), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6196));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5610), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6283), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5834), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6019));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5851), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649), .S0(a_exp[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6406));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5681), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6199));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5619), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6387), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6006));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5619), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6213));
OA21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5681), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6358));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651), .S0(a_exp[0]));
CLKINVX8 DFT_compute_cynw_cm_float_cos_E8_M23_1_I481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I482 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I483 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5657), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I486 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5657));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I487 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5890), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5850), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5890));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6265), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6228));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6366), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6342));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6003), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I493 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6386));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5768));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5936), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6195), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5747));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5919), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6176), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5726));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6258), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5902), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6158), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5707));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5816), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5590), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6258));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6003), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5816));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6053), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6242));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I503 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I504 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6415), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5934), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6415));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5744), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5917), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5855));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5934), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5744), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645), .S0(a_exp[0]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6319), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5645));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5941), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6132));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5751));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6217));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I514 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5770), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5573));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6189), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5957), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6026), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5770));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6189));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6230), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6376), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6230));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I519 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5741), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5738));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I520 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
CLKMX2X6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7280), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7287));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457));
XOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7264), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7284));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7528));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I529 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44974), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7289));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N650), .S0(a_exp[0]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N652), .B(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071), .A(a_exp[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45061));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I535 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45051));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45019), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45064), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45045));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45046));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45043), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45032));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45065), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45016), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45043), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45031), .A(a_exp[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45065));
NOR3X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I542 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45015), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45070), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45031));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I543 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45067));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I544 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45050), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45040), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45033), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45025), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45068));
NOR3X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I547 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45052), .A(a_exp[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45050), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45033));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45072), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45023));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45020), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5750));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45036), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45072), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45020), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45071));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45055), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45052), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45036));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45015), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45055));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I554 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I555 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512));
NAND3X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44981), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I557 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I558 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N706), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7447));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I562 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I563 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6275), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5603));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I564 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45473), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5897));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45454), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45456), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I570 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640), .S0(a_exp[0]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I571 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6168), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6350));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I572 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I573 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6022), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5711), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6183), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I576 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5666), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5711));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6345), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6094), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6311));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I578 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5666), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6345), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5788), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5974));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I581 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5968), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6235));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5608));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5968), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5784), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5818));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6299), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I588 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5975), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I589 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6184));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6102));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6302), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6071), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5991), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5884));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I592 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5628), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6299), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6277), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6304));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I595 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6277), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636), .S0(a_exp[0]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6390), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5701));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I600 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5576), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6300), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6408), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6300));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I603 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45439), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5814), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6046));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I604 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45439), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I605 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6005), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6198));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5955), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6232), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45460), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5955));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6334), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6044));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45460), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45451), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5865));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I610 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I611 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I612 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I613 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N649), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N648), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I614 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7478), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7333), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5868));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6140));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6063), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6327), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6063));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5583), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5825));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6234), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6048), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6240));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N645), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7365), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N646), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I623 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7365), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I624 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I625 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7423), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7428), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7423), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7348));
XOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7391));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I630 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7570), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N640), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N639), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N642), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N641), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I635 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5926));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5977), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I638 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5977), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6018), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5753), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5729), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6018));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6404), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5781));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I642 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5804));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I643 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6208), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6014));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I644 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5924), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5688), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5617), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6371));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I645 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6116), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6208), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5924));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I646 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5729), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6418), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I647 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N637), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7424), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7533), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N644), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N643), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I653 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7565), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I654 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I655 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7366), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I656 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7366), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N696), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7549));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7344), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7454), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I663 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7373), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7486), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I664 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7477), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7457), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7404), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7477));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7404));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N698));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12808), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11882), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7402), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7503), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7416));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N705), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I679 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7346), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7394), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7559), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7559));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7401), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7508), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I687 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7411), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7378));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7450), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7450));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23276));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7332), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7547), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7522), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7480), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7480));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N701), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7354), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7388), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7325));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I703 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7337), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N702), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7337));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N702), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I710 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7949));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8780));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I714 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I717 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I719 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8231));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I720 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I721 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8161), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9050), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8161));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[21]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I729 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8122));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I732 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8703));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9127));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I738 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8782));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I744 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I745 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I746 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8407));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8330), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8985));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I755 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I757 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8536));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I765 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8375), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[19]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I766 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9026));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I767 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I768 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I769 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I770 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I771 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I772 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I773 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I777 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I778 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I779 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I780 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I781 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I782 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I783 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I786 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I787 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I789 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8804), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I790 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I791 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I794 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I795 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I796 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7961), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I800 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9059), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7961));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I801 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8345), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9059));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I802 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8345), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8605));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I14394 (.Y(N23925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I14395 (.Y(N23926), .A(N23925));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I803 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I804 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12838));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I805 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7432), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7543), .S0(a_exp[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I806 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7444), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I807 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7535), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7512), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7535));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7513));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I810 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N699), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I811 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7499), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7532), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7437), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7467), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7370), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I816 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7370));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I817 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N700), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I818 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[16]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I819 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11849), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I822 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11849), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I823 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8554));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I827 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9075));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I834 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8478), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I838 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8670), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8106), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8670));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I841 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I842 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I843 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I844 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I845 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I846 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I847 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I848 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I849 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8920), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I850 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8223), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8106), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8920));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I851 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8743), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8478), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8223));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I855 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8828), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I858 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I859 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I860 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8624), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I861 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8743), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8624));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I14396 (.Y(N23927), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I14397 (.Y(N23928), .A(N23927));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I862 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I863 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I864 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12225), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12869));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I865 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[41]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[40]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12225));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9028));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8210), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I870 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8037));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I871 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I872 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I873 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I874 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I875 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8323));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8853));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I879 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I881 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I882 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8677));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I883 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8192), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I884 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8252), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8192));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8748));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8252), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I892 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7934), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8909), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I893 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8306), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I894 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8024), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I899 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8151), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I900 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9046));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I901 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I902 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I903 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I904 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7888));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7907));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I908 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8465), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8151), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8024), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8465));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I910 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8210), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8040), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7934), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8728));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I912 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I913 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8652), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I914 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8389), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8676));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I915 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8831), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I916 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I917 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7968), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I918 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8652), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7968));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I919 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8898), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8774));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I920 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I921 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I927 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8080), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9067), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I928 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N761), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8898), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8349), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8080));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I929 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N761));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I930 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I931 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12932));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I932 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12719));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I933 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I934 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12261), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12898));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I935 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7460), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7536), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I936 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6226), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5561));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I937 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I938 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5672));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I939 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5846), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5624));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6032), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N635), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7321), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7475), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7546), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7460), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7566), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45504));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I947 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45771), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I949 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45771));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7426), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I951 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5853), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6037));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I952 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I953 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6307), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6333), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6146), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I955 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I956 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I957 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I958 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7510), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7489), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I959 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7438), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7349), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7510), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I960 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7438));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I962 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[10]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I963 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12835), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I965 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12835), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I966 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I967 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8678), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I968 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8164));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I969 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I970 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8083));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I971 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8875));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I975 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8597), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8749), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I976 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8058), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I977 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8977));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8396), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8506));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I983 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I984 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8635));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I985 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8058), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8484));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I986 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8597), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8325));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I987 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12994));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I989 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12916), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12581), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12261), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13146));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I990 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[40]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[39]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12363), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12916));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I991 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[40]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[22]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[40]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I992 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I993 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8806));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I994 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8462));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I995 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9111), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I996 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I997 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I998 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I999 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9053), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9111), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8919));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1000 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8392), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8195), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1002 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7995));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8584), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1005 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8584));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1006 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8821), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8759), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8936), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8992), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8821));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9053), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8759));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11913), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1013 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1014 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12658), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12866));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1015 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7368));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5737), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6338), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5660));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1017 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5737), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1018 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N633), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632), .S0(a_exp[0]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1019 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7463), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1020 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1021 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7436), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1022 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7379), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7492), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7456), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1023 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7379));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1025 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7833), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N693), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23275));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7568), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1027 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5961), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6151));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1028 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1029 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1030 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6394));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1031 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5733), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5602), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382));
XNOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5766), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5733));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1033 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5587), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6382), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6118));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5559));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5766), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5587), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N632), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7408), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1038 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7563), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7376), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7400), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7324));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273));
XOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1044 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12863), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1045 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12863), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1046 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1047 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1048 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11894), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12962));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1049 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12422), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12066), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12658), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11894));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1050 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1051 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13186), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13023));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12298), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12931));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1055 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12127), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13186), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12298), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13297));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8186), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1058 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8657), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8186), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8783), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8657));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1061 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1062 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1063 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8950), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9010));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1065 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1066 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7977), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8444));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1067 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9076), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8950), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7977));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8905), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8783), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9076));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1069 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8351));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8419));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8085), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8248), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1074 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8085), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8248));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1075 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8353));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1076 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1077 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13057));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1078 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13130), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12772), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12127), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12785), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12066));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1079 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[39]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[38]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12581), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12422), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13130));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1080 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[39]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[21]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[39]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1081 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1082 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8654));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1083 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8502), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1084 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1085 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8502), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8074));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1086 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1087 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8286));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1088 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1091 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8057));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1092 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8925));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1093 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8767), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1094 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8844), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8138), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8767));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1095 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8158), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8844));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1096 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8701));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7967));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1101 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9123));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8333));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1105 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8454));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9142), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8158), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8411));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1107 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1108 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1109 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1110 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1111 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12895));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1112 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5775));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6257), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6251), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6257));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6065), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5772));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6068), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N631), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1118 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7351), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7387), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1120 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7387), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7322), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1121 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7524), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7343), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1122 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7524));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N691), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6260));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6368), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6179), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5777));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1128 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6368), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6179), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1130 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7551), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7453), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7544), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7331), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7521), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7469), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7414), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7544), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7469));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1135 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7812), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N690));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1136 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[6]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1137 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12892), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1138 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12892), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1139 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8483));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1142 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1144 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8579), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1146 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8575));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7984), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8857), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7984), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1149 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7895), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1152 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8000), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8857), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7895));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1153 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8579), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8000));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8773));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8169), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8519));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1158 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9101));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8123), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8169), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8425));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1165 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8370));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8904));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1168 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1169 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8618));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8537), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8273));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8377), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8537));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8377));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1173 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1175 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7918), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1176 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1177 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8448), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1178 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8448));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8513));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8711), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8338));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1183 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8705));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8399));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1187 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8146));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1188 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958));
AND4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7918), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8026), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8711), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8562));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1193 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12078), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13188));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1195 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11813), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12078));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1196 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1197 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12439), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13122));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1198 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11905), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13196), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11813), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12439), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11750));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1200 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12816), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13088));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11931), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12990));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8798), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1206 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9089), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1207 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8798), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9089));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1208 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8259), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1209 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1210 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8259), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8522));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1211 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8317), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8471), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8739));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8173), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8317), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1216 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8846), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1217 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1218 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1219 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7989), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1221 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7989), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8586), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8101), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8218));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1224 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7937), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1225 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8586), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7937));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1226 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8173), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8432));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13257));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1229 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1230 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12960));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1232 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11721), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12331), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11688));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1233 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12551), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12186), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11931), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11721));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1234 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12477), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13151));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1236 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13222), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13053));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11978), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12721), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12928));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6075), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5886));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6075), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6286));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7495), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1247 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7398), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7487), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7531), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7466), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1249 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7412), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7357), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7487), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1250 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7412));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1251 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6186), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6373));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1254 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6393), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1256 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6393), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1257 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6306), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1258 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45756), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6321));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5614), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5836), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6111));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6035));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1261 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5801), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5614), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1262 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1263 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7441), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1264 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7341), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7434), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7473), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7410), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1266 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7557), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7434), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7355));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N688));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12926), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1272 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13219));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1274 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13304), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12115));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1275 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13168), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12800), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12477), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13222), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13304));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1276 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13265), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13168), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13105), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12186));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1277 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12635), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13196), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12551), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13265));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1278 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[38]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[37]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11905), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12635));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1279 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[38]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[20]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[38]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8112));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1283 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8671), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9066));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8633));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8571), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8528), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8571));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1291 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8744), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8921));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1292 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8671), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8744));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1293 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1294 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8053), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7884), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1295 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8107), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8053), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8107));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1300 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8625), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8867), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7903), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8590));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[14]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1302 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1303 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1304 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[15]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1305 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10403), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[13]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1309 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10403), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10442), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10576));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1310 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1311 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10851));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1312 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[12]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10457), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10855), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1318 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45499));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10920), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1320 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10666), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10529), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10493), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10855), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10920));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1321 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10425), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10457), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10666));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1322 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1323 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1324 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10778), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1325 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1326 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1327 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10737), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10778), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10992), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10592));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1329 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10737), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10809), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10529));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10838), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10892), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1333 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1334 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10554), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10401), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10838), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10892), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10936));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[9]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10653), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1339 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1341 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10988), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10842), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10433), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10410), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10573));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1342 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10819), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10710), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10653), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10988));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1343 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10610), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10554), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10819));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10933), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10441));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10716), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10586));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10939), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10939));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1350 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1351 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10793), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11023));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1352 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1353 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10447), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10568), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10435));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10774));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11029), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10786), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10917), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1359 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10515), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10786), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10917));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[8]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1363 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1364 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[7]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1365 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44729), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1366 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44729));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1367 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1368 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10782), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10656), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10981), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10763), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11008));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1369 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10629), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10515), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10513), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10782));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1370 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10629), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10401), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10684));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10649), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1374 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1375 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10675), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10543), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10649), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10640), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10497));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10702), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
CLKINVX6 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1377 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1378 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10862), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1379 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10870), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10655), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1381 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1382 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10566), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10417), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10655), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11005));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1383 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10946), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10702), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10862), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10566));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1384 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10427), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10675), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10946));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1385 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10427), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10842), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10492));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1386 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1387 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1388 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10424), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1389 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10848), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1390 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1392 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10832), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10424), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10848), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10724));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10996), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10583), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10715), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1397 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10443), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10935), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10583), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11026), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10715));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1398 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10480), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10443), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10417));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1399 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10601), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10455), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10543), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10832), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10480));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1400 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10601), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10656), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10923));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11010), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1404 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10598), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1406 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10717), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10776), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10598));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1407 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10726), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1410 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10960), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10824), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10726), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10512), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10739));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10928), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10439), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1413 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10686), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10928), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10439));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1414 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11000), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10853), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10960), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10686), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10935));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1415 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10748), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10621), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10717), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11000));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1416 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10748), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10808), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10455));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1420 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1421 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5806), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5993));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1422 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5830), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5978));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5639), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6353));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6099), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5909), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N627), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7385), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1428 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7541), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7318), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1429 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7375), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7419), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7501), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7375), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7555));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N687));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1434 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10452), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10469), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1437 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1438 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10925), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10454), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10469), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10792));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1439 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10613), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10483), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10452), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10925));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10860), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10926), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1442 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1443 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10581), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10860), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10926), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10833));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1444 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10881), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10740), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10581), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10557), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10824));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1445 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10644), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10505), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10613), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10591), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10881));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1446 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10644), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10974), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10621));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10807), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1450 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1451 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10893), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11019), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10807), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10528));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6291), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5620));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6403), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6210), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6106));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6403), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6210), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7516), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7329), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7362), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7516), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7320), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7552), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7448), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7320), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7498));
CLKXOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23277), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N686));
CLKINVX8 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10597), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6412), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6104));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6097), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N625), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7529), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7462), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7496), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7392), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7518), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7446));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23273));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[1]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10805), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1479 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10544), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10597), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10805));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1480 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10845), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10709), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10944), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10544));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10660), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1482 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1483 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10593), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1486 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10811), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45621), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10660), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10593), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10569));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1487 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10495), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10811), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10784), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10432));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1488 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10530), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10470), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10845), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10495));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1489 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10853), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10530), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10505));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1493 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6410), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5720));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6216));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5928), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6083));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6023));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6040), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6153), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6271), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5844));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5832), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5564), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6040));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N623), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5643), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N5832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N6400));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1503 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7360), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N624), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N623), .S0(a_exp[0]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1504 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7360), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7472), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[1]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7506), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7372), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7407), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7468));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7506), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7443), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7390), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7335), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7464), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7390));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N684), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23278));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[0]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10551));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1512 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45631), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10556), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10673));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10476), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1514 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10458), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45584), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10476), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45631), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10750));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10890), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
ADDHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1519 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10558), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10890), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10609));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1520 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45595), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45581), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11016), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10913), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10558));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10445), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10541), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45774), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10877));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10671), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1527 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10825), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10671), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10902));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1528 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45624), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45608), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10827), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10445), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10825));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1529 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10729), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45612), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45595), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45624));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1530 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10759), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10635), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10709), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10458), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10729));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1531 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10740), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10759), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11028));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10731), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1535 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1536 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45583), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10731), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10722), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10645));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10987), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10922));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10620), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1539 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10787), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10661), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10987), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10620));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1541 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45611), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45598), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10787), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10560), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10408));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1542 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45587), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45572), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45583), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45611));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1543 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11013), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45621), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45584), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45587));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1544 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11013), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10991), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10635));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1547 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10633), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10461), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1550 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10434), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10927), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10451), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10633), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10461));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11001), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10972), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10823));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1554 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10727));
ADDHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1555 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10398), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10895), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10972), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10706));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1556 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10711), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10582), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10907), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10398));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1557 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45575), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10883), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10688), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10711));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1558 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45615), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45601), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45581), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45608), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45575));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1559 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45615), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45612), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45576));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1562 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1563 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1564 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10679), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10548), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10683), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10804));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10718), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10814), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10542));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
ADDHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1569 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10918), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10775), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10428), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10538));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1570 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10951), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10815), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10718), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10814), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10918));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1571 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45620), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10661), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10951));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1572 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45604), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45569), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45620));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1573 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45604), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45572), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45601));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1576 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1578 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10625), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1581 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10865), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1583 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10500), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10865), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10970));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1584 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10617), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10477), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10533), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10625), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10500));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10889), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10894), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1588 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10449), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10889), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10430), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10894));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1589 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11006), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10617), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10940));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10444), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1592 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10839), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10994), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10444), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10775));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10516), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3809));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10619), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1595 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10967), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10516), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10619));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10797), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1599 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10801), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10670), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10416));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1600 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10720), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10596), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10797), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10670));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10590));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1603 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10574), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10423), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10547), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10708), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10801));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1604 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10487), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10720), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10449), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10423));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1605 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11006), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10700), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10980));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10973));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1607 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10604), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10895), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10637), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10574));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1608 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10872), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10732), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10839), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10548), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10815));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1609 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10487), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10462), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10732));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1610 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10636), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10582), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10927), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10604));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1611 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10847), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10872), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10496));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1612 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1613 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1614 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10883), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10534));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10436), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10517), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10979), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1623 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10764), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10517), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10979), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10882));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1624 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10885), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10743), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10829), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10764));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1625 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10596), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10885), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10858));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10540), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10788), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10600), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11027));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1630 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10930), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10693), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10600));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1631 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10412), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10788), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10930));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1632 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10412), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10477), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10743));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10450), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10962), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1635 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10676), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10765), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1638 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10817), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10681), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10676), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10765));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1639 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11020), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10422), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10817));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1642 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44730));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1643 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10415), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10634), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1644 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10734), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10415));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1645 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10585), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10438), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10523), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10699), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10734));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1646 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11020), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10789), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10438));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1647 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10639), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10585), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10909));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11015), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10431));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1653 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10898), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11037));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1654 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1655 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10465), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10898), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10605), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10681));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1656 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10606), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10874), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10465));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10510), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10867));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10852), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1663 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10627), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10749), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10852));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1664 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10510), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10627));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10481), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10810));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10587), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418));
ADDHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1668 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10587));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10840));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10861), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10878));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10790), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021));
OAI2BB2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10982), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11021), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10861), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10790));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10816), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10984), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10489), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10982), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10414));
OAI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10584), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10692), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10816), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10756), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10399));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955));
AOI2BB2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10966), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10550), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10955), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10584), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10969));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10525));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1679 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10650), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10618), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10966), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10479));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10663), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10714));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10950), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10888), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10650), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10745));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10850), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10561));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10691), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11033));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10871), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11035), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10803), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10672));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10472), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11015), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10950), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10871));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10536), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10511));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1687 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10975), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10450), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10472), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10942));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10975));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11036), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10626));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10540), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10747), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11036));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10674), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11017));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10761));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10453), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10674), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10945));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10906), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10798));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10937), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10484));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10623), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10518));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10658), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10903));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1703 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10406), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10667));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10768));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10891));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11038), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10728));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1710 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10864), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10579));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10758), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10705));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10900), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10958));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1714 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10880));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10575), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467));
OA21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10701), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10575));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1717 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10697), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11014), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10837), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10697));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1719 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10519), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11014));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1720 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10690), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10828), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1721 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10723), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__115__W1[0]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10836));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10941));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10478), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10562), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10502), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10413));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1729 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10968), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11034), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10887));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10859), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10802), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10721));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1732 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10873), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10440), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10932));
OA21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10545), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11018), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10873));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10978), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10678), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10698), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10545));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10659), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10486), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10978));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10961), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10785), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10659));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[32]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10723), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10961));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1738 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13228), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12514), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[32]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13228));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12514));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23314), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23314));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1744 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1745 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13019));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1746 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7963), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8238), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7963), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9061), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8281), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1755 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8076), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7922), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8076), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1757 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8756));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8941), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8868), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8868), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8607), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8941), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8504));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1765 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8200), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8607));
AND3X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1766 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8238), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9061), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8200));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1767 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1768 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13325));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1769 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1770 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12850), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13120));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1771 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12373), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11971), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12992), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12850));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1772 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12246), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11873), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13010), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12373), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1773 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13262), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13085));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8264), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1777 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8415), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8722));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1778 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8108), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8264), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8415));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1779 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1780 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8203), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1781 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8849), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9070), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8203));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1782 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1783 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7885), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8803), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8849), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7885));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1786 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1787 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9055), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1789 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8972), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8673));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1790 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9096), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8803), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8972));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1791 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8108), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9096));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12651), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11712));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1794 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1795 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12510), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13184));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1796 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13207), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12834), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13262), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12651), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12510));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11738), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13288));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1800 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12369), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12987));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1801 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11751), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1802 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11759), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11738), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12369), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11751));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1803 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13076), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12726), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11759), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1804 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1805 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11680));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1806 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8751), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1807 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8751), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8651));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1810 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8981), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7946));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1811 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9005), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8440));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8551), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7909), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9132), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1816 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9003));
NAND4BBXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1817 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8877), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219), .BN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1818 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7943));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1819 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8060), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8809), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1822 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8595));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1823 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8327), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8382), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8060), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8327));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1827 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8287), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8382));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N753), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8014), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8551), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8287));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N753));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11776));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12006), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13051));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1834 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12620), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13028), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12290), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12006));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12009), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N3808));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1838 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12751), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12957));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1841 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1842 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1843 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1844 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13251));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1845 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11885), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13177), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12751), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12145));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1846 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12283), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11911), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12620), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11885), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13046));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1847 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12159), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12283), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12008), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12726));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1848 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12950), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12611), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11873), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13076), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12159));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1849 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12337), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12888), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12246), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12950));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1850 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[37]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[36]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13204), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12275), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12337));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1851 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[37]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[19]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[37]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8508), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1855 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8013), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8013), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1858 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1859 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1860 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8612), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1861 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1862 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1863 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1864 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9124), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1865 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8393), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9124));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7993), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8393));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8243), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7993));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8508), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9068), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8612), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8243));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1870 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8052), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8137));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1871 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8695), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8543), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1872 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23415), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8052), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8695));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1873 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9095), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1874 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8477), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9095), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1875 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8589), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8477));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23415), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8589));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12710), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8775), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1879 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8775));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1881 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1882 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8081), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1883 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8081));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1884 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7926), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572));
NOR4BX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7926), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8720));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11994), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11022), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10527));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10499), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10638), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1892 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10665), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10791));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1893 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10952));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1894 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10800), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10471));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10539), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10800));
MX2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10411), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1899 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12038), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11994), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1900 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[36]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[35]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11974), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12710), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12038));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1901 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[36]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[18]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[36]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1902 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1903 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1904 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11775), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13321));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1908 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13016));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11814), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1910 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12224), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11853), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11775), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12399), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11814));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1912 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12880), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13147));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1913 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1914 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13298), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13117));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1915 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1916 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11745));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1917 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1918 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13216));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1919 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12015), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13298), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12684), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12547));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1920 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11667), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12224), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12880), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12015));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1921 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12181), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13284));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[4]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[3]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1927 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12984));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1928 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12567), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12200), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12181), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12780), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1929 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1930 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1931 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1932 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8402), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8901));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1933 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1934 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9135), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1935 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8660), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9135));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1936 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8402), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8660));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1937 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8208), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9079));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1938 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1939 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8515), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9013), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8293), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659));
OR4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8906), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9013), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8293), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7932), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8515), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8906));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8208), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7932));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1947 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11837));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1949 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11710));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1951 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1952 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11804));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1953 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12041), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13082));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1955 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13283), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13062), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12324), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12041));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1956 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12730), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12378), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12567), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11921), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13283));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1957 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12406), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12047), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12254), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13177), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12730));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1958 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12982), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12645), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11667), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12834), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12406));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1959 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8485), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1960 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8165));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8307), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1962 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8307), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8615));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1963 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1965 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8326), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8969), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1966 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8596), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8980), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8326), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1967 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8808), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8596));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1968 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8485), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23407));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1969 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12906), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1970 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12859), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12524), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11784), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12982), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12906));
OA21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1971 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[31]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[30]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1975 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1976 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1977 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13045));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8214), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I1979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8214), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8796), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1983 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8987), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1984 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1985 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1986 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8170), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8620), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8994));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1987 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7951), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7897), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8987), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8170));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1989 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1990 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1991 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8044), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1992 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8044));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1993 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1994 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1995 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8126), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8686), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8275));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1996 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8932), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8428), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8126));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1997 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7951), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8932));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1998 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I1999 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11902));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2000 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12920), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13181));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2002 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048), .A(N23926), .B(N23928), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12434), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13048));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2005 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[1]));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2006 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13013));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[0]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(N23926));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(N23928));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12775), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2013 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12084), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11707), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2014 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13079));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2015 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12392), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12775), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12470));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12909), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2017 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13095), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12737), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11874), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12909));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2018 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12349), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13213), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12920), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13095));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2019 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11791), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11853), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12349), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13313));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2020 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13113), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12959), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11791), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12047));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2021 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12072), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13113), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11911), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12645));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2022 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11943), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13067), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12072), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12524));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2023 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[35]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[34]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13331), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12859), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11943));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9102), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2025 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2027 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2028 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7996), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2029 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8268), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8433), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2030 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8114), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8268));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2031 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8679), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8534), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8114));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9102), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8372));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2033 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[35]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[17]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[35]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2038 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9133), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8292), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8555), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9051));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2044 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2045 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8639));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2046 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2047 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2048 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8401), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2049 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2050 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8658), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8401), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8232));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2051 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8148), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8555), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8658));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12711), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11772));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2055 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11807), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11677));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13145));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2058 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12873), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12540), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12711), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11807), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13335));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12583), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13249));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2061 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2062 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2063 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8342), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2065 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2066 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8300), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2067 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8300));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8135), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2069 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8196), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8135));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8564), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8891));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8196), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8564));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8963), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9141), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8155));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2074 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2075 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2076 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8236), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2077 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8236));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2078 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2079 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8030), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8764));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2080 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8842), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9017), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8030));
NOR4BBX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2081 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8665), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .BN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8842));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2082 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8963), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8665));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2083 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2084 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12843), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11972));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2085 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2086 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11963), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11865));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2087 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11962), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13253), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12583), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12843), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11963));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2088 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13054), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12200), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12873), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11962));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13100), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11741));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2091 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2092 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11834));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2093 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2094 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13114));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2095 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11774), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13061), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13100), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12358), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12074));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2096 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12216), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13317));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12572), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12812), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12744));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8435), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9093), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2101 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8865), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9093), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8865));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2105 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8261), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8474), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8525));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2107 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7902), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8220), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8474));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2108 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8175), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7902), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2109 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8175));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2110 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2111 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12034));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2112 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12714), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12357), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12216), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12572), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12503));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2113 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12683), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12323), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11774), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12714), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12737));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2114 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12139), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11765), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12902), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11986), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12683));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2115 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12532), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12165), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12378), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13054), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12139));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8124), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8538), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2118 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2120 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8815), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8858), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2121 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2122 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7950), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8611), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23399), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8815), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8986), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7950));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8124), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23399));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2128 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2130 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8514), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8400), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8835));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8952), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8656), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8086), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8952), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8656));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8951), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8784), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8514), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8086));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2135 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[16]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2136 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13125), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2137 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12193), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11821), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12756), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12532), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13125));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2138 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10971), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10736), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10879));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2139 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10971), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10687));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10608));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2142 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10475), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10475));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2144 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10616), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2146 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10854), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10754));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10849), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10498));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45208), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10648));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2149 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10595));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45200), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10572), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10509), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10421));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45208), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45200));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2152 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10849), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2153 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12798), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12798), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[29]));
XOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2158 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12188), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12949));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10818), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10957));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10652));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45206), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10777), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45190));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2165 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45530), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45206));
MX2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45526), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45530), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10552), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10682));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2168 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2169 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45195), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400));
MX2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11779), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11779), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2173 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13244), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12165), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13084), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2175 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12365), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13174));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2176 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12894), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12188), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13244), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12365));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2177 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11844), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13140), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12193), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11694), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12894));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2178 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12205), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12718), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13111));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2181 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12778), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12431), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12718));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2182 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[34]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[33]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11844), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12778), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13235));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2183 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[34]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[16]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[34]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2187 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8801), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8147), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2188 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8966));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8794), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2193 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7896), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8794), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8254));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2195 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8212), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8732), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7997));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2196 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8305), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8212));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2197 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8305));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2198 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9033), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8580), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7896), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8426));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2200 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9138), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9085), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9138));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8887), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8960), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8644), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2206 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2207 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2208 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8153), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8644), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7957), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2209 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8960), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8153));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2210 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8352), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7983));
NOR3BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2211 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9085), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8887), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8352));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12415), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11936));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2216 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12951), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13212));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2217 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2218 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11842), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11706));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2219 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11802));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2221 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11809), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11842), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12392), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12745));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2222 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12509), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12147), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13254), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12951), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11809));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2223 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11740), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13027), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12540), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12509));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2224 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12842), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12502), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11740), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12706), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11765));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2225 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2226 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13009));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2227 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12316), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12415), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12842), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11812));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23307), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11744));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2229 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23307));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2230 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12004), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13242));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2232 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2233 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12002));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2234 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13178));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2236 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8321), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8048), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8321));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8439), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8439));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9063), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8648), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8944));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8202), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9063));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8873), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7965), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8873));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8179), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2247 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8241), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8179), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8896), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7965), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8241));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2249 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8056), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2250 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8507), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8056));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2251 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8771), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8771));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2254 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8202), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7924));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2256 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12097));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2257 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12546), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12180), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12874), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11697), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12136));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2258 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13224), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12849), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12357), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12546), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13061));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2259 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12476), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12114), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13224), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12323), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13027));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2261 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8360), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2262 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8864), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8360), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8102), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8706));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2263 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2264 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8316), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8260));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8655), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8316), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2266 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8109));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8472), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8413), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8532));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8174), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8472));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8864), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8655), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8174));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2272 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11682), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2273 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11920), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12476), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11682), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12502));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2274 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13018), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12867), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12004), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11920));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2275 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11980), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13275), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12316), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11821), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13018));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2276 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[33]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[32]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12431), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13140));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2277 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[33]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[15]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[33]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2278 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13075));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12716), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12716), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[27]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2283 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23303));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12858));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8630), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8530));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8110), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2291 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2292 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8851), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2293 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8574), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2294 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7994), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8851), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8574));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2295 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8973), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7994));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8368), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8110), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9099));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8368));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11766), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12156));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2300 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13245));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2302 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2303 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11969));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2304 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12368), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11766), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12986), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13290));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2305 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11769));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12391), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11864));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2309 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141), .A(N23928), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2310 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12110), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13141));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2311 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13300), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13133), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12391), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12110));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2312 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12333), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12368), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13300), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13099));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11996), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11899));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12614), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13280));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2318 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12250), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11675));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2319 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12426), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12845), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2320 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2321 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12537), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12065));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2322 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12582), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12217), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12250), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12426), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12537));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2323 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13261), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12882), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12614), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12582));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2324 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12297), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11930), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12333), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13261), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12147));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2325 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10588), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10899), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10400));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2326 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10588), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10757));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10733), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10794), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10812));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10603), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11004), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10459), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10916), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10857), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10773));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2333 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10949), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10603), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10459));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2334 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[23]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10875), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10733), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760));
BUFX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[23]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11683), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23226));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2339 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13185), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12818), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12297), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12114));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2340 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12653), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12289), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12925), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13185));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2341 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8346), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8075), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8283), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8827));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8895), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9062), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8075));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8388), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8455), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8008), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8388), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8503));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2350 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8346), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8895), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8455), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2351 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12630), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2352 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8398), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2353 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8398));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8247), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8315), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8315));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8182), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9128));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2359 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8247), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7973));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8512));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2362 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12218));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2363 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2364 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12774), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11831));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2365 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2366 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12648), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13314));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2367 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12613), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12249), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13055), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12774), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12648));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2368 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2369 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11737));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2370 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12589), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11876));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2372 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12803), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11875), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12589));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2374 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12910), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12031));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2375 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12996), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11732), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13209));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2377 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2378 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12171), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12126));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2379 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13334), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12952), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12910), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11732), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12171));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2380 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13068), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12613), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12803), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13334));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2381 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13034), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12691), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13068), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12180), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12882));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2382 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12999), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12661), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12849), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11930));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2383 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2384 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12588), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12921));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2385 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12263), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12630), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12999), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12588));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2386 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2387 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13295), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13311));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2388 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11702), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12263), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13295), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13215));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2389 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12106), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12653), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11702));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2390 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[32]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[31]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12561), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12106), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13275));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8938), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2392 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8071), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8162), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8384), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8384));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2398 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9113), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8473), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2399 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8386), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8647));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2400 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7901), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7901));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2402 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9113), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8133), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8823));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8071), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8496), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8610));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2404 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[32]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[14]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[32]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2406 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2407 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8046));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8404), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8839), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8132), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8730));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8956), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8839));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2414 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8786), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8371), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8956), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8067));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8404), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8786));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[29]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8582), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8549));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2420 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2421 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8913));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2422 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8582), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8687));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8378), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8128), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8276), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8215), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8640), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8378));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313), .A(1'B0), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[28]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2428 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2429 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[28]));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8565), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8031), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7920), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2434 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8409), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8031), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7911), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7920), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8892), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8841));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[27]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8565), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8714), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8409), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8892));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2437 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544), .A(1'B1), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[27]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2438 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8437), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8662));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8222), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2441 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2442 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8050), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8501), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8176), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8222), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8050), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2445 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8437), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8176));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2446 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248), .A(1'B1), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[26]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2450 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8588), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8227), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8588));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7966), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8459), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8348), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7966));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9065), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8096));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2457 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8650), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8626));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2458 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7925), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9065), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8242), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8650));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2459 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8113), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8079), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8459), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7925), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8897));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2461 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964), .A(1'B1), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[25]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2462 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412), .B(N23926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[42]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12810));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8975), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8308));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8369), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8975), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2469 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8632), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8886), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8369), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2470 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2471 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2472 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8531), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8924), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8531));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8772), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[24]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8632), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8747), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8267));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2476 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[24]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9007), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8958), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8018), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2481 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2482 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8121), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2483 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8755), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8121));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2484 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8880), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8755));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2485 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8834), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8880), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2486 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8854), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2487 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8064), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8489));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8553), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8183), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8704), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9131), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8834), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8553));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[23]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8018), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9131));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[41]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[42]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2493 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[23]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[41]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[41]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2495 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2498 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2499 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15513), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2500 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12918), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11700));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2503 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13139));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2504 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12965), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12626), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12918), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12749), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12818));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2505 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2506 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12826), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[23]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[24]));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12826));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12046), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12769));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12397), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13206));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2514 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12791), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12447), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12661), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12046), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12397));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9097), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7886));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9097));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8675), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9071), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8204));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2519 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9025), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2520 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8627), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9025), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2521 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8922), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8725));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7941), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8971));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8319), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7941), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8761), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8723));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23391), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8675), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8627), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8319));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23391));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11898), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2529 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12155), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11782), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12919), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12217), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12005));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13170), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11799));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12284), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11704));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12646), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11915));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2535 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12837), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13170), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12284), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12646));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11933));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12573), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12094));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11897));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2542 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2543 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8423), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2544 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8517), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8272), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8423), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8464));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2547 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8272), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8251), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8856), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8251), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7933));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7892), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8355), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2554 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8811), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8856), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7892));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2555 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8908));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2557 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8682));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2558 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9106), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8811), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8983));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8120), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9106));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12280));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2562 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12647), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12285), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12573), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12427), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12704));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2563 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12400), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12033), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12647));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2564 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11800), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12185));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13020), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13278));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13328), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11999));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2570 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11696), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12985), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11800), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13020), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13328));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2571 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13107), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11696), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12952));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2572 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12857), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12516), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12400), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13107), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12722));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2573 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12123), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12155), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12857));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2574 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12979));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2576 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12088), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11711), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11898), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12123), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12220));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2577 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12053), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11676), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12791), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12088), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11893));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2578 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12438), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12081), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12965), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12053));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2579 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[31]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12438), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12677), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11728));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8160), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2581 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8524), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7976), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7971), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8160), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8939));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9080), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8505));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2585 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8524), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8568), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9023));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8361), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8357), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8946));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7883), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2588 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9090), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2589 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7883), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9090));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8361), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8103));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2591 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[31]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[13]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[31]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2592 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10986), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10490));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2594 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2595 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11024), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45780), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10760));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2596 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10841));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2597 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2598 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10611));
MX2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10954), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10464), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2600 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13252), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13252), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9126), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2603 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2604 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8395), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2605 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8065), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8613));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2606 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8802), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8065));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7970));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8779), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9009));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23383), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9126), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8779));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2610 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2611 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2612 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8702), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2613 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8244), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8702));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2614 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23383), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8244));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12821), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2616 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12823), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12481), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12691), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12821));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12579), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11763));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13093), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12245));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2621 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9015), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8643));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8191), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8491));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2623 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8445), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8336));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2624 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8295), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8191), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8445));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2625 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8884), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8233), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2628 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8916), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8884), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7915));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2629 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8295), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8916));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2630 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9015), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8560));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12340));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12804), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11862));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2635 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11957), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13247), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13093), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12350), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12804));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12352), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12655));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2638 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11916), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11767));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2640 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12870), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12352), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11916));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2642 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12207), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12153));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2643 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2644 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12063));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2645 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2646 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12069), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11967));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2647 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12679), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12207), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12942), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12069));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2648 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12433), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12870), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12679));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2649 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12189), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11815), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12433), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12249), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12040));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2650 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11938), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13231), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12189), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11782), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12516));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11846), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13041));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2653 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11901), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13192), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11747), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11846));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2654 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11863), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12823), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12579), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11901));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2655 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2656 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13274));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12824));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11827));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2661 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12632), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12269), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11668), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12037), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12213));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2662 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12601), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12632), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11711), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12447));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2663 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12761), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12411), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12626), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11863), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12601));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2664 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[30]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12761), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12991), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12081));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2665 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8480), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8696), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8480), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9043));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9045));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8674), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2671 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9098), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8999), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8674), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9098));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2674 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8282), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8009), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8999));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2675 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8696), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8282));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2676 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[30]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[12]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[30]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2679 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13142), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12779), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12497), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12285), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12985));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12738), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12310));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2683 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13208), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11828));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2684 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11836), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12215));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2686 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12707), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12351), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12738), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13208), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11836));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2687 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12472), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12109), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12534), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12707), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13247));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8914), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8964));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8199), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2690 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8469), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8199));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8862), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8469));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8666), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7919));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2694 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8666), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7986));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8099), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8899));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8845), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8735), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9037));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8862), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8845));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2699 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2700 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8312), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7923), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2701 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8420), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8312), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2702 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8429), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8420));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2703 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8172), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8429));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11987), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12401));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12463), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11929));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12606), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12124));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2710 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11990), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11987), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12463), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12606));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11672));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11926), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2714 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11734));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13285), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12292));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12904));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2717 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12202), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12319), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13285), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2718 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11731), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12680), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12202));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2719 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12221), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11848), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12472), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11731), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12073));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2720 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12889), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12750), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13142), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12221));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2721 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8726), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8576), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8912), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8726));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8271), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7890), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8793), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8340), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8576));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8847));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8544), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8907));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8535), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8422));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8855), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7998), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8855));
NOR3BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2729 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8271), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8535), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7998));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12121), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2732 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13108));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2733 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12666), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12889), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12121), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13138));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12958), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12885));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23421), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23282));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2738 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[22]));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12784), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12690));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2744 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13333), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11669));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2745 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11717), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13003), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12958), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12784), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13333));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2746 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11685), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12970), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12666), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12481), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11717));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10780), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10921));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10402));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10680), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10820), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10426), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10577));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10820), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10813));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13149), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13149));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2755 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8334), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2757 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8931), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7913));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8838), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8334), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8022));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7952), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9084));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8838), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8622), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8707), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8497));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13031), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12058));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2762 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11976), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11815), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13031));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11891));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2765 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12456), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12095), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11976), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11841), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13231));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2766 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12417), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12061), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12456), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13192), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12269));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2767 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13323), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12938), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13157), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11685), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12417));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2768 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[29]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13323), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11676), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12411));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2769 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8394), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8302));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2770 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8144), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2771 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8614), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8144));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2772 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8900), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8829));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2773 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8082), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8552));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8778), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8245), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8692), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2777 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7927), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8778), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8245));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2778 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8614), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8900), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8082), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7927));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2779 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[29]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[29]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2780 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2781 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2782 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12619), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12947));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2783 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12743));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2786 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12948), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11730));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2787 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11753), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13039), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12619), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12440), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12948));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2789 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12384), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12372));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2790 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2791 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12276));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12836), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11895));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2794 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12940), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12603), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12384), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13127), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12836));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2795 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2796 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12028));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11954), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11795));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8766), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2800 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8280), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2801 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9060), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8280), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2802 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8197), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7921), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9060));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2803 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8766), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8197));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2804 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8715), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2805 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9117), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2806 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2807 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9117), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2810 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8136), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2811 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8452), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8344));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8715), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8452));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8033), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9019));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12465));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2816 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13158), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12793), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11954), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12757), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13281));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2817 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11768), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13058), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11689), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13158));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2818 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13180), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12811), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11768), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12318), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13022));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2819 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12927), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12592), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13180), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12779), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11848));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12777), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13171));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2822 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12696), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12339), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12554), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12777));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2823 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13162), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12796), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11753), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12696), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12306));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13132), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11960));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2827 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8680), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8733), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8826), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8468), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9087), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8572), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8548), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8619), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9035));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8045), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9087), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8619));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7985), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7985), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8219), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8668));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2834 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8376), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8213));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8733), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8045), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8376));
OAI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12329), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2838 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12240), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12182));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12091));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2841 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2842 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11995));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2843 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12027), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13326), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12978), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12101));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2844 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12505), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13286), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12027), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11829));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2845 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2846 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12430));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2847 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2848 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11964));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2849 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2850 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12640), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12151));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2851 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12271), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12023), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12498), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12640));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11830), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13218));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12412));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12026), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12528));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2855 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13195), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12825), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11830), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13121), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12903));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12765), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12338));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2858 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2859 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13248), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11858));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2860 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2861 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11867), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12242));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2862 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12973), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12633), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12765), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13248), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11867));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2863 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12740), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12271), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13195), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12973));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2864 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13217), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12844), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12740), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12351), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13058));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2865 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12256), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11888), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12505), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13217));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45518), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45533), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10407));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12152), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[25]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45525), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[26]));
BUFX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12152));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2870 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12432), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13239));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2871 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12010), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12256), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12432));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2872 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12490), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12129), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13132), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13267), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12010));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2873 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12239), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11869), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12490), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13003), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12095));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2874 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13126), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12768), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12970), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13162), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12239));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2875 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[28]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[27]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13126), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12232), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12938));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8373), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8421), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9048), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8028), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2879 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8061), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8373), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9048), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2881 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8752), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9105));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2882 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8328), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8752), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8928), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2883 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8061), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8328));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2884 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[10]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[28]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13007));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12610), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11793));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2892 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11786), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13078), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12592), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12255), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12610));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2893 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2894 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12795));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[21]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156));
CLKXOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2899 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2900 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11892), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12600));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2901 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10631), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10514), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10654));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2902 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10631), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10546));
NAND2BX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2903 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[18]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2904 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11803), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13097), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12793), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12603), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13326));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12025));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2908 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12122));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12056), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2910 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12939), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12560));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2912 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13043), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12056), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13155), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12939));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2913 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12098), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13011), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13043));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2914 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2915 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13163), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12307));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2916 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12507), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2917 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12871), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11925));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2918 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2919 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12277), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12212));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2920 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13006), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12667), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13163), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12871), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12277));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2921 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12770), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12420), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12098), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13006), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11903));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12448));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13225), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11998), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12495));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12762), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12846));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12398));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2927 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12308), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11940), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13324), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12762), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12418));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2928 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2929 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11723), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12060));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2930 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12064), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12308), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11723), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12825));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2931 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12541), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12174), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12064), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12386));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2932 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12291), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12141), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11803), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12541));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2933 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12961), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12622), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12811), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12291));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2934 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12727), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12375), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12079), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11892), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12961));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2935 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13199), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12830), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11786), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12727), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12339));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2936 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2937 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12771), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12022));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2938 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8070));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2939 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7960), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8788), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8436), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9012), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8436), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8693));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8499), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8684));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9115), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7960), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8763), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8499));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[6]));
OAI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13260), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2947 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13308));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2949 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12049), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11670), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13260), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11888), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12071));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2951 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11701), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12855));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2952 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2953 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13187), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12660));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2955 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11883), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13072));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2956 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12758), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12407), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11701), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13187), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11883));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2957 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12527), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12161), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12771), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12049), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12758));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2958 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12279), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12527), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13039), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12129));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2959 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12945), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12605), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13199), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12279));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2960 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[27]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[26]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12945), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12061), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12768));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8294), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2962 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8955), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2963 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7980), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8955), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7910));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7914), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2965 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8201), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2966 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8403), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8335), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8997), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2967 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8250), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8721), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7914), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8708), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8403));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2968 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8294), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8606), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7980), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8250));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2969 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[27]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[9]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[27]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2970 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2971 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13237), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12861), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12375), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13306), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13078));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12424), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12086));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2975 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12248), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11855));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2976 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45786), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2977 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10863), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11009));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10755), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10725), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45786), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10599), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45792), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10843));
MX2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10897), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10460));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2983 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2984 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2985 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12272));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2986 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2987 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12797), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12370));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2989 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11760), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12089));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2990 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12832), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12797), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11760));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2991 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2992 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12462));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2993 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2994 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11991));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2995 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I2996 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12179));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2997 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12131), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12062), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12533), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12673));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2998 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12799), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12458), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12131), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11940));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I2999 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11839), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13129), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12799), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12633), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11686));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3000 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13258), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12876), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13097), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11839));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3002 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[18]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12659), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12506));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3005 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12995), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12654), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13258), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12844), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12659));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3006 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11824), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12424), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12248), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12995));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8968), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8458), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8533));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8526), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8090), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004));
NOR3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8800), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8859), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9064), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8526));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8848), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8262), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8848), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8917), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8741));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8414), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8598), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3013 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8719), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3014 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8414), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8719));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3015 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8968), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8800), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8262), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8669));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[5]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3017 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12543), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3018 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3019 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11695));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3020 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12083), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11924), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12543), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11692));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3021 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3022 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12713));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3023 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12993), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12915));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3025 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13176), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13136));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3027 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12786), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12993), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13176));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3028 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12563), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12194), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12083), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12786));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3029 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12312), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45350), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11824), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12563), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12161));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3030 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12977), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12639), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12830), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13237), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12312));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3031 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[26]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11869), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12977), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12605));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8012), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8837));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3033 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8127), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8911), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8012));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8621), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8098), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8860), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7978), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8098));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3038 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8171), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8539), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8734), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8621), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8860), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8171));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9110), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8383), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8539));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8127), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9110));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3044 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[8]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[26]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3045 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3046 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3047 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3048 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9116), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8949));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3049 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8569), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8498));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3050 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8604), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8116), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3051 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8237), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8039));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7988), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8745), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8005));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3055 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8237), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8893));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8451));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8343), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8604), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8324));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3058 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11872), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11923));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3061 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12068), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12144));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3062 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12265), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3063 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12703), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12347), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13193), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12265));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12966), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12142));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3065 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3066 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12525));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3067 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12864), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12529), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12966), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11684));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3069 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13200), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12336));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12453), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12428));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12238));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3074 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11948), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13241), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13200), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12453), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12313));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3075 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11909), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13202), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12698), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12864), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11948));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3076 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11870), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13165), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11720), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12667), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11909));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3077 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3078 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12575), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12211), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11870), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13033), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12420));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3079 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12342), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3080 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12296), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12569));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3081 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12326), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11966), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12174), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12575), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12296));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3082 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11856), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11872), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12068), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12326));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3083 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13276), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12897), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12407), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11670), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11856));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3084 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9122), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8460), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3085 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8872), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8776), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3086 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8594), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8185), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8609), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8631));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3087 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8805), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8974), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7958));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3088 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8390), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8700), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7906), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23375), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8872), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8594), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8390));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3091 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9122), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23375));
OAI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3092 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11806), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3093 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3094 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11761));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3095 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13029), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11806), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12983));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3096 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12652), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12976));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12475), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12767));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3101 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13203));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3102 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12118), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11742), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12652), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12475), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12809));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3103 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12596), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12654), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13029), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12118));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3104 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45345), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45394), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12596), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13115), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12194));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3105 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13012), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45377), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12861), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13276), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45345));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3106 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[25]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[24]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13012), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11907), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12639));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3107 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[25]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[25]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3108 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3109 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3110 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13166), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11989));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3111 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12332), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3112 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12167), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12057));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13050), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12148));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12482));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12971), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12484), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12883), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12590));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3118 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12096), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12492));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3120 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11762), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13052), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12347), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12971), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12096));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3121 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12675), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12314), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12167), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13050), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11762));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3122 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12642), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12281), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12675), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11756), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12493));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3123 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12607), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12243), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12458), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12332), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12642));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3124 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13293), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12913), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13129), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12607), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12211));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12206));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3127 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12819), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12479), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13166), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13293), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11687));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3128 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13315), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11705), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12441));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3130 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12395));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12702), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12209));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12305));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3135 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12501), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12135), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12829), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12702), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11944));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3136 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11725), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13015), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12529), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12501), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13241));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3137 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13263), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3138 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11691), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13202), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11725), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13263));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3139 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13329), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12946), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11691), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13165), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12243));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12822));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3142 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12469), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13272));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3144 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13064), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13329), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12116), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12469));
BUFX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13137));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3146 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11979), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11932), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12627));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8397), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8416));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3149 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7930), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8397), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8055));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8903), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9130), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8995), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8016));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3152 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8948), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8962), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9086), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8953), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3153 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9073), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8948));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9044));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8274), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9004), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8461), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7974));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7930), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8903), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9073), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8461));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3158 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[3]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12742), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12644), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11823));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3162 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12361), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12000), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11932), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12742), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12644));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3163 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11896), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13189), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13064), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11966), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12361));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3164 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45389), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45721), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13150), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12226));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3165 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45371), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12897), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13315), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45389));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3166 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[24]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45342), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45371), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45350), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45377));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9024), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9069), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3168 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7938), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8095), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8279), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9024), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8117));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3169 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9041), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8998), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7938));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8427), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8304));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8221), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8527), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8364), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8188));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3173 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8587), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8035), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8364));
NOR4BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8318), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8221), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8051), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3175 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9041), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8318));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3176 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[24]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[6]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[24]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3177 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3178 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12461), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12117));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3183 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13339));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12637), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12330));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3187 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12183), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11810), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12461), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12105), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12637));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3188 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11934), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13227), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12183), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12000), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12717));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12099), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12173));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11729), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11727));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3193 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11718), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12556));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3195 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3196 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3197 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12491), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12459));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3198 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12321), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11959), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11718), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13190), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12491));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3200 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11794), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12119));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13086), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12176));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13238), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12366));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3206 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12344), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12270));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3207 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13025), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13086), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13238), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12344));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3208 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13210), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12321), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11794), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13025));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3209 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12545), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11910), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3210 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12467), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12103), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12314), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13210), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12545));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3211 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12429), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12281), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12981));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3212 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12922), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12099), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11729), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12070));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8374), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8785));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8813), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8154), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8167), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8001), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3216 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8636), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8167), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7999), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8683), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3217 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8488), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8813), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8636));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3218 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8488));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3219 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8982), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7948), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8374), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9032));
OAI22X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12029), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3221 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13273), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13223), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12686));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3224 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12282), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11887));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3225 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12394), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13223), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12282));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3226 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12881));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3229 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11922), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13104));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3230 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13102), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12747), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12429), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11739), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11922));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3231 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11973), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13264), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12922), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12035), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12747));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3232 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3233 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12792));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3234 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3236 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11752), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12586));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11743), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3238 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12489));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3240 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12969), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12629), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11752), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11743), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12526));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11983), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12334));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12478), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12708));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12517));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13004), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12457), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12519), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12615));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3246 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11927), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12478), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13230), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13004));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3247 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11708), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12997), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12969), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11983), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13220));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3249 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12732), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12234));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3250 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3251 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12522));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12862), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12425));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3254 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12656), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12295), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12732), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12130), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12862));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3255 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12112), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11735), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12656), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11927), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11959));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3256 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12814), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12474), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12682), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11735));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3257 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12989), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12649), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11808), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12840), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12814));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3258 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8540), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7940), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8006));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8550), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8762));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8645), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3261 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8820), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8125), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8659));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3262 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8736), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8608), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3263 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8380), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8736), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8930));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3264 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8094), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8216), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8380));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8933), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8820), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8094));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3266 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9036), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8187));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8003), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9036), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8685));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23367), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8933), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8003));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8540), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23367));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8446));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3272 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8023), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8481));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3274 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8516), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9014), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8023));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3275 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8790), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8583), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3276 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8709), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8646));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3277 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8049), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8520));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3278 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9081), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8269), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8457), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7981));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8089), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8709), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9081));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8516), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8790), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8089));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[1]));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3282 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12237), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3283 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12251), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11880), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12989), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12237));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12274), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12390));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13005));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3289 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13234));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3291 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13205), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12017));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3292 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12955), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12617), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12841), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13205));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3293 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12007), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13302), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12251), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12274), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12955));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3294 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12287), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11918), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12135), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13052), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12112));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3295 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13173), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12805), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13015), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12103));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3297 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13026), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12944));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13214), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13167));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3300 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12219), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11843), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13173), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13026), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13214));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3301 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12941), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12414), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3302 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12893), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3303 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12848), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12739));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3304 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3305 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11912), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11956));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3306 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13135), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12941), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12848), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11912));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3307 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12884), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12946), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12219), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13135));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3308 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12693), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12335), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11810), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12549));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3309 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45718), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13227), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11973), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12693));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3310 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12853), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12913), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12394), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13102));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3311 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45711), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12853), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13189));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3312 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3313 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12975), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12267));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12288), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13037));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3317 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12054));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3318 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12150), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11778), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12975), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12288), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12802));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3319 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12628), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12264), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12150), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12687), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11742));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3320 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45692), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12884), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11778), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12512));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3321 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45708), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45695), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12264), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11934), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45692));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3322 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45677), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45718), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45698), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45695));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3323 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8879), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8812), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7959));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3324 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9008), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8879));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3325 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8331), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8832));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3326 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8442), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8362), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8209));
NAND4BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8290), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8331), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8178), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8442), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8066));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8063), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7898), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7945), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8184), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8194), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8063));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8978), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7908), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9119), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8184));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3331 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8017), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8290), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8978), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9056));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3332 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45353), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45687), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12933), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12628), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45711));
ADDFHXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3333 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45380), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45721), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45687));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3334 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45677), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45700), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45713));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3335 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7929), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8876));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8418), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7929), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8934));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3337 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8976), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8418));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8545), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8077));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3339 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9074), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9092));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8163), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8463), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8777), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9074));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3341 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8266), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8163));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8852), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8365), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7893));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8634), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9027), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8603), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8852));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45391), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8976), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8266), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8263), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8634));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3345 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45400), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45353), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45394), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45358));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3346 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45380), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45391), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45386));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8150), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3349 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8663), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8150));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3350 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8091), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9052), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9034), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8663));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3351 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9030), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8750), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8870));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3352 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8799));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3353 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7947), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8297));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3354 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8616), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8789));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3355 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8616), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8270), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9139));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3356 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8038), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8770), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8727));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3357 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8091), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9030), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8038));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3358 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3359 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13017), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11790));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3360 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3361 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12233));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3362 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12044), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13337), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12805), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13017), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11722));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3363 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12723), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12371), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12776), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12044), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11843));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3364 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13159), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23315), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3365 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3366 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12146), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12852));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3367 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12075), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13159), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11918), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12146));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3368 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3369 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11904), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12452));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3370 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3371 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12380), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12303));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3372 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3373 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13277), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12393));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3374 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12688), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11992));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3375 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12555));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3376 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13040), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12980), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13042), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12643));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3377 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12389), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12030), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12688), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13268), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13040));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3378 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12059), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11681), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12380), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13277), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12389));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3379 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12444), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12087), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12059), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12295), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12997));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3380 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12746), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23286), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12192));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3381 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11890), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13183), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12444), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12746), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12474));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3382 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3383 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12833), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12082));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3384 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12783), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12437), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12649), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11890), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12833));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3385 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12752), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12404), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12075), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11904), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12783));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3386 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11783), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12585), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12752), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13302));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3387 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45668), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13036), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13264), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12723), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11783));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3388 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45684), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45668), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45679), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45705));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3389 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45720), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45684), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45724));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3390 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3391 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3392 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8874), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8320), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8713));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3393 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45383), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8874), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8758));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3394 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45368), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8084));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3395 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8180), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8943));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3396 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45341), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8180), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8824));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3397 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8890), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3398 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8653), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8043));
OR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3399 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9121), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8593), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8699), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8322));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3400 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9121), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3401 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45397), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45383), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45368), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45341), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45355));
ADDFHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3402 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45400), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45397), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45342));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3403 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3404 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3405 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3406 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942));
NOR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3407 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8296), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8021));
NOR4X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3408 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8843), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8441), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8523), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8717));
AND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3409 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8453), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9077), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8825), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8434), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8181));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3410 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8453));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3411 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8410), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8303), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9104));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3412 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8563), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8888));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3413 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8157), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8843), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8410), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8566));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3414 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3415 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12504), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13303));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3416 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3417 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12325), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13070));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3418 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3419 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12676), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11852));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3420 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11851), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13143), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12504), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12325), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12676));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3421 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11818), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13109), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11880), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11851), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12617));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3422 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3423 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12137), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11693));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3424 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3425 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11961), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13134));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3426 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3427 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12317), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11919));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3428 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11673), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12964), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12137), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11961), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12317));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3429 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13310), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12930), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11699), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12437));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3430 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3431 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12359));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3432 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23308));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3433 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12828), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12580));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3434 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12409), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12051), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12669), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13183), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12828));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3435 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3436 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12896), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12455));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3437 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3438 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12162), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12553));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3439 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3440 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12016), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12362));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3441 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13098), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12896), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12162), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12016));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3442 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12764), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12416), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12629), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13098), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11681));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3443 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3444 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3445 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13154), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12764), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12032), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12087));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3446 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3447 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12133), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12201));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3448 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3449 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13201));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3450 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12935), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12599), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12789), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12133), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13255));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3451 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12943), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3452 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3453 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11787), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12612));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3454 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11965), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13287));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3455 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3456 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12564), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12518));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3457 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13229), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11787), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11965), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12564));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3458 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12178), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11805), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12030), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13229), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12741));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3459 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11833), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13124), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12943), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12178), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12416));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3460 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3461 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13063), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12972));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3462 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12229), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11859), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12695), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11833), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13063));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3463 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3464 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11951), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11985));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3465 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3466 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11764), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11758));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3467 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3468 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12311), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12419));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3469 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12021), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11951), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11764), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12311));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3470 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13119), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12759), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12935), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12229), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12021));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3471 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12377), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13143), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12409), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13119));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3472 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13270), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12891), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13109), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13310), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12377));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3473 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3474 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12515));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3475 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3476 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13008), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12299));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3477 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11819), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13112), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3478 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11773), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12912));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3479 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3480 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12140));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3481 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12625), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12259), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13154), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11773), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12496));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3482 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12593), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12223), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13198), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13008), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12625));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3483 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12557), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12190), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12593), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13337), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12404));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3484 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12520), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12157), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12371), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11818), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12557));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3485 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[18]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13270), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13071), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12157));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3486 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[18]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3487 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[19]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12520), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12335), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13036));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3488 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[18]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3489 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3490 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13035));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3491 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12241), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12755));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3492 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12877), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3493 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12591));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3494 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11946), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12671));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3495 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12423), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12067), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12877), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13307), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13077));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3496 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12905), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3497 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13316), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12421));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3498 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12304), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11937), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12423), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13316), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12854));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3499 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12879), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12544), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12241), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12304), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11805));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3500 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12571), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12204), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12712), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12879), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13124));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3501 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23313));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3502 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12487), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11679), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12968), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12638));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3503 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12734), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12381), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12571), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12487), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11859));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3504 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12196), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11826), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12964), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12259), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12734));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3505 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13080), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12729), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12930), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12223), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12196));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3506 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[17]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13080), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12190), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12891));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3507 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[17]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3508 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3509 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8927), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9140), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9134), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9125));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3510 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8379), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8130), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8991));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3511 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7899), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8724), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9022));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3512 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7899), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8159));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3513 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8935), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N9020), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8097), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8628));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3514 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8313), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7887), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8207));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3515 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7953), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8935), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8313));
NAND3BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3516 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8277), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8309), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8456), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8002));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3517 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8672), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7882));
NAND3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3518 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8819), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8363), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8689));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3519 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8277), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8819));
NAND4XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3520 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8379), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8492), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7953), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N8234));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3521 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[19]), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[19]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3522 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3523 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3524 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3525 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3526 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15524), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3527 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444), .A(N22905), .B(N23646));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3528 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15035), .A(N23051), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3529 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3530 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13047), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12327));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3531 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3532 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12356), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13101));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3533 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3534 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13336));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3535 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12689), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12328), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13047), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12356), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12538));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3536 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3537 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12868), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12113));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3538 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3539 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11884));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3540 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12235));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3541 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13233), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12548));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3542 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11746), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13032), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12868), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12705), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13233));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3543 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13060), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12709), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12204), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12689), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11746));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3544 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12536), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12169), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13060), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13319), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12381));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3545 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3546 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12934), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12485));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3547 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3548 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12195), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12584));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3549 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3550 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12641));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3551 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12175), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12570));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3552 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3553 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12595), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12550));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3554 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13038), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12175), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12595));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3555 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13131), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12773), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12934), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12195), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13038));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3556 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13161), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12405));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3557 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13002), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12664), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11937), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13131), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13161));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3558 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11968), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13259), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11785), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13002), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12544));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3559 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3560 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13243), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12052));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3561 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12450));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3562 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11942), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12542), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12177), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12483));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3563 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12355), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11993), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11968), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13243), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11942));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3564 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3565 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12875), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13269));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3566 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23302));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3567 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11757), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12266));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3568 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3569 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13056), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11820));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3570 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13289), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12907), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12875), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11757), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13056));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3571 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11796), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13092), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12355), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13289), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12599));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3572 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12900), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12566), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12051), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12759));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3573 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[15]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12536), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11826), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12566));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3574 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[16]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12011), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12900), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12729));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3575 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[16]));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3576 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15141), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[15]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[15]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3577 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12454), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3578 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12214), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11840), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12773), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12067), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12454));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3579 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12045), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3580 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11997), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13164));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3581 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12093), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11716), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12664), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12214), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11997));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3582 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13096), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12203));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3583 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23344));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3584 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13116), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12435), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12499), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12697));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3585 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12039), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13332), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13096), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11671), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13116));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3586 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3587 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12227), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12608));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3588 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3589 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11857), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12668));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3590 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12387), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11832));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3591 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12787));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3592 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13148), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N10622), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13089), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12724));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3593 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13327), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13123));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3594 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12860), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13148), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13327), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__61[2]));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3595 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12460), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12100), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11857), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12387), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12860));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3596 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12748), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12396), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13332), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12227), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12460));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3597 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12128), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12039), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12748));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3598 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12917), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12578), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12562), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12128), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11840));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3599 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3600 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12700), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12388));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3601 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3602 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12172), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11724));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3603 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12794), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12917), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12700), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12172));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3604 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12480), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13259), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12093), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12794));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3605 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12143), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11771), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11993), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12907), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12480));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3606 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[14]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12143), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12169));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3607 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[14]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3608 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3609 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12170));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3610 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3611 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12348), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11952));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3612 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11866), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13160), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12531), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12348), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11716));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3613 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13191), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12820), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13032), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12328), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11866));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3614 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[13]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13191), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12709), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11771));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3615 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[13]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3616 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15456), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15155));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3617 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3618 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12164), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12231));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3619 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3620 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11988), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12014));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3621 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12720), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12364), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12164), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11988), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12578));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3622 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23304));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3623 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12092), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11715), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12449));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3624 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3625 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13291), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13232));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3626 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3627 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11788));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3628 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12003), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13296), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12343), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13291), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11801));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3629 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12604), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12236), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12720), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12003), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12451));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3630 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[12]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12604), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12120), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12820));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3631 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[12]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3632 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3633 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13094), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11847));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3634 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12665), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3635 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11811), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13106), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12396), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12665), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13312));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3636 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3637 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13282), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12080));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3638 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11906), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13197), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13094), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11811), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13282));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3639 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11719), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13340));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3640 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12956), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3641 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12908), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13301));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3642 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12827), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12488), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11749), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11719), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12908));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3643 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11781), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13066), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11906), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12827), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13296));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3644 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[11]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13160), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12236));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3645 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[11]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3646 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3647 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11792), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12294));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3648 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3649 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12736), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11914));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3650 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3651 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12574), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11690));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3652 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3653 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12901), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12138));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3654 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12552), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12187), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12736), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12574), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12901));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3655 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12636), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12273), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12488), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11792), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12552));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3656 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[10]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12364), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13066));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3657 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14950), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[10]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3658 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12974));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3659 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13083), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12914), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12577), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12354));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3660 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11939), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12618));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3661 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3662 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12208), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11755));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3663 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13169), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11939), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12100), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12208));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3664 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13266), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12886), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13106), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13083), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13169));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3665 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[9]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13197), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13266), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12273));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3666 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[9]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3667 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12036));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3668 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12568), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12199));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3669 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23285));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3670 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12856), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12253));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3671 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11941), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13236), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12856), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12523), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12410));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3672 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3673 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12385), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11981));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3674 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12247), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11871), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12568), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11941), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12385));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3675 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[8]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12187), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12247), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12886));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3676 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15038), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[8]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3677 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3678 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12024), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12048));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3679 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3680 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11835), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11817));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3681 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12184));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3682 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12486), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12125), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12262));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3683 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12670), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12024), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11835), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12198));
ADDFXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3684 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[7]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12670), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12801), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11871));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3685 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15403), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[7]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3686 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12154), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11881));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3687 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12602), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12443), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12763));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3688 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3689 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11879));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3690 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13074), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12154), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12602), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13128));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3691 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12521));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3692 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12108));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3693 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13069), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13175));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3694 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13305), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12924), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13156), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13069));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3695 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3696 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12766), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11950));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3697 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12367), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12807));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3698 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13299), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23290), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3699 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11845), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13299));
ADDHX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3700 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12587), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12367), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N11845));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3701 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12374), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12924), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12766), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12587));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3702 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12160), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13322), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13305), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12374));
ADDFX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3703 (.CO(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[6]), .S(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13074), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13236), .CI(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12160));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3704 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[6]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3705 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15492), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[5]));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3706 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15201), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[4]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3707 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12309));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3708 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12609), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12244), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12166));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3709 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15580), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[3]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3710 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12468), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3711 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12013));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3712 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[2]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3713 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12104), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23296));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3714 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N13073), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12725), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N12077));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3715 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15519), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[1]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3716 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15144), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[2]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3717 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15129), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15519), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15144));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3718 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15270), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[1]), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[1]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15284));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3719 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14960), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15129), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15270));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3720 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15429), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[3]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3721 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15453), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15580), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14960), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15429));
OAI22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3722 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15199), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15201), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15453), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[4]), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[4]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3723 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15345), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[5]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3724 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14974), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[6]));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3725 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14994), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15345), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14974));
AOI31X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3726 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15068), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15120), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15492), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15199), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14994));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3727 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15257), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[7]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3728 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15023), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15403), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15068), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15257));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3729 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[8]));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3730 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14970), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15038), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15023), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15556));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3731 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15177), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[9]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3732 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15498), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15322), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14970), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15177));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3733 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15466), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[10]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3734 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15097), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[11]));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3735 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15327), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15466), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15097));
AOI31X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3736 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15485), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15234), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14950), .A2(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15498), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15327));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3737 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15379), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[12]));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3738 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15560), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15531), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15485), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15379));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3739 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15011), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[13]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3740 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15298), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[14]));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3741 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15311), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15011), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15440), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15298));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3742 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15084), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15456), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15560), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15311));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3743 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15590), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[15]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3744 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15210), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[16]));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3745 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15000), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15355), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15590), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15210));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3746 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15141), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15084), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15000));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3747 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3748 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3749 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3750 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15297), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15378));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3751 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15412), .A(N22772));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3752 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[17]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3753 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15033), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[18]));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3754 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3755 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15171), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15316));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3756 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15461), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14945));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3757 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3758 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3759 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15089), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15230));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3760 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15373), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15522));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3761 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3762 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15006), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15148));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3763 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15288), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15433));
AOI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3764 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3765 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3766 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15376), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3767 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15584), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15062));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3768 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15205), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15349));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3769 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3770 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15495), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14979));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3771 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15124), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15262));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3772 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3773 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3774 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15407), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15561));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3775 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15041), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15182));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3776 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3777 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15326), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15470));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3778 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14954), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15101));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3779 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3780 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3781 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15044), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3782 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303), .A0(N23646), .A1(N22903), .B0(N22875));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3783 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15384), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15238));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3784 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15535), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15016));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3785 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3786 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15159), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15302));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3787 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15445));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3788 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3789 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3790 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15216), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15076));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3791 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15509), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15359));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3792 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3793 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15133), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14989));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3794 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15417), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15274));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3795 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3796 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3797 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3798 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15051), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15572));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3799 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15335), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15191));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3800 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3801 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15482), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14964));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3802 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15111), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15248));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3803 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3804 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3805 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15313));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3806 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15544), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15394));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3807 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15167), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15027));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3808 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990));
OAI2BB2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3809 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15424), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15455), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15309), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3810 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15032), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15575), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15424));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3811 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15283), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15172), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15361), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15032));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3812 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15553), .A0(N23051), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303), .B0(N23049));
OAI21X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3813 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[49]), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15035), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15412), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15553));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3814 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[49]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3815 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45117), .A(N21282), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3816 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3817 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3818 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3819 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3820 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3821 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3822 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3823 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3824 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3825 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3826 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3827 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3828 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3829 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3830 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15143), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15547), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15219));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3831 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3832 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3833 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3834 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3835 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15400));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3836 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3837 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15565), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3838 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15574), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3839 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15488));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3840 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3841 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14995), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3842 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15362), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15598), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15221));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3843 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15514), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15279), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15136));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3844 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3845 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15196), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15422), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15055));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3846 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15114), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15339), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14968));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3847 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15490), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3848 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091), .A0(N23628), .A1(N23630), .B0(N23103));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3849 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15254), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3850 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3851 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3852 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3853 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3854 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3855 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15409), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15320), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3856 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015), .A0(N22793), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091), .B0(N22791));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3857 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3858 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3859 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3860 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3861 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3862 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3863 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15081), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3864 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3865 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3866 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3867 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3868 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15391), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3869 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15137), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15541), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15391));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3870 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15399), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15280), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15137));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3871 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15001), .A0(N23640), .A1(N21688), .B0(N23638));
AO21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3872 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15366), .A0(N21470), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15001));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3873 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45155), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15366), .B(N21279));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3874 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45117), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45155));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3875 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15064), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15464), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14973));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3876 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14999));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3877 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587), .A0(N23101), .A1(N23103), .B0(N23099));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3878 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181), .A0(N22889), .A1(N22891), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3879 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14966), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15090), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15231));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3880 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[28]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181), .B(N22648));
CLKAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3881 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[28]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3882 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15550), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15427), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15096), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15281));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3883 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15352), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15255));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3884 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15207), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15094), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15117), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14948));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3885 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469), .A0(N22897), .A1(N22899), .B0(N22895));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3886 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15397), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15374), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15523));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3887 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[29]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469), .B(N22621));
CLKAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3888 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[29]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3889 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15360), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15511));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3890 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45835), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15050));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3891 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15338), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15244));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3892 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15019), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15588), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3893 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14940), .A(N22850), .B(N23620));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3894 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15539), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15410), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15437), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15268));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3895 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15195), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15082), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15106), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15599));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3896 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15457), .A0(N22850), .A1(N22852), .B0(N22848));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3897 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14940), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15469), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15457));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3898 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[45]), .A(N22626), .B(N22624), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15056));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3899 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[45]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3900 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15079), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15217));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3901 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45829), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15273));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3902 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15054), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14957));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3903 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15386), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15295), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3904 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15312), .A(N22835), .B(N23601));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3905 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15241), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15128), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15153), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14982));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3906 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15573), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15451), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15477), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15307));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3907 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15166), .A0(N22835), .A1(N22837), .B0(N22833));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3908 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15312), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15181), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15166));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3909 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[44]), .A(N22585), .B(N22583), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15426));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3910 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[44]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3911 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3912 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15276), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15418));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3913 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45847), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15247));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3914 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15332));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3915 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15507));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3916 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3917 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15013));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3918 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15178));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3919 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3920 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15518), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15253), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15597));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3921 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15346));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3922 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15521));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3923 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15265), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3924 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15112), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14949), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14965));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3925 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15029), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3926 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14942), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15546), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15458));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3927 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15463), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3928 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15430), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15370), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15286));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3929 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15260), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15202), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15121));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3930 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15127), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3931 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383), .A0(N22866), .A1(N22868), .B0(N22864));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3932 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15099), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15039), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14951));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3933 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15591), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15533), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15442));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3934 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15448), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3935 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15413), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15356), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15272));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3936 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15515), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15246), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15188), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15108));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3937 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15113), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14997), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15515));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3938 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15369), .A0(N23608), .A1(N22919), .B0(N23606));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3939 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972), .A0(N22682), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15369));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3940 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[47]), .A(N22561), .B(N22559), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14972));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3941 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[47]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3942 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14990), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15134));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3943 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45841), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15481));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3944 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15049));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3945 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15212));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3946 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3947 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15557));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3948 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15380));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3949 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3950 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15226), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14967), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15306));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3951 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15061));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3952 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15227), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3953 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14981), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3954 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15395));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3955 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15336));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3956 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15315), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15250), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15168));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3957 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15175), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3958 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15145), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15088), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15003));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3959 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14975), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15581), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15494));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3960 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15499), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15232));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3961 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102), .A0(N22858), .A1(N22860), .B0(N22830));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3962 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15467), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15404), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15323));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3963 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15300), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15236), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15156));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3964 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15161), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15069), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3965 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15130), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15074), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14986));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3966 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15223), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14961), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15568), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15480));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3967 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15487), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15363), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15223));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3968 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15086), .A0(N23615), .A1(N22826), .B0(N23613));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3969 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342), .A0(N22672), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15086));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3970 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[46]), .A(N22554), .B(N22552), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15342));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3971 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[46]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3972 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3973 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3974 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15536), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15017));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3975 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45811), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15301));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3976 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15110), .A(N22873), .B(N23646));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3977 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978), .A0(N22905), .A1(N22907), .B0(N22903));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3978 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14963), .A0(N22873), .A1(N22875), .B0(N22871));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3979 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15110), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14963));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3980 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[41]), .A(N22599), .B(N22597), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15225));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3981 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[41]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3982 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15483), .A(N22978), .B(N22793));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3983 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14985), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15091));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3984 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15334), .A0(N22978), .A1(N22791), .B0(N21688));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3985 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15483), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14985), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15334));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3986 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45805), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3987 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15534), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15239), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15385));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3988 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[40]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14938), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45805), .S0(N22594));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3989 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[40]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3990 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3991 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15160), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15304));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3992 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15075));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3993 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15135), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15047));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3994 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15473), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15208), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15377));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3995 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15393), .A(N22800), .B(N22910));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3996 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15235));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I3997 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15152), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15057));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3998 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15008), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15554), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15578), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15402));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I3999 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261), .A0(N22881), .A1(N22883), .B0(N23137));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4000 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330), .A0(N23041), .A1(N23043), .B0(N23039));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4001 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14992), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15540), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15566), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15387));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4002 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15249), .A0(N22800), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330), .B0(N22798));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4003 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15393), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15249));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4004 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[42]), .A(N22547), .B(N22545), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15516));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4005 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[42]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4006 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15446), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15596));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4007 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15508));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4008 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15420), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15331));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4009 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15105), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15009));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4010 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15028), .A(N22814), .B(N22985));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4011 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15367));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4012 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15435), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15343), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4013 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15290), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15176), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15200), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15036));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4014 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562), .A0(N22843), .A1(N22845), .B0(N22841));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4015 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14956), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15503), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15528), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15353));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4016 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15278), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15162), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15185), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15024));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4017 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15543), .A0(N22814), .A1(N22816), .B0(N22812));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4018 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15028), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15543));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4019 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[43]), .A(N22540), .B(N22538), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15140));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4020 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[43]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4021 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4022 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4023 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4024 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4025 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15100), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14955), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15103));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4026 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15190), .A(N22992), .B(N22866));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4027 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15505), .A(N22868));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4028 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15052), .A0(N22992), .A1(N22864), .B0(N22919));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4029 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15308), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15190), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15505), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15052));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4030 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[39]), .A(N22636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15308));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4031 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23358), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[39]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4032 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23358));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4033 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15325), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15328), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15471));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4034 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15571), .A(N22828), .B(N22858));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4035 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15354), .A(N22860));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4036 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15416), .A0(N22828), .A1(N22830), .B0(N22826));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4037 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15026), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15571), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15354), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15416));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4038 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[38]), .A(N22566), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15026));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4039 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[38]));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4040 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4041 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15123), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15408), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15563));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4042 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14988), .A(N23601), .B(N22889));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4043 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15071), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15154));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4044 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15510), .A0(N23601), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15587), .B0(N22837));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4045 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15107), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14988), .A1(N22973), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15510));
XNOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4046 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[36]), .A(N22728), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15107));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4047 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23255), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[36]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4048 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23255));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4049 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15559), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15042), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15183));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4050 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15275), .A(N23620), .B(N22899));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4051 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15211), .A(N22897));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4052 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15132), .A0(N23620), .A1(N22895), .B0(N22852));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4053 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15390), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15275), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15211), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15132));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4054 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[37]), .A(N22641), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15390));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4055 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23324), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[37]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4056 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23324));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4057 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]));
NAND2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4058 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4059 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15372), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15585), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15063));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4060 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[32]), .A(N22651), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15015));
CLKAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4061 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[32]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4062 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15444), .A1(N22772), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15303));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4063 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23433), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4064 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15147), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15206), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15350));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4065 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[33]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15567), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23433), .S0(N22575));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4066 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[33]));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4067 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4068 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15583), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15496), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14980));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4069 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15078), .A(N22910), .B(N22883));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4070 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15441), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15530));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4071 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15594), .A0(N22910), .A1(N23137), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15330));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4072 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15187), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15078), .A1(N22708), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15594));
XNOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4073 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[34]), .A(N22533), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15187));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4074 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[34]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4075 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15358), .A(N22985), .B(N22845));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4076 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15589), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15012));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4077 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15215), .A0(N22985), .A1(N22841), .B0(N22816));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4078 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15358), .A1(N22764), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15215));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4079 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23439), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4080 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15348), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15125), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15263));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4081 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[35]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15479), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23439), .S0(N22530));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4082 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[35]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4083 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4084 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558));
NOR2X4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4085 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4086 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14944), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15289), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15434));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4087 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[31]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15383), .B(N22611));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4088 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[31]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4089 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15170), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15007), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15150));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4090 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15102), .B(N22606));
AND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4091 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[30]));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4092 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4093 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]));
NAND2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4094 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4095 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15419), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15173), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15317));
INVXL xor2_A_I14398 (.Y(N23929), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261));
MXI2XL xor2_A_I14399 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[26]), .A(N23929), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15261), .S0(N22491));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4097 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[26]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4098 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14991), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15034));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4099 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[25]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14978), .B(N22616));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4100 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[25]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4101 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16497), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0]));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4102 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15192), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15462), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N14946));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4103 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[27]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N15562), .B(N22580));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4104 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[27]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16220));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4105 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16534), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4106 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16552), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16497), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16534));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4107 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16522), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]));
NOR2X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4108 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16542), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16522));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4109 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16562), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4110 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16493), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16542), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16562));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4111 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16537), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16552), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16493));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4112 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16548), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4113 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16569), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16548));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4114 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16500), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4115 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16519), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16569), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16500));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4116 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16489), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]));
NOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4117 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16509), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16489));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4118 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16526), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4119 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16546), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16509), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16526));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4120 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16488), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16519), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16546));
AOI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4121 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16516), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16537), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16488));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4122 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16535), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4123 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16554), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4124 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16486), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16535), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16554));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4125 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16564), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4126 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16557), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22]));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4127 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16514), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16564), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16557));
OA21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4128 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16553), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16486), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16514));
OAI21X2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4129 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16516), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16553));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4130 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548));
INVX3 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4131 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0]));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4132 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4133 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4134 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16556), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4135 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16506), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16529));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4136 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16525), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16512), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16556), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16506));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4137 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16515), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16538), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16558));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4138 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16533), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16498));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4139 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16551), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16567), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16515), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16533));
AOI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4140 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45547), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16525), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16551));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4141 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16541), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16505), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16523));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4142 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16561), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16550));
AOI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4143 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16492), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16531), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16541), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16561));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4144 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45552), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16492));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4145 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45547), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45552));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4146 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45549), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0]));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4147 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45549));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4148 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4149 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16517), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16544));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4150 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45000), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4151 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16508), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16565));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4152 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16545), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16503));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4153 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16566), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16571), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16508), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16545));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4154 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16504), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16528), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16511));
OAI21X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4155 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16566), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16504));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4156 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16643), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4157 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16643), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[0]));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4158 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45000), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4159 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4160 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4161 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23240), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4162 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23240), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
OA21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4163 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23239));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4164 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16663), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[22]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4165 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16719), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16663), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4166 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4167 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4168 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4169 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4170 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16662), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16719), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4171 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N548), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N549));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4172 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45854), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551));
OAI2BB1X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4173 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16646), .A0N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636), .A1N(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45854));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4174 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16646));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4175 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16754), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[4]));
INVX2 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4176 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16754));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4177 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16727), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16662), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4178 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0]));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4179 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4180 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4181 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4182 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4183 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4184 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16742), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4185 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4186 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4187 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4188 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4189 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16684), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16742), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4190 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16684), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
XNOR2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4191 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16636), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N550));
CLKINVX4 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4192 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[2]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4193 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N683), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16727), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4194 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17223), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N683));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4195 (.Y(x[22]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17223), .B(N23924), .S0(N23918));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4196 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[2]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[3]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4197 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[4]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[5]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4198 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4199 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4200 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[18]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[19]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4201 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16790), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[20]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[21]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4202 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16685), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16790), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4203 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[10]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[11]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4204 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[12]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[13]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4205 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4206 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16789), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16685), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4207 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16693), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16789), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4208 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[0]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[1]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4209 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
NOR2BX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4210 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4211 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[14]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[15]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4212 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[16]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[17]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4213 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16704), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4214 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[7]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MX2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4215 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[8]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[9]), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4216 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4217 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16809), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16704), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4218 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16809), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4219 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16693), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4220 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17207), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N682));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4221 (.Y(x[21]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17207), .B(N23924), .S0(N23922));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4222 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16769), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16677), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4223 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4224 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16810), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16686), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16757), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4225 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16728), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16796), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4226 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16756), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16810), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4227 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16817), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16756), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4228 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16823), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4229 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45002), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N551));
INVXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4230 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[3]));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4231 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4232 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16705), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16777), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4233 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16749), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16816), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4234 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16775), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16668), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320));
MXI2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4235 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16775), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4236 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N681), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16817), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4237 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17267), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N681));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4238 (.Y(x[20]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17267), .B(N23924), .S0(N23919));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4239 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16734), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16802), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4240 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4241 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16776), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16811), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16720), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4242 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16694), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16764), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4243 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16718), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16776), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23322));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4244 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16783), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16718), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4245 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16795), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16669), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16743), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4246 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16710), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16782), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4247 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16741), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16795), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23321));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4248 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16741), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4249 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16783), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4250 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17251), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N680));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4251 (.Y(x[19]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17251), .B(N23924), .S0(N23921));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4252 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16703), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16763), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16801), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4253 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16703), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4254 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N679), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16750), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4255 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17234), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N679));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4256 (.Y(x[18]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17234), .B(N23924), .S0(N23920));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4257 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16667), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16726), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16768), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23320));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4258 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16667), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4259 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N678), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16711), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4260 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17217), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N678));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4261 (.Y(x[17]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17217), .B(N23924), .S0(N23921));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4262 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16794), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16692), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16733), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16681));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4263 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16794), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4264 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N677), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16676), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4265 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17202), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N677));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4266 (.Y(x[16]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17202), .B(N23924), .S0(N23919));
INVX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4267 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23318));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4268 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16724), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16781), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16822), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4269 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16724), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4270 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N675), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16699), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4271 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17244), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N675));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4272 (.Y(x[14]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17244), .B(N23924), .S0(N23921));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4273 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16691), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16748), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16755), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319));
NAND2X1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4274 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16691), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4275 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N674), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16788), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4276 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17227), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N674));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4277 (.Y(x[13]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17227), .B(N23924), .S0(N23918));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4278 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16814), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16709), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16682), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4279 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16814), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4280 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N673), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16717), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4281 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17211), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N673));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4282 (.Y(x[12]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17211), .B(N23924), .S0(N23920));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4283 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16762), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16815), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16698), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4284 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16762));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4285 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16746), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16675), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N23319));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4286 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16746), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4287 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N672), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4288 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17270), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N672));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4289 (.Y(x[11]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17270), .B(N23924), .S0(N23918));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4290 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16673));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4291 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N671), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16739), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4292 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17254), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N671));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4293 (.Y(x[10]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17254), .B(N23924), .S0(N23920));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4294 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16767));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4295 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N670), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16666), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4296 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17237), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N670));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4297 (.Y(x[9]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17237), .B(N23924), .S0(N23922));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4298 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16697));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4299 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N669), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16761), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4300 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17220), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N669));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4301 (.Y(x[8]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17220), .B(N23924), .S0(N23919));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4302 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16786));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4303 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N668), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16689), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4304 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17205), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N668));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4305 (.Y(x[7]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17205), .B(N23924), .S0(N23920));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4306 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16715), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4307 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N667), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16780), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4308 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17263), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N667));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4309 (.Y(x[6]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17263), .B(N23924), .S0(N23922));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4310 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16805), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4311 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N666), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4312 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17247), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N666));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4313 (.Y(x[5]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17247), .B(N23924), .S0(N23919));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4314 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16737), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16800));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4315 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N665), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16798), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4316 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17230), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N665));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4317 (.Y(x[4]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17230), .B(N23924), .S0(N23920));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4318 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17213), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16731));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4319 (.Y(x[3]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17213), .B(N23924), .S0(N23918));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4320 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17198), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16820));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4321 (.Y(x[2]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17198), .B(N23924), .S0(N23921));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4322 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17256), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16752));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4323 (.Y(x[1]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17256), .B(N23924), .S0(N23921));
OR3XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4324 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17239), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16680));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4325 (.Y(x[0]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17239), .B(N23924), .S0(N23919));
OAI21XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4326 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16343), .A0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8]), .A1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45128), .B0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45139));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4327 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N585), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__68), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16343));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4328 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N595), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N585));
AND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4329 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[30]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N595), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N741));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4330 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N713), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[4]));
AO22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4331 (.Y(x[27]), .A0(N20596), .A1(N20746), .B0(N20748), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N713));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4332 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N712), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[3]));
AO22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4333 (.Y(x[26]), .A0(N20596), .A1(N20746), .B0(N20748), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N712));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4334 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N711), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[2]));
AO22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4335 (.Y(x[25]), .A0(N20596), .A1(N20746), .B0(N20748), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N711));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4336 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N710), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16759));
AO22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4337 (.Y(x[24]), .A0(N20596), .A1(N20746), .B0(N20748), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N710));
OR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4338 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N709), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16722));
AO22XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4339 (.Y(x[23]), .A0(N20596), .A1(N20746), .B0(N20748), .B1(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N709));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4340 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17141), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[6]), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__19));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4341 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7494), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7381));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4342 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N708), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7494), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]));
NAND2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4343 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44986), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7395), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N7525));
NOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4344 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N707), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N44986), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[5]));
XOR2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4345 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N493), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N708), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N707));
NOR4BBX1 DFT_compute_cynw_cm_float_cos_E8_M23_1_I4346 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[31]), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N17141), .BN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N493), .C(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[8]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[7]));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4347 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45115), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16770), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16808), .S0(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16725));
NAND2BXL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4348 (.Y(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45148), .AN(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N16991), .B(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45115));
MXI2XL DFT_compute_cynw_cm_float_cos_E8_M23_1_I4349 (.Y(x[15]), .A(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_N45148), .B(N23924), .S0(N23918));
EDFFHQX1 x_reg_28__I4378 (.Q(x[28]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__I4380 (.Q(x[30]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[30]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__I4381 (.Q(x[31]), .D(DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[31]), .E(bdw_enable), .CK(aclk));
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[0] = x[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[1] = x[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[2] = x[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[3] = x[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[4] = x[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[5] = x[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[6] = x[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[7] = x[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[8] = x[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[9] = x[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[10] = x[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[11] = x[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[12] = x[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[13] = x[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[14] = x[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[15] = x[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[16] = x[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[17] = x[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[18] = x[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[19] = x[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[20] = x[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[21] = x[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[22] = x[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[23] = x[23];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[24] = x[24];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[25] = x[25];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[26] = x[26];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[27] = x[27];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[28] = DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__42[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__195[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[18] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__197[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__201[48] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__210[30] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_0_inst_inst_cellmath__215[1] = 1'B0;
assign x[29] = x[28];
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

`ifdef fdeQ_A_bdw839185604_bdw_COMPILED
`else
`define fdeQ_A_bdw839185604_bdw_COMPILED
module fdeQ_A_bdw839185604_bdw (
	D,
	EN,
	CLK,
	Q
	); /* architecture "gate_level" */ 
input  D,
	EN;
input  CLK;
output  Q;
wire N8;
EDFFX2 fdeQ_A_I0 (.Q(Q), .QN(N8), .D(D), .E(EN), .CK(CLK));
endmodule
`endif //  `ifdef fdeQ_A_bdw839185604_bdw_COMPILED

/* CADENCE  urfwSQnfoh9N : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



